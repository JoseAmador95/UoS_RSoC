`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Rp+DsHUrhAzxP/56vtW4aNpp/zu9s6ahaH7x428jDj9XKjNdq3fC6jpsidnR4fSCPXi80rH8vori
TrlJC5qZ3g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qvYoXgg1nOhU/NXb+rt6QgJJZKiUgeZ5UTBgfRDN1RaVSht+Pv31eM39uQUJOGuNRBdR20L2Y+Lc
FOb1ZOy8jRDaZnkfjg+U1zhz7AE9WOw/n0hhgV83S0TaVkNb0sL8SGahBoFZN5HZCJc6I6Czcy9r
OmPtfJjVaiKmU/9VPXE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uQQ7fUdn5jlignLBLwCLlA++9HTnI3hzv/Y2Gz+Qm703h9gQpdspxrNiIRx5hz0k/zwG2/dTD4rs
Hb51mJxGp8br8Z4KsNfiGZfRf1AFSUJ74/bdvdXf49ZioYhZKdRf9fiNorue8QAU6nXQOfNz18yq
j2V6/kCIlRRY22+Sjefz8s8CkJ7uDibyL3yD918ENcsMTH71O2wdHSccb0ArcL8950VxiSdwB1dY
SnPSUI8S9XmuYhJJaUIP7lNU+DuXS0EgdJZS9zVgI8IFS4g6Wx2gAWjhleN9T7xJIofE78qV8jpD
PpL60g6edT+Dr+RnQIQ0EqlwtY1UoFb/pmhHIA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LR3KYP6gUamfjjwvA27IVgAXkj4qSg+w4fDuW9kJIkkfiKx4zGyhJq9eDw5P86qvqfF4WDaIObco
St39dl5VX1va2a3fpCQvWLAoK8MRZ9S1pkUygcsmEfwvW69BIQWHHnzvFx6IU6pb5Wwj+iiDTQya
vSV1VdyjrJcUeqrH78RrduZz6sLj6ScxsnkT2CYMfVUuXbtwvs6RurW83YyhtlkmgACCsEXSmB8B
nf0YeS9dMXtIiWAaYF40xOHWw5vmdOUvndz8q5B23VBIWYZ878eoRa1rzF7s4NgcOiHAqb71bMjx
KsFiHu7mxrg5MXJOIz6KchGysDwxWQVSp0/CDw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RtK6li6VCymQ6/2AY6Z8sYVvFjwFRNQNf5OEl60JRkHwTHkLn9nJbLME2u3BYGmt3Cg31iDqZepT
BUJD//F2b5eEcV8VVVZ2rrwtuyU5BKjAgn1oq+XTFRxqluxA5syqL1GjimWjlaolmTnnZJothPHl
8W2sf8awcAuB0OVaICrq70MmTioKsmIyBYG+n0OR3szlktMcYoJUWENj22Isa7AhF7VYi1EpI7FU
i3WzMpTH2PjXRIUqaRsekoJwkmgCeRJcAOVZxPuL71iJrZalFWUYHbUIaomcHtQn6vd73iQ1C8dM
Tin2x/P69mNdGk8gIQjigI7V4wwPgXbRypNaKw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HKNzCjJC+GBAuCUEPEzhx59o6OLlBluyEiT/PXyp4dkr8Xynwjm/wdOAOj7BApwApstI7Z6QW2uQ
7Vcm/5AsAg1RVk7W9fwB47/lsIHfZNt5prsjqgG0wdxF7OZkc9eGwCHhti//lI0w/lA1D5w86QND
ipFaH3O2xKs5eIkPmko=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HLcBvYLQ3QNOA+nkrLp0XrM2kns/P1QwkwGWYvWu0xdVdjFtPNz0zk49j4YATTHw70LqFG1Mt17g
NwNw7dBXKMBx3OPguS/enpbOu9Lg4TmPowPaRpKsYNjpb9ZxJ+idt3VCjA5mCXFr2Hmfhvhg9F8K
fxZ4s352bT4o3mN/vFqhYp/otSUNm3SVcpARTEt2KpEVisOvSJcVCw7v9bQqQ7kM1JK7UMsSavYD
FOR/dq1EwasYWmm9M8uV4JxROgZOOsF0J1gMwrHcbNQeSaK0ACBEZn9YyAaC3oZPTLwsH6hFtkun
HkiWM3ZGvzW3lgSUls1AQ9+2DiYcWS0CaLrtjA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BF4Uj/645t1QRNO5C5i3qTLp+gWuAVZgeZUoC3kj4NE4aXABcHISqpmlbr7qGgG/Zix8eGWcY9WC
73NvYjs9Vq3XSMFWfWEGyeMaWg3cC9r3H19WbzRkeS4IwLtIvvihDGEwK+cQxiq37iV4Vs5LSYuf
rEendDB34vYVJmGNPkC/GRj6/BqZ/VwuPUUE+9Wqxu+DmXoK5WQPNwQzNoYIVPsg7wzc5hPA+NQ2
Sxuhk9BzhrgBiN1hSKglJmgxvCoAL43KZ+eigPDlBRv4IyZz6332XWuxmtc9vA/sezLtdY2Zk6pD
UrRgdKsIEM2wuQ+f9KnDXkf84NhM4XhUEdukvg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1559120)
`protect data_block
chrhmNL8XHPD29EwnkNNCRAGUfhQDhesnNS8cPLW9ylOp8bkWodbzGXf5J5HNCAwOgqiqQJJYSQp
uNpNgIzAqbsKJ6AGnULt28cMprL1jyTR2MlA8ve8SMzo0Dg41pR3ltav7uSBoSkfrLEVaPcGczz1
vrdLr5ZxPinxcKd6MNHcdHInLhsk5D7y6zxE3+894V3JJkjZ7vgCoMK66I02l/hvNOzUValPyAQa
hE/Heg4TDfjrrYF5DRbk7lOnLq7KSjB09Z/zXzPWC9m2LLfcAw7wfUsZQKxypYTOQkzU1AIKsvjR
/QxXBLJIPVXnHH4Hav8jIcy7m79XMHsTvLSmrtKODe+RPH7Z7gquY7cs03EDIw0G3aYncntVXKNl
32NEIwUxXZFZFuGk7H+PDJGANys4KhpoUougqgwLpT06TSipnFsWOAik+73W5TFC6oy80lrMm8C9
Uc+nMpAzJNOJxw6TTU06G9Cv2kPWgfVOGdwUKipIC9JhVSqK1RRDhByQfkyea+6zhGAkWQoBAyns
b+QgBtPXg5y7VWCASLCD0cTMpE8qdOOXuuPZuH6OgzEtRQu2Vm2xODIQcaHnPcJexKY+iNlsoEZO
T3eI1twKS8okro4hwtiyETQQ4cL8OQAPNi7ImW12KPmg4Waacd+JcBhzvkXlCJS3mr3JgRrU7G56
2LhZFdGyYykrCR1CJWdXiFuV/BlNxYqmepTrHF7k0XlNL31eSXjGyIaBuxwM6mEVOa3WBI1G0GMx
Hh2vGeCcVCDkOu5r1G1TVLNlKPbs9K8UkRnnLHKfoTy+pUiHobjHu72E64fII9EPqddRBm9Teapa
M/6kAv9LyDt+M0bsCUw7iJVt0L0vAco7YcI9vuluhJxShCdDomEWmeJDAMy6qk9OO92+thfMBNZ7
uQsIUHFp0uZ4ehIDLceLjSCwN6C3Nd4hQjWoOrLYcBumfBKs8Q/2gAweEdB9sarWAcBw4f/VfIJU
OmZ+4mioJRJRxtGFdJ5F/ZbD83CUzqFq41kzKApacgyl+g8Lj06aKiyC/eFTN3Irz6IU7mDdc/Uw
DrR971Nx8K67vZfRILBK0JrXN6tmWGs0CAOC48szLiuEP2CJltwIWTN6my+4TZE08aD22F4TGkjw
VvIDiu4VB5MXnPOx0jLOCbXKuj840S+THJcXouWcL1y6c+iA0BkM957U3c8bQBb9id760pIrWGcU
GGWBndVaZ54fzbKPi8IRHRm/3f9hlhYAW3DkVbJzDPKlheYawEgJuQC6zUnAWFHhtgz+imRSlWiZ
Pw4v9sdyQxgII96v24Fin903kJvYfgvyEy8xFQv+Pnj2MDSJqxLwqM9KGwr4lhcqq341XzlQ5GmT
rjGPsmrV132AcfTHhWb4YLb54urxk+ykCXDXFXTCM9JozPOqDn+lBueNA9QiIoOfChWG2T2K87uj
lZBLCo1RRW1YMHDN7uYvC+EA98JFVGtBs1CxmPOmkn+J+GzuNALT6b69zIcAWpd/2M/hhBVq7E5q
WBiaxHGPTvmRptNBnePQlhD3CA7z9xElv6rZRGVt2LZ1v0Wz5D/UZu2LTt7gvU1zVv9hR7oz7g6e
3ZYZj/E1kHPgVGrut5J/JvN3rVVD//5Put+9jFI/z9pNp6QgaH2dh7JgaDfQlpmT3d6ZrL93xOjY
fWgQRMPab2LoDSBUjsqwrl1LqnffTDysZRi6E5870dcO4TiYeaCjtSTMYnvu9IRpqMOqkHY27yGq
MYtZVF51Xit82GoMiqbmJnfugNxQ/1CTQ5Yfp/1KwIPrv5pp+6Z1Jc+ZxobPpL03eXyVtWeQDx1y
Hd92WK6mJlAjXDJAJ49isCWhDEahgsfejVlJDOWs5Quenv0Lg0BHgSMsZCrdVERyQ25D0hi1w0F0
8U3PtmU9Lo6RU7oe16n6TT/HYEsqj830XWOSVecZD0d3h07xrMATaeAPrp7vwJG1InwczyE0fIMm
dVtqAjAQup3QroaooRelVkeMTqJyA+Wbcs4DYAzXMe3lmkBZWwySRYLzmFy2nEBKXwCSvYWb48dr
tCspV/g+DENVwWFQ6g1VpR9pU5vwNWMLG8G3MweVV/99d8wg9LoGXfjx+851dPd5CkqxC56+clOj
0eCDCB3KMMvRUxVKwX9jIII5bK6HN5ejWXDOXg3sUy89mvvZK/h/HcWTaMCA13aF/7sadOuqwo6q
K58IkF5xJ7pppeRMWmrotvI2wlOl7HcjQMSi/P2ppwq1WuOmW7jh1SGElFlFTqIMvvoPQo5QKApr
g2W0PmbbYMg9PoJMhReB3m+OrGZPjgNCFceP0kuJK1wdykJwN5+CJMallMqp1mS0iAv6RUCKyJyF
v00usl1a80V8ybr0JgfDDxNaTkbCyCAoTm1LkZVVxZ6hp/01XDA0cqhesWWvgI/cUTd4t82i3Em+
fmV9pCbscSx8lTw/CePPn5LOC/M9tD8boTRjXsckmeR3vo3V8y+otKLK9/yyx1wxw59VlYRxaGrm
okHGTXY1Wl4Ou5bEstUAwLERGANUHx5ed9ehNpdUGvccVyC2e9z5nKgtKBlnWWAnl14ILUtvO1T6
Ar++NPX1UBWzap68wtgKwzoL7PswaECVwW6th6PnT8TyEqxcTybh67q4Z229B8XggkWaFW8+ZvMh
XC13BR9gkDne8hkEGZu5eugN1WsjU62dtel9Xx6o839TgahPudALswFzLDzyTAcAsQfxcI3zoN31
zbL/UCwruwACGfBwacQOMh593Hm5usLMCkmxVG8QYNzNg6hR5hPTsVDo+E5mXXxv/cdQ8hiE14N5
rLY937vdgfWvdef7/Jm77lu9iL7l0YMbGden/deaj+4kOoOmbpr3lzGQ+11sJNXZMPYszOB61pBD
JETwaVvSJGxHd7TL2pI/p0DBHQ6Jh7KjyZsWaRlMAnSsbcjCayGwIaqBdpXKVqfkIYnNDwVv36SX
YQogapbBm/AWgxQnjyAyYkRWy0kr2kSPaolIpvbmJ8roVZXlfYzX3DL99XdVWgiyxJ7U5O60KyYu
pVRk0KjnDHL+Nzs9WWq+zsL0hapko0FrbI/Jz+xbm1gOKmk44h8cGzinoq2EiJPYvBk3um4W5sqE
YHqKXJLsgVQ6gdz+/ocG1EjW8CJt2+lLSK7mSQsGr/CgRN3HQE2oGEzffXPI9TkIJyKkZxkc6gEU
QuyyuZHw6OouwiDxAXZ/YlqgXv32cPbuW2IQBscfSZv0P/9jCcKd7QyHwqsLk9+QB9aHg9QmQmD0
SFZbFCOKNrAO+fJX0VofVEC1s3XUA0xr0ntSkVsQFdKA8XumkCesKwQGrKSPrjHvgwhswj8miSDG
m5qwni6XX9sdNggGA72aZotQA2bsoFS2IWifmApLRVy+Rxya2p14Hz8ChzZSKhtIlruruhLuxj56
Vb2SNi6wAUT7QawyCPzXIbB+K63gsFUTPigeOVLAaDb5X1T7+M+exPq+uOtbQ2n55Nr/wRjx/8Kn
WaoQiAVxLAHH1fFwm0Q/Bc4VRJ0yIXQcqI7yZY5YqXj2fd6Y6+zh4exncS278wNd9gD25SyGGjFn
wwDsWwJMiAk6Hkxv1RMdeTx0A4cRl8SwWIwngrm+Dlja70YVM+U1Apm9EfF9zkefvwreGqQozPz7
CLV4tb9lFgtP2r42G2YBNY1VtqqujNE0DZL1vAdZPmFgYguqE9a7kffBBmJsL3AW33J9T+MAtQLY
4kQxZXbGLb53CV23lm0GaI7MA7n6Ks5h0OPWidbLlEHJ1mffr+pNCOmHbZH8PVcYnrC7TKdNPV0a
aUb4w4+5n3+joe6lefSFZYNdwp29uL5SZAQUSJklPGC3d55R2BzlDpayV04cU2ch86SNAOMCrrm5
7PtwTE/wMoQjbhX1Hz2DveUETVXOE7l8aoYDvyJaZlqubQsBZ183sIvsRY39GytOH1FwKidmJI3B
xqHbOtqOhwGUU3wpuujoAHeZdh6UqAj6JM1ZQA2ZnDrPOMfOBQ4t9RNDR6yv5Vekh7nzz1JmdMBj
JZJxZxolq3u2SNw9gYDK5ZRSTXx1lEbbBk6kl12M1JVMATr4QLHIRY8+qAg4H6mhrSNz19lQctzH
5mzQBXzChxf2wRl7294O8YAO1ePX2pDiR8NZ8S1Yi1DWSjPYBovLOn2A502CrICOj2X5yOfKRMXN
6g62fRzfxfGN0kn7osarC0cjL8wzgoMlswwstv8CGg/Rjlph59gfGcnkpOPbxX2dA8CuHhzboZ4f
62XlSa168hMOMxCUxMtrzWYWOQFc9SqbKb+QKGY7rBhPFu/QRvzg5ZhYuu6UJG/S2YbOE30jzh9u
vG6JPYWyRfi8FGSQm4uoZ20gsj2JZR95gDyKyTMspAza86j27FL2P+992MM6DJKIkMtwl/v2EYaP
5t+K0HDwyESLhhJNmCPeBAK3CfJc0eAgHnC6NdlpmceQRPS9N4gefw6Qk7v2ADHicEOzV4jbYTm6
ZTq9Se6uyj3HwpWafw7Bw/Q3bxdxKXoSHq0u678bqUwKefT8XWylw0MrdWagaS4vjPYORN32zU1A
s44RK92aJ1BGpinFmUHKhQB+AxEfbtwqHbRVULWEuPPWPTrar6OrBcSkKPTuaBFfkziLaI0MvKPC
yudntMnvXAoyz3M9PC4ykYQnhtPBf/GeJVdo/qneZiQRoiD42+llLorgHCYDOmqjJP1oYkwrBJOJ
4E+feo3R7PYXPjk2dGvl3z6oH8mNL1QU1h2SZPh7LSb1cM8gi8hhpiAL/6xJaCAbJJYHnoUqAa6H
PU8xzG+xPw0KuS5IXWggNPYV+k9eFbxDGly9NUfVNySfuoasOi3AJy42eTaSpRT6nYezJsdHX5VZ
oVkxYc8bbv6SqBwFOgp7S/10QEHGnGozyXLClpqeWz+hoO7eDP2FO8swE+mYr/0E3zww7nr2VO1v
zk5fqVeD320Rmts9zQWjkTBzqBs0ypWVufLx/P0FdA1PcddUsZWZsPG24iyd7Wck1jQf2t0zibtD
v1Mp3NIR5fruXNQ5Rg51BBgMlBeeGB54j2O3WexwMvIITrq5bwICHo2OXCqcZ6GFg0DECNQOx5uB
zS0XdJc4GkZXNlquKMKAq+H6dP/L4JRv1qW0H4hjKBAbLSl/+MqCNx2e+peHum7oGiu5IH9MISLQ
Je+SBqd6uhlZYbUdTe9e/sP+ZlYMGvZPfdaNTXJQQ95gVetBjpIHbrmRqll+WfyZ5JbfANbyTq3O
K9D4O/28lnYM3yi9zVq9/KMmMGmZ9wV7IgVS0Fb5mWZ305Jupo3WgVlEbEuHoO27DINpAnaGGc9/
QxaIjBQ4o+BBB1WOBJBxHvC8z6SDu5VoygV4oDPRcHlQir9HB1fjyIgdyTNOfiX7u95AAQyvYZ6T
0tvIEcN0/qGjNIPgerHbOvKssH95/GFTuHuXzSOpJnC0LLmxbGlXtQgV/m8pBQqfQsTeB37NNqnI
5NFrXfsi9x2a3sPdJ0XX58lTvckJCvAohr7avZ8yLvfHLwgSA8jf4a4k0bPssIrH2QKG7Bt8uyvk
pPGlDNlP7+mWuKDx/qYTNqHv8s5WYx7M2f0JYMWA4C/DobkIgfTOHuuOEKbI9PQvW9AshBiPHmWy
SpmIdzFi01gBjPRuQ5b02ilk91JhxeFT/puzGluPHJRLl1VaOcA8zalhQ8a+d+7HscsAvQqADLy8
l8SLAA8b5BytmTS8p/auoVZgaqgGCwkixg8vE9m2IJeZHbIoS/Cy0PThfSehFt4EyHJXqlYlwfKB
sT2LDFT1Pv19fBexDO3rBXFbU/6kDRXNJO1gRP5yRbOfHPOIKLOGX/Sqo1sXdnMvNPGqdIl0a/Uu
bO1V+etvvWnXxOEsJ0lA5KFGdDybsucdRvAptPECzMGzonjFNHdoCQ8ZSL9orH/iEcYFnZI3ci2r
1AarSzMpuQAmR3IkeDbAdExXWAiuntf+83lS+4I6CKkqiBg0becyo5JFnHfEgeTbwCopkvYGaL/w
5JrOz/l+qjkKqjm/ojft19jKecBVtt0z/MLytUzRjjm5oidytB0NKMqhRF8uom82X9sl46MtQ7OX
g9bdNRr9ZMrDqsB8KI5CrKBoqF52YSU4+d/reR8xhxhnQH1Sox/ZLstbj/ElXSYtr4MCxHR+c+e1
iJV0wMjxuubBL8TViV4wDbCUHNtqvMh3+XwWdba8ESLT8CkkQNucoFbKR9wwiLJVcyhDRNLdXoWE
Beh6iE8kEJyXBO36cC5QHFfe0DGPEnk5et3oHG+LKFoPv5Oy3yqC1rU09apfl7ChMzIKiFvy9Dbe
tM0OlCrZOsF8GlXgFkjqSx3HyMgoH+9XoYvgEAQ21F/MuPpgLFNGnI09R2ZLE9Zw59Fv0Y2nRN02
BhymzQSBoT9ZysuwdfAKpgwnnXhMQ90xHn+F5iP/PL9w7vLW9VDylgsOHaH+NCqq+LI8uxQG4SPn
ArB2Vmrov7I0hsvfC91Vagjwyoa4UDRUhhgRV6LwXkiFF2SuCe27gWVkWwupTlz3V0uC741bKths
fhXgeSJm7LnVWKfV11IJOJMZyUBz786+Ke6i1KagYxIKY9FaKiXWOUwrtCsB97UjFMWBgPjc0Qyd
GXrmrl+EA0UmxH4bx86UF8/SrWMKVUO9dgD96sA7wQNWlOr9M1r54fkf/VaeXwGB6gp8T/AFhr1p
u74A0QeHBLD7tQHoUtFNhVFDUg6Gjkio3YvwT/osVYSyGAA3ORi4Eynn72q9ADc4WIpJDacMjaBU
tjj7MwjUF6UBvijhRXgf0s+vTAQiu4OhoXl0Enr7LkQ4Hw9nz0lgy+5o8MgNX/yEwarJx7gJZ9FY
pgqda0NxQnmkIlLyeSBdGZXjZ/I/4Rf6f+Fr2h3eViovgxyyMEPXE2WyYjuQ3Z6cL+oG1O+hMPKr
XZIwbBaNoU4nkYe0e1R6+GZfSjns0lpngXxof2y1Zdu1d+tK2BOWedwhOtnLZANlynVzBL8lR7LU
Kz8BecS9UG/ifEIc2Sy5zO7HB3/9LbkSAz6/SAt6L2Cz+vYCrYxW85gKJX9B6ZL6UtCFmTytmwsH
uuqpR3IbXfVTn50l6CWBEvNpeqoT3BENcR9sLyV8NclaFpXkc0LauStBn4ImKCOOgF2EiXQwETcz
PybHZR1JiwwuXXQVH4wG3x1s9273WvgbePOn9h8kZABn+aMf20sdeApcdt7Nzk1jF0PWz5opIg1v
GqiccMwjDmoc6JEpaGiU8eZVV8tMlTn/CR4GTXkrPopNH7/wP4qv6PgMgLrOG2Gj+0uHsYLA0juC
xJI9Hmzf7ul5/5iAQ/py+eUCK3x/RAFAfA12IBosKWZMMI9OBW9h8ON0KncvpZB0j7ouuAP3fB3H
i6X5Gg9k34Aik+6/37S0skrW9GgMfh7XIJRPw8ApmQxyePb6Zi8ISAmUR5Z5zL7Jv72KJvZzQOqQ
OUA0HlrBKOdPFRyqlZs5F5Y7w3uy/Q6rgmFMd3V6cndcga2udWx9g2NYiIbVxVPETzSKoLC8iB3E
OihMmU091Co2Cz09CVZJkiU58jKoMTvRbGzOWYAqq6jcpUFg1N7g+I+fbelMrlanTg0qAd/79SBU
fuuPsZb2MEds8dIVEFD2lt7B8vrn/vmr+ZEjhLu0dhmFTzxYTx2PO9jQSMy77IsJqZzyGJU/Ovrk
HvwTjup1Jh43JsHmWBngQVa2PmJkfCTxJPH7qGn3lJs2bQ4sonrgv+h7KT39eAHU+wb6WLLWLEJN
Tz/r1+7B/pD1oF2lmyQ7BCq5Ap7rQiNZHotLzBjpHhW7JcTHp1Hw2V/CMQYv2EMnx+w0dQ9cPyGi
LRNCjXKmbgn0wueQfRtr8Kx6PRMzNCIj5jPp07+89h3s6rhwJK3y8dZIjcoBzeRTSbhFI9JXVRSg
OZlvA6ICyX3rGbwbVxszS7xbTGuLEtseOy9lGm19Chcjg39Rcl5XTIYHjW71asi/G8jEwHxbsAgj
JMWW1B79ve25Zpv3opRxqS/xEh+woGY5wLahgihDfh78K8Ppwa8NR8wTdAXavIvPJhvAlL0j87w5
T50lHX/2U+P0O1kdBG7rCedTqPwUFYwke6Z2ZYg2yxwdEoEcmJAzlBITJiFA+TpFSIpk7AklnCqr
VPp4C0nBgYn1zlCpwDU/R0tsPJ1dKYtXPf+/5M7uLqmQYFgIichCMkUDSVB8yEX37o0iEDsXHU11
u5eUDf94DyloMwZXQmQ90RYVR2EMmmCpKul45tOwLDiluTdw6CODaZeIXuCxd1eGGiAa9AYtTywK
oC3KQE93klxhoumA9adE6wkEzF3aWoHKK1/1e1YOj+5OhfTS3XfiBOqsE0FULXuKKj0KhuX5WDyt
cGKQzQMpwtWs+ugOCa3s2+6COJ8UhkzRXpNOaZZGJEJSSBdeZiZhhmWRv6Jyp6DRWvXfio+NLWRM
eoP5ly4yPfnOOw2rGjcxIRA4YZwHIxFteuZqfkwIi1SIVIdEME0YQtNh0wSIOmMPxuhmrCr+ptUZ
h4X0VnONrxYB8F24KWLFIm4P9TZ6CuIiIMLFg69HWZe4cPhEuDKk68Tm2IeDoKHrtrGAxji/3CBx
/hR0XKLyK41PivAX+5Wtw9oG4hvGm5kX8DElkC7fuAV3vw7tEmvYgBbjl3hC3ryFSGaihfeRxI/D
4kShNyuXUEAt/Nk2G1gXDBbPSrVkRKYuKv5qTP6HkNAOElfJqHxVc9GXXhPYJIhrjdWpuZWVLdQ7
1zs2L6CSBRsnmqTkxqGWZ6Y592wqKp1Y5LJyJ/0JHz0B2ybmsR0H8GCcE2BdvcjdKnzzh2s3tyWc
S290WcgrLWyG70R8rqodLSjBUrxUPhty8+0mStkzE5YqiGjuku60xkXCkBtUHGPYFjOfk4o/oNF8
ae/9ufh+r5WOcmicZhaqfaooOfpNBvBPbHSiLLlrGxO0BfR/Abzjv4mzEp6plL70kwvqPu1q3RZo
EC5n+g/iVMv4+JU2VWUVv8ew0XGNiiYzVyOFjFbn8ctczgNlS1QA+i6dFb1ITiCXn5k9AuZzcAqC
zz7CHULNgHwppGJaDQxmRf9Iyk6MCGmz2qiPrhzPYexAgdAwJLfNmjHOt/UXjIOpFQgKoLTPmtg1
Rb5eSTKWdHNIc9fNemIF/TEvUGwCxMKuXqPdyhfQO1uZvyre7YB7dLx1fX/N19/y/uQx/YoA3Jrq
JwbDn6FaYSu3FhiNlJikpuTo/DJwqqo6ZRB/4CZ0St55HxuYl0JA9zCl2RCe0GhJYsWwm4WXA52z
i2/hgZqJj5YZxjAY3GDfCpVnc2EqZ+7250kBLuxDDcSknDiOpFelwvzDDRvo7dl+nGm5N3pEx932
JyguOC7NuzpTYqsY9buhoAFrqpN5blLnKS7Pf9Qa4zTqai7AcphPmqh7VznHhr0WrtQ9z0ymhVqu
jPARc6X8b52ldKgs/EpCR+JSaNipdJMhZMuYn3ZFf6f5aTbCa3RIyryTH18P2OCv2BWE0aUa8ZfU
KoCd4qoxDc3Erdzx3VxpDe4raI4z1+v8dS0N66P2mfp8/DI7C3SHnYB7RW2Gkminyb4PIFpnks20
4eI7q5YaWQxs7sBNKt47gycnOEckmcDmpaC2/TFmNC4mKAjEMkc6c3Hxn6HK+eZAUa7LWmj49WxB
nSqX2na632Fz/ciuLHutGYj+qEoq3G4J0+1wGQLAd2rwD8eGje888e8iPEP00EBDhIplwQV4oy9Q
w9s0txakCPzNS0jRzNy7rDlREozxrzIRhlWgykkBboZBBBTv/uwVXzUqBFUayasoK6eGXRtEEkPW
Vt8BtFMByCUmAT5yl9sBciakjD+2IuDUaIZQAf6NripdDk5FFddRyNqPDKmPXMWKyD05hk2BecZn
dABGRyLdEo7UPNy3Ik6YgZa/bEjAZO6fTF1sIF9JjXsqjMXud6dMZZX5kHPqqQAKYxrmEwPGln0m
iQzDScCjnmnoATIelWFSc2a8rBB94JsulRZdyAYqPyRV7Y+bQxNBaqTVlljQvVebKUE9Y/XRACB5
W+uXw1XeYK31NKCP6Y+hhecmzX0gT44k36KDprNIYwf/DxyZ4tlsLTaAA5KN1llLrqFT3hR6h9y8
pFxraxGLaU3Qet/tnazyAUI0ktBe3qZzJElows3vjsrmnsNz+aIwck2b80Wy4zDEmcYSK9xCrBGw
/se00AZufX7YsA50+4MPsFTDZVfLwLQmCDuHqI1BwO7dvIrbBLpYei7x/umD31vcf3RG7ovUBYO+
iIiDKV/b4XrfkLoR9b+y9155pCXAtSG6EMJe+NotcfN71EXx/iVFoWRqIYUrLd1peBoIqgW+I04n
59+0DPe4xK22U8ORJqowyW32SOshyuZ1J/RQK8DTtjFRZ1jpU4SXpzSW8J4QeENFTo+Fc6mGOycS
ulX3VnB2FWDz10S57J+Pb47S8YNI/EYbWjDE4+SnwnLInefDEtRLjpamTCc1NdKvP92ALv1v8uEf
nU8CCuXWvXG8LbCqY/tQalkWrCCIVLsKwbqQzwREHCbLukMUzqBCX3sf4wmUOiJTfBJpcuOWSP+n
URL8ACX05wMzryFoYXEM9IZcrWUwF4v2iIa0g7OYjKM+Y59p6uFpQIc5xR+nptrRTMmw8YKJxlRs
GajG+u1Xule1Gpo05513ymI+hLrBplQ5z7jHF9MhlNrZf/cXqvkDM7TLS4mmvGczH93VRDcjwrLK
15m6EyYe7/fZPRB79VstoY1t6ulkISbInnHR9x6NcbE1MbWJEP4mhZ1o2+vVdyDYQY3DtDkgITvY
8BrTTuWt8poqHIK5VV4zjQUz62rf+4W5mavyqs/IaEdUbbbjG4hpJUAHG9N1lUh9qykOOP+h86gn
aTBGAfYpsAAefFMoIU/WYrzDfBgj4kH+OqnTk9ljl3jJcLUNloZCjHgHFxocu23yvFxuKkQhfCMs
yeuiFT15NKAgv9nSAzVu7RQFDsPDfTScI1vZVIK1SlgGUCg2DyBo6uEC7FrvhmiyhvRtnszxhG2a
0eXHfNrf3M1Rka0jab2yA6/qQHd2Ko80SPlOybaJJQAPg+7EBSGZYu9hB0+L5Dczwqt8KmKgwMBa
75qOeRBlc1yEOWwZdDJVWoPF4QzQxaKv7lYN6gR3K8Sk0ubByewCMyZK8JFxFKPZUfr6AGW2nRHY
1zabkWErqX238RLUep4220evxTgwelYJYFVnV5gjYKCwHUZ2iFASHvg1CERmbR2BiWSrYOA4xdnl
LoBdu7BgxYG1oP5Ab+Mm3SobPCYgxqoHlDbgmFMLZ7DOQy7kf7xjOWecpekqwSJGZn8JlG0lk5FB
Is4v0L5xJAZyGmGjDqXZxlSElW759t5b2AUNQliSkG/+rtayHG3aKxr/1ihouo9L63AuRYI9a4dC
QR81/bpnEv1l7siuLLyJYVe7KA3GYLbDYaW/e55lQ0HALR6Nnlmt8pYnWA/8LKgp0O+hNVUj3E/L
F8X4qi+ehWDgWMwFebLHB1L+QoVCKz4v50KD8kRI3rCEVZuMX48YKC1R6FeF6FuzVlsmLesDc83z
MBLjZgnJ0dkejzqGrIlY7+qL7wsf86DzLsouT3dvd2Y88wgHhoEECrd10nEEQSs5Fxwodi3jDhnQ
y1qAlWDr9QmnM99i9kgNLk1WvLFhtx7iiLcglnbE2PhQHdNFKdh2CVnq2VMQ39PX4TrWaAgBSISn
OHZ6+FZ/n2p9GZ977lyBnSfongW8+mH5Pc7rL/VKqJxsLT5ww0ZhGp4m+BJgeugQMGz5J+annHa1
FI/Ng3Jmn35kOyQ++/t0OugXx4AOQwO0iWjkPkxoDc4SoOSiChma1l4NEq9DAN5pwPwOcOavQTwl
nA5BUtUlGwYHQqjqvhXacHw5ZD///4m9Z+ZuM6ekX7cGV9Z3MlbqBSQNnevjoCw/gFViVI4UQFoE
eVNYiJkL8wqED0Pf6qIb+tRA3YPZH+w44rWhPjAptSVbIiTJosl53sk17qi9Eu+KK3ZkkHsBqWee
dOSyW70Ol0Nc4iBJLGFJOW+1D9tdpl0jftBVMy9u1JMhTq/Dh3uLFIXAnZZD18LYjpLUk/yQC27n
sPuzagYHK9qG6FUakC+1g6pA5UBFgX22ME0IuhWPEXREf3rUeYdFIoSWwD6A3Q9pTaZsJWTS2tIZ
zlSzul4Lu3nXhrTRxdYGaZ0BWEa87ePctDLqBLvEHDTTIXWrsCYojJdqTIAtfCU7pYrxirTctaby
1lGO6PDmEcxDNSV95FRW+Sq4a3DpQ1jciLTWo3HJYzJi85M+1nJFoBh1+XJchVcevcnTuvlz76Mf
0VnBYO1qrAvQ+b7tXz3jfoQRsh1hCAXNJ/L0FCloQQ5MLiHuFqiHl6Ohw1E2bDCSabtzxJS/+0qL
NUdKUjLDTSHpUc65AHx7Ksn2HWXUR1gKN4pFYpbX7UPRwYbvHe7aiQFEKjjYt+ALuCpcTlH4e2pU
tUgEKwG2SN0OG+Q7od7Slgw4MUftova/Q4k+zEVcMAuksUMiDJ7cutmMJBZsB3GqV+DPRwFe+Z3e
EiC2eR2aH0ZsCEWrHAXs02SSJaUxzmlLHT68gBrZno32QrvQcCyjCxkuVpaqYQyfOy79OdkNq9qW
U0uMSsYAyhV2DOduG9iQ9+vsPmHbBIKNY0eJfi8jvzfI5cPkEdFgedkWYR6zMC5wRJq9ujinrNJT
CUzLizXMdHNTufO6m2odvSMs/ejqcL3W3ihbLAFOSSPGA9Qi6hZoQ8PLz7tUEzhJCjp7kCc1RPIU
0oqgK86QY9FgeL/LPhE38g9q0JCNqR4XaT6Gd/UzSqAJdRMFKQDyNuPQq05ff+zNxk58WAPdMIHj
QuIQg/lWXuGO7rRsFgYp+Mku+jy37jX3tbZ3SMJGHV9+nCCjM+JetZHGIqdHddpczw2HZrUcl2s4
ChfKYw1q85VqdSwWU7xQC7y8gL++EQ3LGadLYsCCwJmfmR56SLUDB5vIVseh41zJZZVa917qiwpe
h5PnyFOEw+ZktqNEYcWhWE+X2gFMItvgPkcw3RqnfZh1jO/ObEXIVzlN8iGJAdQO1XWwEIzNa3d3
UC+86OW4qN4gxVmmJi/s6Uv4BQsvmtc6rguNzH4i0tKI/aW1LLkN7PVUHUG2DFbolMY/nhBVqqwc
D/CRU5sH5wAgc6Q56Z0kkb3EY37cb7MRPjrCu2nJSPwiDc+56JikaLYRXthNNB/RvbvOd+jtLCrd
srlgLz8ArGECl6GUrLO9JLujtHqg/VI84x7256sGv3XIlonmDgEV16aYjIybJe4cJnJNGNwt8Nr8
qjbzFz7l7hFe0Uuy+oLj+M1F+MJbhNLLKRRPz0lY6cWFmCf1RILYI6vRwijEFkfo3+lvE+QkkOFT
eWN/ZFOJq37D/VOFCcudmGPDZI/krUXy9QPsIitKjcwsI7mIZHyhUub3nAr5vim9ogd11ZMogdPU
rCVbuJvwwS4RWc0GIC+vxEKvDZ8fBsF6XD2dWjb2Dw7ODq11u9osS8uo1uQ9HVIpc+C3GJGLMidj
NpB0XehjxQFMz0fDOpWDmwXWymO+y3hY6GX9AuKT3kOQh7jBieuVMCN2mEPsLrGiWoO23+OmD4vr
XqDmBTIhEEKoXU5jBKjM30mxneSW9FCLsBL9Lv2I68Er3jWoVsP8tz0j2vP56LbHJofNeqVYQ9cC
ET7kDn2JbjEY8nOVfhc7asIDnX9oswtMQwxa3W2PIAJ0m1vAh2ow8wYdudcLDr+yheomNbWCOpwo
7FUsAqlW3RKyTOOAM7/5KAWkno9Il/ubNjnOM36IGBMsWXKh9+bukB0IZadz5hiTrGvjHs2pLy1a
6leJeDlRKmSBRtOM9+3JLOMJ9j8IAnRhaGWRYy8GddyQQ9KOyWLoEVVz05NKN6qf4g/1PYbXs6b6
B/7w+Surl2tvk52z9uf9c6JNbbBI7mmw4O/0Fwc9Ee1mRzHr6R7LUshvm4SgoIFADqjq7M6WrYA+
QsANrH1NhW7m4kCcR+F4tQbLXbcKw5o1s3EcGcx5Av5ent78Ps5ZAq6CbTXBlD7JuNC+8Eho7Mwn
l9rUGyNzNf8EFyAOtfoThev0XorW5Ae/YFOXiufA9MZgRth9zMNhyKmfD/+Eu3oBw6EiSCXu0Eze
sw7O9ARXEH1BLQqME5f2IKVPDkCr/9MtCCWfIc80kdQUTGhL2YLg5J4ILvS8sP2m+6H9hmGxB7GR
QcH3Qv1cCdqiBzkelzjO2lHiwQf+ZibzNjCIJSjasyoNOglKzZOT+NGHtYVvbGrYMP+bzRWRKYpc
7X41TiYl+iXuImx9rpargRtvFiENSBc0bcqbVme0JONhK/Yi57+f406rUWoP+mU2AXc3i1B14twJ
7EFtwTTIYpksVmd7yFPmLjCvUB1eCY9J2j6W8raWgqZI3f1z1Z7hcKgSCYlBlP6VwIkWglrhTuML
Exhpc0p/2c7v0YhAec6AhaeuLtpqil4j7pUBOkemZ3ojf98AqDaX4g96HMfU6sIfpQxEiL+AnTP8
LFCyxWB7Z1Z3mJ3Y+PYSOGjoM4UIxg3gBL+SZ9MceRNRoG124n1Ie60UcAGveAZkErMDNfyNmICT
0Hv5Sgslhohv+W+s93zsy7zW2qKVJe88UL/zKGcipc0vTMcVmBB1CHE7n2sLXHwsy/+T8KmImN8E
WFjnzxo3EWLArgU4KBcdJhXOEvTT7bYMgxxJDps9J9O5p0zGlkr5kEeXWPsjr3ZbZBOdlvDP6SxI
SOIc38PeQcvyCbwdfn8R/pShCOnTr/46FCJOIWttqUwzPoAHUMNqUb/oEWkDxVyj9V94FNByoyxr
1KPDwwaA77Z7nbxXjAZzmzKRPAk862EE3TqkCtrTE7KNf7LkNb4Q30I7GVqlxskDlNdlLlHgZYOP
MPzSigMeqQWJviqAnA2laykLaF/8mPlxSu0VQXbdZmc06wREUshcIYQGgPYGqmpXC9vrsKBC0o2n
5JQ4mR3k/oN85sjFN0LyPFdwMsJ4jGB1CdHFebBRkYIniySV4UT/b0JOiHPwkxjJuxe5zM6AbE68
LPJyUkRJR1FUDtN71zg3afE+u200g6eJlFoHvm5RsWwqy97FgbKVXi64VsmvnE5SAlxO1RgOCqCG
pLfMtWmjV22Mcq+L9V8I5Vkrvc9f9N9UNqgMdpl07M3mumBJRrrpksqFijcnZgi5cva/So0p6odM
Hq09mVfK6drtlo9hA5aosR59DSx5asgUvPkwO5x1viwJkSzi1unrSoePMr3bTv+dPcumwn23mKYA
iqCNqpno4iZpLae1Mj/lX+mEHA7DggTG3eFrZiokjsRWFQhP2VJIypZ8f7svYGxH8sLj2mYwnugT
6SHZ7YOuhuoEMzVyHLRYOABAyRsqHvYFkV2iBOuR0Ac6GLgEk4sGoDlELw+Z+uUyXP8r+pIzityh
hOl5Gg0ZXut+txUnggX0bSf3oF7QgLtlLHpeDmNDr/TuHNIDm5FgbMjFEJ2KzQVIUmmqYPa3iN6C
kYC+MiIK+bFg1NyZX2qqZ00OX299PF4OXtpmCYYYTJ3HLvEQL6ipWq8MQp3Q/AsEWAAcRhBa8aSw
hy6JrnE55GYZ1rwOZRDjBexWYFoLDSUlqx+edcIF6TkZPoGxXBjVEb7k3pkmCNrDMovfViY3tuHZ
yvzLI4JNDHunL3QlM3/gwtXTxKFzVRYYYVDRr6R2XIplgjcA33kL4+pe0oZYV+HBJIXwWyf/V+Ak
3hjRKN8xHteSaC/LthNSY7/CDKeXyQAYRgFaK7/wUe0PTjnpcXHYMpZx8cDgKzIvCPehS2o87rSW
fs6/09EDqWF9Pf048zyptz7+Y2UmwNOIaHwMqNeA5ph3KZ+IqBRJ8GRFdrdCvwNmAb92XsxRv5Vb
Z1SQcsmrx/yXNqiXk7WK7DYaG+32xF4UXV+5IoVGsGUU15O4ymDIzTS94yV0vX/XRkxy7Pin3IqP
D+KYYDzHbSq/T9j6NIXS9I6bLcwhTyR81oV4UQH9qiLarb75MgIx2tX7bgvg5XMLvYJsElbM5+2Z
Z2YEXRm9SJTZFsTkEtikdgmfUbAWDKPyir7WHm53TFErBLjwVNJ5DuI/EFBKbGpDPReI1n6g898h
IMKV/ga4k4QLPYfQ5yDj90P3F4NIkN2fQT5ZnYhg/7pXNRXhHJH5w5yi4KN6yDpSDW44Mdmqgi+A
tuvWSNDue3CvmYINJupF5ULOJS6Mq6zaXuZ4cIpb2tAYdI+/ZriGYuI3XRQhVgEYqwSGenTjVATh
7N6I0VIz4ycy4mF8ZYM2pwSKX6s5AFmVisQIS5rmdwYO5GAuLefbLGIhdxx11dXsB6gbVzCl267u
lBYt8yQ1vyh6kvRMVlq3DI0Q6IMsjJS+fqRxm5PIle/BDPn+MO0TFXArWN+0siGSwXhel47KC8Nn
Z0LGg0wO42tjL9hduZk4rcqEHzO3VL1d9bXl4eGa5xOC02honEzBOZ5DJ8EEP8Z7hJlehDlsg8aN
1tVLc1bhtnus08Oed3/BJaQKlrF5v2pv/Qi0CGcB2Rm/RxICnTb06y+llruj7nnp+eJl+CE17FR8
bbAQU5cz6VHOE/pSEXZgILPdZfF8aXToEO8KoSBsI+eho57lpdFKedvb4LlXXeQvtaMuNSY6ff7Z
5KMxPqFjbrLS4VLhVSkNQjpLF5bDfnkmwBuf3QFVSnYKvM7cgbtnp54FEbaGkzs7JRHuIQmxTy6c
qSQ5QucgHIkjd7EK/5GNTRpAXbdCjR3KpWxwk4+Odi5Z/MTBPJ0j1GqcYJQdlqCuV8sXLSXZXnWY
61EiBN1KIGvaKqeW8LWPmcK/MfF6O6Bt1M/QVanBDhSwee6YAAmlhQeAKWOHGbm65NiFtqHCj/Re
SKv1WfcVVKtftLObPfRE/2E4WMFKbb7hjClquN2bG2IfNLXDrNvpBeXXASX4ps7i+Q6cFw+8EdoG
vGXd46IN2UTP+98OIWZ7oT8wSQ0zRihx9PesSPmt8kwzUGlWl5aweO2XFAGmFciuxd2zkzqqjUdg
dAuWEZF12ZVyDavYMa0rAtGRDG8nGIpOkmQpD9aS4UcZU4KQ4z5xhOIGOHphub2PhmitB/cabZv3
wJxT0ENU58nS3v8wnFfo7N/a9grOGhuFbRKZ0AScI5xHS51mwl6RqWjULMJGStf4jA5p2LRC5sFy
O7wmdcDznf2yn2TxFfXXBkAsDuBeby6y8+nROCfqOeZ11Rys7SwUISISEDvcMi/j65+kyNiJVIlC
NyZxVG7JJy4V1bqFblIpUfzEcjd4vk0+UKyuc3Us9QTvlOoNnENK/ycyFA3d7V3jzVKYauZPIn26
VPMMoCWNM1KLsJue57N2RAkvBnxA0Rp2d3500C/bRrXpVWF4tn4KoQOAyQVMvi5r9yPn04RKSyEm
LzN8VhLs4yhhCLRw3egD18OtiETLQ0+uWXa7G46f1hmyizuiJSv2z154HDcCIob3MYdoLu3OOgTM
BRit9lt4yY0RdjnKw8zhKStBE2IC/w4THcoktfuWhXHK5WTYdsOSklzsJlHayHIPsFBw58aepyjr
Ixmup4nA65iIJ3S7ZVyRry05R0bt8pRZaa742+zPf2XCOjM5C6nh2pUD1x0XeDZ/3RkUBfB3YtdM
c8GEIgERJb4QVpO/5vTCSM2WJL1kNn5g1+eh3xdDP8z2OfglGEibw7gui8PGxu9PTosRgsDDrjRj
/wvsOM58loc0HvUVsjQhdmY0N7awKEtjl12ZGml/leNmbr2u1rOhDXnCljflAm1c0ACW5KI7kNWY
mOcOV/10A/kj7WPSe1oApSrFWkHJiKry4X2AyHBPlG0i/1nf58lzauREi0wesHakPWyx4rXny9Ll
y2ifbr5tMwGQU58ZHbyGI4Zpx0KHTQ/Ips/SofEhPsTQHf3vjojl9rz/2tblTCJBel/yveHyAmv/
rAxLcKCHh24yAUmx6xgLgmz5AcjGW+UXXgcvNMeZPf/YiMkNiZmxN1YHcP56s57LMBuCiNNKr/Fq
6XK0GMgR8/NpUV+VliVpX9PGa6EfdW8shOiq3a79TMeRpzHsat10nH7QtfEnlwQxb2GHoJgKBeRz
fKN4r5SLirgohRvWynHTP1dQ9Zuqu0yJ95CxbVQm3p55QcTp+AVef2vC67JZGzSXb1lbFdY0HNkn
Q5I/MmLliGdBTbIKTQ6AOshtreK/An6ki21PvQZRLLZjy3A7UrRHj6wSYEEOPH1EBvgv+Ru1HUzU
fqIMq9bGrGXgOnw2GxHC63f7RQBromrRnXf4ukY98EsGftFeE0ZLlOPPRv9BECbwYvOP1RNWW1K3
wSPGUc6U1zJymHBDQ3ChUji90maBAgjUskRbS7W0zn2/0YxB8+LHI1bMpaopWk/p+bUm8pZyiZna
Hs1Da8cgZMfrwv8YiFY6hg/zwPlva92C0F3fr/TIZVzgcxYTFHA0KKjt2SsNY+lSjwJIdrERoBYD
3Se8WUBuuRpH6iSxxfCfMLjodF4mPiftMYe7UP/pSJyNr8STimroR8IxA4HJ55iu5zXA5KyJ/PYk
grl2IG21g2atdSV3zh46JpRcbQC8U/VWXCEeemnosUpeZt17RgtQ6K6rjt44Ppj81c/NUWf4fRFl
FLn86g2HS8yu2juEvM5Qzg8cSS/JTAcdlPxpzUezs3JtpubSbVmcCMyCRadQmeCC9hN3fE3DRSMC
H13GfdWrMdlTQIlyfV4jYWkwgpeVGjrp/7zb+8XHipsvgrDwXnRgYazO2VlBLXxsuMtt+oZXoN6M
DIDH01sfKP6BB3q9mJN8nQizmBLOie/wf64MUHiD4EtWUsZka1h0L9aC8yZn9Aaq/5hFXYijXZRA
qggvWEsyU4RIxAsfW9Xikt94CNGdg2AuWRxgNXA1+LJr32ztzIKi9to6gN9Ew/QX6PnoOYTajDFv
DSKwCgCce/ctYiv3QcC7xGIQZ2Usk8RPNjOkfulWT9VnChvXUzxawJWZeo2GKY1fw6W8Qg8fLVAD
JmiKugkFyDowv+y5uzWAojzo9SlM98pRR+gHOZ+Rfgi+9qv0kKy2OjCq4KvQycOMz/aN89HeHJq6
e4pBO43xkHXwHDpWCe1ZaYbzhKVTdzf4qaaCt6sIgtEDNKrDr8mHjM9Uq/3bjmOBuaNVu7uO1n3Q
Gf/pnnNx6TSjsrPJop4u8YjDQTvpBino8DVG2fcHhW8XVTHeMPSqQ7h9vD3Ihh4Y722r+wYoFlDe
3AqIHAeCWHcxjhxghUrBje6AGfqJBguqfgJKnYGbU/bhQoaVIDycD6ubCXIsTQON9B4rj7m5WX6p
6y6nNhsSkVGWnvbDEQbFu2sRmYOPCmfoNCcNOlyKeCUruBxqKsAw5sNIRK9Stp4xf0aJeiHIJdFb
A7mv5u+0Fq4PoiDog6s2YmaKUB0a94+g86DYPyqWjiI9eReDH0K5wdyscZPE6yYwO2or4hy1Nc/H
aj3C2rrmcmFB7BKAl1bBwUtQKVuqoi/0llm2JyWqq/j68Nvq/NxLqkdDnWVDrIzjMavxH0+U76+o
AyXxulDf5RNaEg++5FkgqEdJIgvln1JyS2CM3RfaAtDmLjIVlxQtOFIbPLLVuqGZYikoILFiG3ym
hfKJyaa3WVPEz7jvWyZ8Y82B3erSrgRf+BZ8f8sKIiEfl4qeeu62NQ0WHTW3aX8TDMGHO0phwSNP
paJOUITbK70sRcs9WrScW5CUlirDjdf4gD8K88qSDQwwRmCKKvIHG0RD5wvLOudHA93CeDw38Sz/
nr0F+F9iNXgMFayVmaIe4X6/dgsY4GQdE0jbeSy6m5yXV1N8InIUjWqfUFqCcLwxM+O1KEnDjh+5
4pnggZdRRb38R1ZsVE+xMbQ0r41KMl6r8uLeXG/i7aWQ3sicztTJzKEQ+P77k0gW6NixOTL9oApu
C7v0XhFvK7n3lIqctUlRJ5PFcbbJSH/pBQHXT7I7aFy8jTsUR6hylU883ZIoONxSxw6oQHJqukX7
j5va7fW14nspV1bSjkZjzdbzmWlhetISBsT+UjoBv076AfsbfQCAvvrkT80c289z6VxzZ+dvVV4C
uVFQCwX9dR5r3xOn9BuaULOG+CztBQrYDbL6s7BP7X8FFEc6tncLNUq/YHqJOvIyS0DHEgQM4wGZ
94c8gJjC3GmUfII4kMSTnNwCzp1pRvFFt86CCcjoFzoK9477Kd71TMTFtpkjxywCw5uzMAUDTHqb
9I8seeHzmqEbJH4u+vGkKc5Ch8S/Cy6NTvxJq+E5ZGPjC0qcdi39f8Mes3rUqyvSsT0y6cOZrR/2
SRh0DRXMz7pR+RJ8+D/F9Y5iyV0VSSvvY/kVhTYWYaIKdsmsFqXeoInZG5ErJiuVfLRN1tQw2vN6
COSNTJyDCAi4DWd4aSDHZCZ4HKQNim3yGfjODKAyr4DnhgLOKDQmwcy0RARMHHO+jUbhCh94W6Bn
Axk9uuY7Fr1E8GZB3yJhW5axSqCocVqr5IqcVznyWrAh3d/eO9s3VgAC4z8zR5FMx/mhTnOKyl3H
+ZsMfydmrAbXxAF4rn4s3E1BHhHo74N0NAVLBEr4glustHKt8NQhT0Pn5ju0jBHYX3Y+xXMXt5e3
FFWmWHVMbT8ctvTsxEvm9Z+ABeZDyY/as10XcYHkL2cEUgOuVj6I1WBtr1M2It9vIXNxExZCL6LE
3nR+GC0r4VSrsut/CTAVLjs9oUcrb6kJFjhdj5NHhOdEwKhLuuuDQmEhWQDPr10nLCCCuoh2aA2C
3wfACgDIIIWss27cjHeV5gBToK84c0Hm2qTIjDarJ+xGuT/gIRxy0nkZvBtwA4/HfL90OIt35Tb8
X398zGsckppskIcXgro++ZAO71AzuKe8oAMMtoT9d/FbojjYlVj+9dwwwuliEAc2f8MGcL4/FviV
IpIjNIYIm3nmS5CB7ewRpxLSlANCMRsYIADY05sKocjapB53DhIckj6272hKJ5nza/1TL4l9w1sX
B+uQZ+jaGm5W8gK+7NXZVXtAAvSjE0tTav/gQBie/PZFA88iCG+ywcANf6EVLmYicsXfMHKnVmJ9
K5FKTksxjUIcCjntiwv+3wx4IC6k1Mtt7QpvpVk0Ef+8dpISi/meRLgMa6WJAwWrr/ZfQFpj9SOL
2VfQPXzB0jFStUMQUSvwWrG59DLkNTN1n1C3bAmP2oabqQARxa1+YQh4xPeZytEPexQbH33aRydZ
S57Vr9intHM7O1nDkDkXdbQ9qoBNeWNCnmBnsdi9bpjvYPjX3PijkBHj+hNnUlFmLmoz+U2mqFTU
cvxuXSXBkB3leTb5TS1XWfqBQwBFO+X5UWfU75xpBBrWlwtZ2DZj+qgiA3QD9QFG09H1YKuODS2X
5rimqQnFp3s83399FH4gL/Axxz6dRqPqM03EMlyB+sbDlY4Q+WSKk5+rugtTyctHVLcJZDSNTv5E
UTHT7y1lZlujID0RGhZXKtLXySWmOtEhuX3sQ9VutrYYL+suZVt9qBoJnPcLj5/4myf7Z4QkKQ8/
YBI/Dfd/k/rfjdrvvpvmuHuhOdXlSS6RdBYXS1RlS0npxFt+oMDSYqgJRLZ/H82sSqKotg3L75EZ
+OS+Dcm6P3w3SCRgyzv5/XvrW6EC7NThYY3F5yDRepgYXr87L9qA3Kio9Ggg1YuGLC2/BkLVxq1+
WBTNpJJaKOwyK6GOoiDhuyY8Te/lAY/XUDayp3QjOw+otz4sBAam5SAx4BtcEC9KGTEep54F0wUk
b6gF5iF7+2OIxYx758hRST2HDqsIh1fVw+vTVkT9aRkoCz5b4nB46bv+WICBImjtsWhdqIeiAeVR
XXRVEs2Q3f232Rw2Xon88IElZR1TimRMdn11GgXg4zGh5v97qNePcE94fePwqvjt5icX7H1JmY2b
GJ+4aA3lTnJTs98n68LoBwc5JriAMtSRWnpr7/e6/2zr5L6ooBWLzBo6PhlKp9kxPOCUvZrmC3jV
Srp3G6DxjCGA5IJdUuUxPZ+98yq9Lt6RN77KiNDkQPtN57tLF5/ZEfOXYKRrXc2IokJHOv1xsXyk
ipLe06PHUl+CnG6CDUVsgpc2MsqIZqCRPWlAIfO6IVrDRBNcCAfYtW7C3Tvnno/s2h3mqO4PN62d
/ebhsbbMo9Z9m64QwwicHZrkkqiJLQsqjhzWNIQV3rRihq6iQibF0BefB0g9lp3mDDuhD+O3r/te
lrWuLvg5/dzMTCWT66ZsggYNzDze5gCKwZX32mLwnWdB8v9ZJywoquDtmxvKx3fZO/I0BDOdPJ+7
0McmLk5VxHs9p1ZkHDb+zqpMJMteUER66SA3wMVIcRfQWSuP50q9VYJERxf/g8+yihxZpl4uuADN
hlr2dh5VGrY9z80SRKZRyWTVSv6yb2lugIWXLqxtkwY++jx/QnINeLO7wTTtdZbvlmCoonGSEmCN
Tx2nfjz6mkTyQC3MYWiPeeoEEA26z+s+e4ZR9bICYT2zM3gqwEYasGOTAmOAzPF9C1MAcWFygZ1Z
HzYTwCVtspZRGV4porIesCrRXNMb+ZjVqyUI2+q5eeFRIEA1zknjM0Atm3czIhrzaLShXTBgR4se
79BdxDJq98g4kKIy/PjQMuBxQyncRjgQODk5/PraYQFw5VEek6Dw3TJgH/wRhkvrxHmyZQHEjOJ1
dMYtwdxsbjK+PAIr6anfAJtFgsj6eh5kCGVxa7+9V7CUSrAQFVVykJrpmfLrOKS9jGryuk2a9Ji1
f3jXu0z+E6S2F4boUxQWDXOk9aLn+Civg/S0N6pRirOCerZsJWNOL20nR8WHqW5NxKD5ndAFXXwt
1LHOC06U10qHOLpmUfvQ9dbHMFlGpj0uEUuSDEBTCLFQQsZJ0nAwJTTUQE0OkHgDRoo6TISwhRag
uVMue30n55+GR0ws4nrf/tbrQ94RyBwexwZYkmk0jkiixos0vu4dbqXv2xX2KCgWoXRG+Qllng6j
UloRlwWrJSVMbR+jaoX6qWzs7FTalLoTkJANYeSrQ97xEU/cjOwTZKlSxrOVDaTntNvV38DSPVmh
1fDOFdRzyIBXr3f4053N19MYpDFT9qjXtk1J++fM4p9p4iKLi4HDDNWKqsC3SvZWPIIF+muk8D8c
OW6F8SCksBTZHur+sbs14O+cG0oXPRog0ws4zlL1VKQ3MZCITOSv+GL2PWfJoEw/WuloTzlpnECB
6i/7tgS4IBxl71INm3wyeyPdJV9FEDiHVvDYeDVObzDchoSqNVrXUOsz4VGTpEQACjYyINdyy6Qp
AWdN3334Ms27hvhjHN+3Y3XOLkptD/JXlQZqAP9q4AChjp+7N1Ec7t5ZsX6SYkRDCoNexZzIEjb2
tbUcbK2Fumg8z+3r0hq7BFZ0bvpFre1cc68wvY8F6DTUN1iXzLZlu6rI4QLnVPY9653OzBpPukcl
wEOz5YqPDY1mhu6Q9neZu3oE1bC2RDQnT8AQhYFQ1UlwxEM+ffLs52XWqDTiKNRrZwapsWiDfSbF
4Vr5D+r9CpzoJnp441ZmCRkBrdMzUSB320c4nGhfgGOE6DDehR1BKHKjvv3xU3ruOfxFo6v78ptA
MqDxr429/NhR/g0qfsZTJdu6SpJJUZ5ZW0bVJ0Mli6a/zeKyd5Jw932qL7NDt0pbrNz/FNwkh+QQ
0Cjy+xDb3vs55uTBoagwgVDuSuRzY56Js/Lexo8bUkUeqQuo0Vr4aE6TQFRBQEno7kzPAb5J4d8M
jn0tXWdASyejQ3Vh1l11r8qedVg4GY9ummw2RqLWILvt3b2Q5ML+lvLtyuxsGHMfQ49AL8ZZ3nCL
EyNEkqyW6cmTU3ruT4OYqRnn0RnFquCdCScI1HDdfpigBMBDVtVjLxEIoOO9q5sSx80/yL7u9ehD
dg2+MeIgB3wNiFFDf/PovO8yRqI31MHkaZUjOi1fHmmjLOszKaqeMjGT9NwXqXn/LmyGpLdbLQs9
Ip1h7S3TfDkmhIOaYOEdGUuV308Tp1uxHmEwTyUYu4/y4IZRfTCW4RC4VzLrPnKjrhrhTlDtDXua
3oKDWx1ThNT/YSNbHjEe5XIeYNJtOMXMGFF88IQbJ/nw4yjNSqZWCf9lwQhefeuk+VUUV9I5/2I0
UVro07uwMGWPczO1WL1kxSHlFtfULhFxFF9BxYgMeRSBF3R3fMDgX//cxY5iZ4T9zQCnKOewxeVF
e+Cd3d3VKxWS8zGM7riXpryowU39Uyh2dQYqcCqGSeu5RomxLjPtPMBnI7qSVV2G3qCnrrJ9379N
aO0/GScCUBSy3HKgIszUBv97lcYUvtXcU06g7Ys2ir/4AwrM3iYAy+KPn5FnDZk5L+ffKhw7rjWE
yYWcdeyXlzEBJeAOJqx6jd08CG20loOU3+AhhyfbWcviP1Efsdx2efeY94BlF5DiO1OKm0IeSQPv
m75OBXX0HX+iE5Pt0qcz0MNffO0DWyDBeWv033RKicKCTBut/skzBLjNGDm4r3k9HWaekoBxU0Dx
FOXZF1XhGBGkQRjlrUrRgFwBT/KnIkrqego72Y030ikZsQRFS9ug6WDko7OnDNREsm2GyLF86T4j
0A5QPbt4UDuZlsP1GGlpydIO0t8ME9o2zH3lcVCvPtjKrpEf59q/VXkK7W3/GWj/736f77OfA9AD
e8o57pvqVkkzlVZej9Z5JDdP5lEcf1u9pwKBnsXeBWkkX0cN3g7BgHDgOVhhLDBfXgzpU4TcnVGa
3xjtSWYL5+2hP7kALkdJbpl7N1wPjgkHC6RgWfAU3d2RJe3FV5AspXTweLl24I0mg5J1bkUS6htI
kdRNx1KvWIGAhm2jnm1j0UI4QA4XQNmUiFL+c8X+bum0Co/xC4U30ojvOeLMCowl1jKUoIbxCjoL
U3jRwrCaqTGeKOaLGvEOTY4zmvNdz8GjW0ddzCeqhmY3JieJ+hFRXP5R45H7ST1MkJCD9yKK66O8
Pa7EIPjmR1nxKpChEQIlZgRlCn4GIYEQJDrKooR77QWdwMKoO1avnGvDiUu/+4ZWrHHvy1tBBAWm
ssXqiuE6uLU/Bng5VBvsFupsuKur/KNakoxDu8SIm/JYx5UNKjViuMOc+A539Wd15mU4GKBihR2D
x+NYT5gvmk6I9v5cEonmWHrpehMnRswUpCla6QTp6DoG+fQdipXntrntYb0kpMd4XPPDJaKDz66g
xW5OTTlR/awvKQRR9Ji9IICg9TzHr5nSJxofKUsk4wcVaLFb/568EL7Rmori9QVY4mlhj4GI5Tlk
FItwXh4vxWe+chvbeWVxuUPHCCzprdgrwS22AUzphSBmnIMxJc++lzMeAEi+51svoG1qWvJoBtIP
pRstXKS3LpUiBLGp0/gMMqyYEt3Aru6rJ5sfN7XB0PKg+p5YvB02gXk32JTBNOc1b+QwWpk6OqzM
UA8Tg669KBzGB/w5tbOIjczb5lLCsfgFs6pvFAScI03zBDLyE9zzxqPYyobKlxvhAp3xSDqOD0Tg
4kxq/1B426dyzvT0NalJ7xEix8yL3ZyBzH0O6bNNn9itZ7Ed6j0NXm4JCTkdfjVQLwSZzrdgbRcM
omQ9HPzmuWkVgBfjEV2THugdvG9RNnm7KUgKfpoW4RuU3ZNkdsSee8eabGcWqrxL1o02zUtagYJj
Dja1mRFckr26ECtDUIu23hT6aI5XFVxGB6hgnJr1I8hdd8obVfSUyyDs2lfrji/D6Eog7bHGgCMl
R2KX02m4dor2bRPQYs8TbFFtLYViL7Kh9VWSwhw9cRtW5vJIzte5AD9lp7CQtW9vlr/MZuxIztVB
ZDJU6fnk+LZrKDJXQ7byq/QAg8mJji8npA045NCOaczfuGwYeMIg41doiyBR96YD0ty3dx8kZQBd
xw65Q0+qPcAjlY9BVXPECsYOnOUk++WhDFpUbPd8ETtsTmw/Zy6+zvSAItC+ESLPYbp/L4RyGZjZ
rjr/CneMPniSUK0ehmqRyAsfQS4ElcnsIOcWe09xzfSWzOiQa7SW0wVY1ToDK33KE+uxJMbMeSo0
vcqwBdXIESi+5vrX3gYPfmyuGRxzwsp9LIfVzBrlj0dMyd1yHYnnMssjjhOcX09wKd3ThDAreivG
ITvbGFh6UktMP/Odisf1edxTT3NXrcVZcEQw2eV1QjK14/L6n+NVXKcZT4qovCplJ/wXSa52wyjX
ROj2bs6yPDT2lJL7WHwxYvs7GWMNUvO6rFotAW47y2je6YhnFNnw3RG9MG8KhZwV8GT8F844pIdr
IzNohMfG5d3Vf5hxxnUG47cRIlyyPCB9Ci8YB6rdB35h7EwBMTTY/gUxkX7MKGG6cYHM8qqZq2O0
aSbF/S4AL/tZ45CBcpxo5k+Xs4XkvVk1se0Wesws6ibGogvuU7CBxWwEtXaryw7Cn42mJz+TZU90
rSwypIqWQUltClYqLnmku8rmr6GQ5Kh6oTlkaO53OU4blF3mzsK6N+bn4vke7WBXaWrPnbbL8OuP
Xim6A77bQSdgqG20ENBmsgZbPI47LJg/2R0CYbqhoXVPprRwgnALvbL8pwI8NBpDpNyCd4PYZ8QP
fJShQ2OdIDFj6FxxKvHPxUhG3mvcU7CKunlHHorNHh2J/2CrIVi3jjJuSOT+q6roXy4GaggnwjyN
Yamf71S/VE5qHEBGv6WC7acA+SJcO6DTS7bNx5UQX85oZKn9wgWnBATIBhE3ZzqDabmyB/3uYuxa
4/oGVnMy+TCzd7BN1UI+mrG8C1c5nyGOeoTzTyDrfaP9W1sUyG2TqaFPUQhDf70N9ffRaddxfNr7
BPJOj8+8Fa7AblR21w8+l6F1L1Rq0MV4ZSwMX+keyGn3yci9ERs+1Y/r8nSCnJTeEvLxkWtQrkOv
1IOM4f63dayaArD52mB1Wxo+20LcvVbDoLCQpfJTiCLxu4d92PxGPU+JWauMDcvfsGMAOKV9E00l
DFbFwCYwGE5gmb4usktwBiJ/vFuNHkLrcVIC13F3mcwcCgsDJ+nLfMDrYmBA3F8jE0ZDkrHvWOQh
dJ+LtZXvYLsd9AQRWSkbMPoZDutx+qWm59RKtwdenIT/xe1tGXgbMRVSzxAUO1cchhzrRcDjPmoQ
MHBJtV1wRxw/zTQQZmWaCRxwxmgQoNhABQzuMK7ZzTalqTBU3MzUfTow42OXJqukAbd4p4UYSrg3
revwuukT2EFQx+hWCV5ia/reY4QjuplNtKT5AIOs9BoDgiqmzuuhjvimP7D97LXQksRcADCwnFRL
EThGnlStpTvY50qDXB4rgy2bAMzFs8IMtxCQUAbMMTNcs0g2ZTkrXrXrb4x+fh5TXJNw6i+iGLKj
+L6R/evWNKS+u1otu8IXIKJz00J/GJlzbj/JsdoUwI03MevQPiIsk1qJnnGkSmliCKF6SBpcA+RC
k1/LEjTxbaEw4mty02yfvJzgUkz3ekj9z2TyergcYXpaYPcAp3sohuz0PNMqZ5tAsG5yjMOFxDRI
nwBnoMPrQQJ5ZCW8/NpImRaEPQMwjND06fyzyof9M5zMtQhzr2luQSDfjsQiYydP5GLic4fII7q/
983w2N5bby2xH+R/btfZRozF+31isEn+9XkGNXytGrjLu/ITWw/OC5m4NGa6Qq9XVvcjgEb+E+KX
PeZXlM5xcur0Sj2jgCYAdOBe+SBvN4+a69RXaySXlZkCMHlWXY3c3Xf8poJeodg4XC8bFlA7aMQE
PWF8aylDcnT+Du2JmdN+0qI9/HrTC8xH6fx2ssg7yomyEwQM6UgygwO1RqQ6WjigHGXMpg55XcWo
li0ibXMDAkJBek4nGxsC+inOvB5fWlXR7OqvS0WFYZypwQbeNVM91sfESAf2zZxd1CRjmZnJjef4
68X38B4jc2qn/2u451t5I1DyjK5bBwdSjmSxoUoYSRTMJ2GWo0ZFh+xokUzBKG62tDMAger6kvBI
PXc5oQRVLkN/gVCX3yMPfgiasB2crfCq3PxwdzziqXqqxv2SYa+0PJs/1Xfvu6zCKVS4h/o7UCo9
8SN0Q4RSaYLvnAZ79JCnQyVYhzGpQUHtqYLBUj/jamcG6XfRs5N1+ZDqdBJMcIp3SRkFNDthBClG
kBMQ4rC7IWuOGNy9//jy/2/vR9WnnWebS5YK3SXVUaNCodOjCpjZRfMYvqmjAUB08qW1bCyCD7mE
p5bz0KKfuLrC+5DGNO818spVgJZnb7PTRB/7e+rYmxDUAnlyy2sSP3fqzZKazj14JLRfxiELwhz5
mP2AJrJeK+q9jSsz/e2EVgtzGxca/yflgEF1nKPtGm/cdvLa5z8ZwCzLb53wsGAEhfMc7kPo5Dt0
4UXYI9GowElPE0E8tPw+ra9s4GDPOWtAMsKdH3WEB5GSlcGdZLpfkrSZH7+NBKICuMz6U+LyZRR4
ooog0zfyCn1OqU8N3ux37r42GyWtZbfGei5potX1ESBZT2Zrbqwxoxqikw/8bV1TLJLTHe9+/lit
mDIk6W29jsDWHBPtityA3uTxyAwbYDeTgYQ8Ke+QlC+WKD7WpjROpYvcTrTwhixmfvBZWm7LMCoN
FebY9p4xY/kCzGGdlepfZjdsAkq0+DEmh+Ouz3Lrjtu0uCocAAjvuojsKmd/oqvC92ybsCZXytb7
1GTBVPcPCNYXg372T8kBP3nUv0WXwodULScZ9A3lfmRAXOF/isFb12Yzsibg/+qb+06dixnbzKXL
2BYclzYg//Z9OHEGH7KvEo9fZ9bmTIm4HuilxMtM8XftoK0K+Nde6DNILbhqEry9ka4bfsGadfYH
N3uQ9p/pFJdw1RK0RF5P4h8bSftiLgdF61jrYhfKeBYXVXFOaY4AMgjx/F2a0Dh5I35LCha/Auul
Ci+mUXdrjW5sZ9gKNPOMnCdCpxiYlcBH1Ly6t8vi/CHJeB9pl1ag6KvyW4HJGR5u6OvXtfMVA/MP
1VcOuF/w7PCL4N4XY7yXYx4VB2u/XotmWfD/6DPYfsruGTRWIGtas9oxepUwVYfEiWoCKxC07hjs
cmzF/CIUJKSKJiccuKyCB32vyIOVGLFzbVdefvZrxpvOjOgmURjmwKhjdSOTuiXqRcL0TKJFMtow
jDA/B9Cmm/d0NQLYxrQG/dccF9Awo/M0M+4qHfqCcvsKqD8CimFWg0n3VoA1/vmmOMdoVxZ/4yn/
sCZQXRWZQ3UC5OWx9lLAtrKoIXJPqeQtEENsctL4r6AQR2+OQggLU6bFxsV5wtBB9BR8UswcpuUD
DQSt2p7Do6T1c2OnEz2TAP2bKxFlWRy+uFpNZ5/nQg+4NW1EBIqMHAjHFNKtxRb7sBETEtTCAR73
zTheYH6AKKN4/EX/l5dhxqEc7WUqnjUTd7QeulBo1fF7QNLmT0MBMsVJZl5KeqmncPpbsZ/7/Z25
4m5qqlTEPxsGg1XFFwbUtaSUhXue2ozOzlTIaqVrT7faMc8ZyNX1WAuB7zhlzZnAo72uaWXDqd0J
BlN1HaVqRR0cGOPO7vOAdj+HjL3UAPlIVhTCJ9LSDB4v42mlbH0vjvFolyPltJ0oxseajdyoxsYI
U0Iz6ABfwOpJPvjZkSuoK4xwpcoklHgfoldIa4Ot7Ct9SThTKANKnQ9jCRQOzHmGzon10k3LsYD9
HSQf0X5tR+xAiidLylGgr2uQpyC7kZD6kUTbu29EeQGsWbOnUZjeCKWnFQ9tLhdeTFmBERfz+P9m
40kJNgr+3LyhdjNPifW+RLmrHt+/Ok+Y+HE3Du2+BBSMbYJc4V+A4JVzHWb+tgfT/3bw1skQkmyL
Bi6YjtfC2nhlMEexSqR5nyR5mqlZFq3WhH1Tx8cvfuJaLW5hXl14NZnZJjgz8tATJhCcROqs/F2W
/lNMPz95vsasIEgY7RYa23cOUEqF7UwXAU7pF6GbPZn5GzENz3PqZgowl3W5xICUs0wQO2vdkwgs
SkugMckrpLY5SL1cnIy4klJAs3gj7U7yun6AzvP5WeNnS32nLTXuhk4Q5E1/e06yTvOFviV0UOFr
yU0uBaYZN+tu8sMjCWHCDIxWin4AmPAz/lGOVTDd4A9kt6MuG32e7iedGIIlDwOYnaVKtb0btAzl
n9O7D7h4nLJ3aCXFbb86PXQHVCaFPEJaoSgGv2qRLEyUNQVEhdrs1zyIt/EJ6ROAF1RowAXL43Aj
EjUCYId/MCdHT4xHfvOTIm0ZHrY2wKcdlXe+IG69GVeVVSKoVMeRC3HVcdRP8FPmBlNK5NHoMPQN
FmiuatmQBhsfxyW7GwOaM8fPCe52tTS23cRqUbYA4V28PzCfuU3Ufvn6MFso+JKBwJjkY8whUMyo
i8TuSHPTqRsYj68zI9MJuJhP03td1Hw3fSMpGDQxxwBJ08XAs0GBxj94XiONS/2H81gRvqgk7Iig
mz3woIpOjKubADmmrBi4eRc9Kvj/E1GImpqPs0PaFDldexhHEYk5uwZhn9vhwRstcmTXuUALawa5
AXp12FXASNfy2VFcav/S8fwN6lG9IHd8YiwO1BsDVJPFH4acd2t2nHukVvUNoREWPtPTOIFDc+ht
2qIwanXXL7OK0laNEkK/Dd/Y6hU00ocAixlZp8FEHICElMQp6pd59SlGUQ6/yMs6ZxfFV/8pfvN3
oIR1DLvOgMZloxeRontR7rhiaKCFKWeCj0Y9/W7dbdE6YEJfzoM3S25iJw5tH5eGUkdq4TqWESPE
EF7y6eUWv3taj/Mm+tNIPy4oTgyuZaML8bspukhGqHmtL8rLAGms5twHkWBfYAOa9hKKLAZ933N5
rY5ssNmvhvdpZy1EMEfSGVBYcLWRDxodsRtuWNEIWu+sRIhRoC1q9Z86lmsKT7RHM1HAqwIdumAl
19kxZuJi/R4L7mOr7dK8UCU5dNYI335wIdafss9XYzxOVeGWiYdpMexAHTe3616skp8U4Np+OwNc
p0UlvpdlIE9rvpwlToIblnc0m7uW4pQkzYf9giixo3NqtY4e75jb9fhZok9G5RQTBfcT4Jlm1n+1
mewmXgw3Omtm8qeQUACFipcw2ubtsWdBe7Hh3431e2SC3F7uvcFQnPAMFibC4RONg+hKSyak7o2U
p9fp7utGo2g+qaLdOI4R4iOuwpioz2PB+YXbRfTNcJQ6630sZlwvXD0qpKvLCxle9KooQaK2JRNG
1zZ7T0TGVl7FHJ21BjL9bJ7NxBLIlb3osEmDC9uLcg9H0gHh/Z1XfmjdPuPfyCPpZg64IGGgatWr
4LBARWdI76KphHaUI9mEYBQ/S10majjgArddXRQSFiLyglXLTmBBx0zxdtZ6uPv34F44IXAknvL+
ruArcO91JFH0qwFkdgVi8G9KK93nmfu/P66kIzxM4JcDOBL2ORcA1i86nwg9uZEfcq3rBD5xOEus
CiQHxi8TLLpmg8HsI/Fio0wpTB7u3adwS7lWWTzpdy6sr8uTCVAe3p4H9CsVSrtbCL8Ir7Tv6z5P
MBUpST4Qz9oqD5YP2jvh0C9/IgZKK2uxFMlQA8GHb76pTdA7WAQobqwNLTPfOCgIlhEc7uVhJdw0
wlCcpAn8j/Sqv/LjmRf0Xs5G4x3ki764qqkNJT4XCYoQunNxgo+cb+sDhjhIzYGcd3YrSX3duFkA
abmqkkX8zVoOw63yg4uhdCXyiEZ8QNAAOvNcNED/LVYenQ/fzLe+Gx03xcFXLeYGtwIGIsK7J0h8
CSqfDDCUk3ocw8/y9e+9WA6CHhxbkRjUmfKi3yRtgZi4jc1FrVuSFw3K6EwoHx7IDA4+OzddOSQ1
NCJ2yGUNgb1c5NA589/Tzh63PaTtilEkZzYkk2rIW1EVoVWW0OkG3tcCQsVSecEWqo7Yrtb/xK6M
2jv6Q1/pGgbD9lFGw6lKKbscmuZ1V9OLXPLefa3Od6ff2ErLocamx0Pke24xcmbP2JRrpZ29uuaU
1tW6exXWdtut851DVCJ5RfENJGO4SrCpbOTBTRFIJ9BD1YwQZ5u5hcBdltT18lPbxPRBCpfXd25/
YJ4gQNpaVtk31qAoLWGclBj0tLluqX3iDLzoMl0FPLqg2qRYZr2Yewx65tUfDCh7gTSJmF9ziXhG
rwjREABr6UlSpsAgtbCTe5dOYptwJxR7AIws2FPIT9NdiwWVDOoNXUdBayerLLlayHS+4NvT55Rt
6rNS7MxF0K4UyNbR9lkFUKfcSS5Z1IzKLXc9u+F/+4Z76ruJ8eSBouGVI3HvKUPoqCc/pWCF/kz9
rYAUH1PW073BiAFBkrwJlXUO/Bw89Lne/IwmwTMWw4umD4B1Dzh+9PfHo1b20IL15R+qg/CY+HhE
WnoGVdONvSJRyKC03354gDgGNoC+HFR3/aw9/hVhI5mb7lAk9+s4B6U7aXnWZYKWcy6EJPy2q7sS
zrRhWOGPEkxKCUGXSXDDxOXcVLlsTa880xEipGtkBN9UNvqOUb8UKoklCXVslDCRQZ5r99xELaCQ
f+Zg6R1it4FgyypOp28GyntUQYoUaHV0GVGs/NTNdTAWj8X8ESpcfqjxDSPHWpOYKow/+0wFpFnu
fLQu7qxEZfAqjQ9/nDvM84JnF8pwEYvecwOOP22LSz9/oVOapSrEvHnjMzDD2R3F6cfGG50dhQWc
W/yO0cC6J53QqVJIAxCJMXDmJ20KY/AA3Zgk8BW7v2CCM+jbnXx93AknfG59Bgnv8OoobnVlqTKi
vBhaOHGRr9QY4UuLIbSV6O3Y3yF21tUr41Ew9bPbM0hSJ8cBnqqSpb7091uEHfCmbVkSpTYpK1bE
GvWnwfqL7zKFUSkmDmWuuHI9xRYhFL2Alc1HEOnknHhMq7V+AM/ciZQCsBp/p8cly+TEhnil0gt8
30qWSfnngl4uXvrllYEASNtEMKJ6TYxNM7YMfYyOPtpAmaafC7fp1EKYqM0HxRUnIcDaRU0vNNOQ
sXLeoIchf+rvIZB1/KQN40KEgsIlQCFEy7emjm90qa/olaYzhY4R7pMxiTZlmrAlSuRSzs2+H/6Y
VXfwTcnD+xPNQ5wJeSUtC0W8QWMVfphLL5nYc6emWt5s7wk53ZKdfYV0fZl60On3RdKUvG2r61bQ
CEZbgZvJ0ZVfycvniY8YXiVoYpOPaFuQq5bDGYuUAkOYpSj87Q8t/GFqLqCB+M66DIfuVJD/wGWO
UtSYTB3vWBCgYHBXF7BfCXn+tJviJnegChxXIgpWWAapfpsvVTDAxzucMACNolGmqO3K2zVS2/eg
C02jqsybHHg38wLM7NItDAPzLzbsQf5AKp/HoX3frmZ8tpRqTshlMsADyupvc/AfWY76+fGpqc3c
j/3S8jiRMBYBA5l6Q0sQGVRT6EXdX4qNY/U1sORYyOPd5L6m7Ir92F5+13XOCAoQJlbgH6mKhfYi
FcwGml9P0F85eXhoiVk9pO8uM+ms1VKHM5DQWdXHNYdm1kwFahW1WyQ/0VojGgK7t4nOy6gfoQlx
2TLUAzFS8tqE1czvxGZwntahsqJ7gtXg4VOy6oWPbbvUCv3Z5HnmmKUOoNuJPK56IOiFTNUegaXa
vOTi3sb+fLLT44tGNuI4uVAuT7EKJJQY0uYJuYiWZki9d5ryXjik9bjsvYBCefz0bf9/56WE+cAD
w+ReNi9xrKqWBEkWk4jQEcaP+w536NSIMFteZQXNJhCIOIbY9Q/kjAX6WxpjfPY3Rd8bCDDMKIcL
GnzO++vQu8EBIgwv9Q11lKUux+lSniAd6HMav4b2UjPnEFWUPGUoquzsXZ3KWE09wdBS6ewRQZOt
9W0SXuXeEm+6LkfLYlN7qXes8Pp4gjiT8E0A4w6WsP6GZR0JkgxrasAbJx4oMT0jVRyGEZsEPYrV
XC6NV/A82WeIHCRd29D1NSwBKqD13fvg9LHVxB9JIdWo8R0zQ3W9bTwYaPbCR5OtEhaM/EwNK2DY
tq5w58fWzVxpmwH6s99kk1c0BsbhgLwDc6oPW3VeaXZvSaVTgFRmyFlKhhYQeszDXH+HZQdJHpKg
zDGzIEDcLgZz77gcw/oEMzjWNk6b4RMjQv8o1GF4YcYDObxKwdAN5w7ttsHzJuPKDRSYgVYFtQFV
8shgrUC9xk7PEfWoANFV9ulrqlsVwfLb3bPlDCUAAPCJYd/y4heMBnrOXcGnG2hiNzqJHn2pF4hL
6fkNrt0l08KiubUdp9MGxsFDMviF+QNzb5udsVh0M0jZcF7u/6CJSWwxMjwMR8Ofpdpj5v5BoM/Q
TZIqE48GHsktLVPLFY+Z74T+DmwZIb3EpEdvVrjb4k6NkHj8huu7MrVuC6KvxOwZt95uIYHLZY9v
03KWYJIbxiezurknkpOzqHpktZ5wZ9kLS+l8uLxsguNdqZ+VaGGfj98jRWSRkFbfYFojpCNUCQkZ
KpDOIE2/6SS7JboEnm9gwvl4eUw73HLF1lJDD3HGNQaw/Q1IuENw654vKRpN3MKSWnQC7GSHjR6s
mxZiFEICrPShy8J4P2bE4l4dfCg8DSGs6D9rkxx249MIOrJLnzRTzDFz0hAYKkPDocgtX3edtecL
dWwUNL48jRQ9WuvJC6ABIFAUdF1MPYQ2ibUPziBOGFxQIF0/iZIzRwrHXiCjyfJQWq+FpNi6yolj
gRD2CtCAwlfS1sGaFuP4ux7Df+WMlBABrXoQH++nkAEZApyRTKEN743igu1QEWGWHb+N6FEpv0VW
VfXVA0eGcfi11nfbaNEyMnD5WWdGtLpZAsgUnDAi+niK8ijOtuTUlpF6+qtrbjbK/UdztqQGXPJN
00NBYk22cr3K77m4k2IHi35DR2VgpWCTqsGLOMdV/37dta0Xtdfs1Uz/bP+heAP0ZAvooVAu28xG
Aa1sxXmz/1hmXHN99E875ttJA/xkyMz7ckkEKd3UugG1zS7EVqJ7gS9dHBr2gn3sw8kDdWe7K0XT
500aK7PX2c8eklOZALhCe7cfh8Lhb0C+U/7ZEyWGXDiYcrEYMQrgjS6X4MMZtUj/U5dItGcKpsqE
3wh6/g8MSkmKmEec9cyq+MkwtYlZW3mKyWhgJ09ByDrVxmOVcd9dxX7NI3qifecpyhas76gLaT/W
khXgzpt6MMj6imKXoVDPCNoPtmG77PKzAFWU5KaBy820fA63uc/C2ECTdYQPuAUo+FoEnsrpTK2t
sOSJnYsnJbMcZLsqaN36xkN0ehGRx6ILYuRV/BLH+Q4GKRFic7uVCHeL3uxlgiBm0M6bm+muD+0J
qIKRJMpn+xJadXAclYD+6f8KeG2iOXZ7VI/Zvjzsr9GFdoPzAYjLg/pHl+EQU4glL/MvfoKeA3en
oMxmgsOdL4qyAJeEJWwH2NG21TB+B9EM/XQVZgUVbF4sDtGUU7I2e5GsTUnzzkPbT2ik1R5XrsYN
STUpaZwN4cHzi6PDCy5NeJxGS3XJxht5aphNP5TgF8hZ2YHsKCUAv5DXHVPlyWaG7lopWpXNmSnJ
q1GSv7qCIBOB8r9I3/zjUl3GAFoI8qkvo5woW+nqGlhnGuCvlsYUh4wMgu+K2YgH9GK98ezQWO3l
EDpjSBhExapRK9FACFRh46nXUqe+gjD6twcSMBneKRdwpgf5uDJuth7jyQiEZTMZ53owvs4L9Ehh
lseN5MXBgsUoBpTCt5TWicK2OGnphnS05BVDpUaPx3fblMk/WpIrSZw4DHQ+YZZx8g53aVVk6jUO
IhGUyN/61WqJBOcaZmSw5J1swrv9o07gypJQvTigoA+sn4+QHqreQr06rcdjIqNq8ZIRGwvlbNAl
wZQLRfPdHs21cAdBQRaBKphx7aQSoV9kngvrQXHf76IavTCowUxiQwJfsWjGfD7by4J3MEMNlnYO
wD+goyEFBXQSS2KkTPZ6s4j1CJqRg4gTBbkLZXxuhr174loxkt8A2BrF/iLXfuA8v4eim7ptWEFp
rPA/bh5pfNX90FpI2mk/48jvnUtVGnG6QaqUwQ1+N6k2WiKTEar1mlIvmOLykMrRNA9s7hFF0+/E
YwHGZUs4N8Tp214yts0/iK1TyYvGeEUlLt7aukHIn1NGUsO4U7YWIaFcm4Zx8gNu34QH3jH+n1nj
Nr4gaDbGvwWcqivmSkdUPtoIKP3s+k1EyWzn3UMqNybK8pD5qYPm4sv8b1+XS88EGKGywuQxvLM9
U/KFlUmDFFLHVQ9mSzJjl4QzUwVEnS4tVYKSSl0dbiI27V0t85ZJW8Bg4qtBaUBLx5L07zOXsv37
VCWPH36mYH3OWdki6fzOFsxGeerksRxzGL1D4sVavNh3xIedUd242BWLMJ1PlJ+VQQena6FiZKqI
jZ9Gek7YvtNifxzkGpmtniCunHmT042YUMLDxFpjBKzZ3XkAu+SeCGXlsKX0rLRkDWtDwkuiLvA8
tx8MocH8Inf8mThhXcaLwIY+mTwbaBrahsUzfV7ZE16I2ES0x0pljU9RLLORjMOjNN81Ml3W7UPE
kAInf7hfA3asRJCJ7mUywCUL2OKPG9ZBehtj+dvWI+MOzLtWnhztbRCxByEYiBb6thMGKS+XRv+0
HJp/8w9i5jfHcoTvXC4lwCc6/rRs+m4VVUlST3Bys/RB2SketKHj+QM51tPsHsZylSkIjKG6mBO+
Vhd4Kr80nNKv+xVrngf74nNldTCZLou30HMoBqNh8MJ6L/qX0BfBTH4PW+sqWYclOCWoRvvI4lmu
MsBGkDdXjKYxijGuGNpF76cz1oOboo1tvmwkfcHtXrbu8w+MYIxK8LI39kQbZHhZHUzym89cD/2z
PgqcqDBNfM5LHazHHPbPEHVvzm2/wO4MneAlc84xTmm6YRvRCLPs76Tv81QAMf8jnre+uXCwlZn7
PIIG9w3ptG3N0GlKJKfQUCpRHEsWj9iVWj7Rdqz8WX7sKNfFg+AWpFgm6A6TZpH9hAtF2KEe6pPP
NZ23LuU8qoZtYsG4ZLpNdVj/7dUMXexsGKqbBBAMWuWp92JD1bDk3n1bC6wnMvtHKQTBfMkLCCR9
ddaSiy8GpSmsDA311zpoAm7iaw0ABR5emVDlgNmm50oCbhh3+7wiDi/TiUG9AsDq3qvndS42csB+
4wkONy/hnbp2r0VmnoUQEMIiUCzcvS2r1xgE+laN9G4/A6Cm1KfsKSSZpFR/EK4vPTZrRrvNEGtR
J7XRq3T+gQS3F+hlBWA9PM9pXII+iGms4XEXNZlPJd9rD2QkRI6H3j2Z4pE7bPBGWpe/SvrW5lXd
ZV4zlVbqQJ3jFh3fQlOvJsV0cUUbRA02ZZdYaZyJdf8ru7Ji4HrWQ6DG6jkJsCPf/IsVtrCQnTj8
xZJSipPum0EkPlBCNZfvpTSKI44SfKnteHqf5mlzTDewEdecOz1wY+bytzUf7RWJT+b3FVuK0sTC
HW7J0/x/tDX9UJHvMCtSec/79gwNLOOCkUjWeX9KwT76AMRN4nQCGbaVLLsgja8ToIFmTXaCYT31
0R4HfEY5qZ0Jwe9zha0fCFXuYiOHs4UlCD5EeJAvX2zWYvk+vV2zuGJtmCNUk77noF1+t3HGkATr
IoYEMoCnTLWpxOwB4cdAaFG8n9WDHF8zNZf0RZ89cEcjEL+BEYFt6nXJGelwLvQzkOsEJeiIt8Vi
8gzQaUNmcDiAhymwhlFjugRNSePW/lnAlKJ85F8ryGYAG0dVhgIB5lyf3yIwFFf2bM59AvkrEKqL
rre20FsRNto/qcfCNhSf64UewnTLwZ7jI6O7wtNwqD6KJ+1flBD/pKhdVl6Vu8N0qFbElVjnzTIk
F+/JlISe8rNf4Vd0lM8pjsjMqfel0stdk4BIjYvaCCP/lFGF8aSTeyRW0/YvjxB8ifg0A/rWgncG
q4ZiNSEZ/IaZkuh8kf6+LnajwSat4fNLO+O5VNP8iUbMGHrRRkxLii3a/i4w9IuIOf9HPABIeOoO
5hLGrWrvDQqmP/fjSCQ5dhbx55WaUsB1Sug0La2HEzJzzslUOSelAg3q9gLR37A+bZjwDryFKHke
yNq5o7+chS7eiybw5lF7zCrknrVezNUUTSNbQyfT/2x9FWFYd0M/NluIswq6yFn7dEnar72wb48z
CePBhe2trfW4HbO+9jzSsg6SPDlLWumtlV9MTfg96V1gyxxdcewfGgzxaQVDjUxiqzOhpKBskzK+
5Iagvt+SACcTZFSShZrpL86X660+nBujg5SCkHM/1uxhx0wBLnDb4CrE0Lz9IHq1c3wI8CvK46A3
wXIuZVsD313sJ3H3uW3CIN897VeqSVCTBhuJgfR/rNW6LtjzsMJybA9EztzOiK3k11qUCE6d04Wa
iZ/lDKRjlva+FrW+ujM0UutRX4Ie1SPJ0NwykwlUJgsoMNvZuKPpRJZKfLxYt4rn+yc6Wn468QAH
oyGuIfUIh9H7voWJbOeWRz4vTC+ig33ZGi943kTwGjhnhSAu0W/BgndeD8OTYyMz2+O7ocSdjxSe
Z3RBL6HkLdTdGbetP72JEHM3nuMMsUzgz/2fireBGOQl1FK33KsCxkUxyPms0yTUV30FhzsPxbtw
z6TzXbaNP9ga0P9NjjapZWlsXFvdI1KzttRncFF0wdEzN9NTKWKue84omkTbPhYulL5OV9VIzJd5
iQxoqs9t/NGwbtQljtb63G11x9A7J7fzPVvaOntkOgcGvS/zrQ9UXRJq21Hi/TqjAP6Xm8xw7DyQ
dmAPxUwaG21vkPGBKSbmYVlfRzvlKmhMcRZOfKSC+IgewskYdtLrnkolZGxZVp9s+EV0K28dDyEH
VST6w5ZsVHUdKe8CXXDYXYOt5kfDiSl5OqDysD4sBF4JWZ8Rq54SBebHKYdD+d8u6xg8M14zEKSq
bkQ02iqiP0HULvZ2KzRJCY4cxlo7gC/qESK519QxUHL1huybvuvSm0gysem7KAQl8F3YL7AxwxgP
Pi6yhGREqYxPKLfWPnFz0+4Fr27AfvxcVWFjw+s2vE0n7m6u0b9zpBMCjaC66GLK5JP6MQlCobeE
+hb42UfFayS8Dty8nY/kUfeXex6ir6LyxHPbW8kShKMLXgPuXAVOvcNWKuZjnHFKZImbXdaDhBm0
dP3IPb9lcHKQysE/mFjTBq94Su+JCTzLvt0zj46zsCsz6/PUwEdAHNzcTqdoMpFxguf8lxq3PN4C
jdUfUUlOaSHlFMOc1YIDpWMaFYXSuq0EQ1XqomGRQlnyFtetw8UcZiveeZI9tSaiQzQaAcpd1Pt+
4yeIHwLog9I6r0g2SxVKVHh72j+IvCKW+KEWdbIAM0Rt9RxGb0mIiR+A80YzfkEh7KVYwrw01sfO
AtzT1JXmEcSnHojnJg1ALHJsVn4I5j4cUcDmcMlHbzNTeOemkq4MSo7dr77Wa9JWutn/P8/3NWRe
AxisJvUWzudIj8mc9Dll3Q4UT47fBNSFMPWdIKzDBQhBl9w9knKc2ScRbqJMOqHWyKvdXolfC84f
dYdpdR7lnPlqjGUGWoDqqqKuYK3OwAiBC8wXqPhA94PbwfHCpHOfc0ZqoMU6/f98s/CY8OR1Zu28
GeEVsBj5csSTvddus6tmSaZ1CTvGDNznzyJp5IoXCRXVodEz/bkNzwG5krvp1emhUe6xMzWoG5iK
TMbw6Rgr5fRdW2BDg4EIc4ayHLRTWZPX3esUC6lmldLbj+UOstMA83Gj+rG93XRgR08p1egD7jw6
1UW50P2C7Gns+9rirqiZnDNhri0/h1IstsBCPGVqMQ30EskEY/lD2wZuyvkQiCeo/vJCz4THqKS8
XKLcfnAHUKzW5ddBIBl1mX6ziGHvjASerWXjTDh4guZtYs8DbNudlbMwo0MrVPK4mtcfkCb3Wdbl
WISiMoDFaQ7YXp/1xXOL4aN6b+XFmnzxV/qckwqgWRdag0jjnQMRE65LmspRZ+4KzR/NHJKQoXPB
surtraOm7XzT8D+/F1Lwr0V26YHl9Tkz8Mx+1jz34Mw3Zo0DW/nxEjFqI8pBNbwBvzY5G5oj+uT9
ot3PG2VeLkPPHRJviALJGZigd7VVSq9FlmwQIn9eamgWshnDzdad3hkR4LG6Z2i4dwZwMcemOpkh
fS6dinX0PjsYSgbLYhjYLH+sDGLEXcUZOnE2S9CTu++Bg/C9Nnv6Er0/VVWW7k1UIeOVhDbdmKND
bpcw5qmVAThjDRMc7ui4vwu9p5VTYASLvoCM9lgaHjpfsU30sdBNzl78U/SBF83nGNizU3Xqj3pv
N+wx+njilW4Meq7TPhgapezW7oPWOfuer2FleLbeFj1WYjfs/YhdOaJGBEZJbtCAUbsUsfnbRmWf
yU9qyL/4adn/PVhlqh7ia3E/iXkx5AvaewLo7H4vKFzY4RBbFHBfi0wVGSxMwrF3Sxbxu+k1rvaL
7IcLhDWsj+3lZbNMGXBWNuYj8kCiLqSv6ao8RSeOrwPcDRX/gqvFFHNAN74DC6i03VhNsQEvBhN0
zjTDKjXAx0u6+7l0gn3R396ZTQf0ZG2O0vDCS674BnNicUbyhv7AVG0DcuTOnh9cAVV2sB7rBxdR
XeKVMiykXbpdoVR+XkuJjfyV6mktEIgspu5tcSMvtw9k+BtoaC19U1LwcqYygWLj6Ou7UxQvir+6
91reR7Kij8Z1JS6zVm+/jxiaqaEVe3xDF3IFdOSm61OIL04nQc5lTcHCv0Q/S4sKj3xcl29xD2Ls
inESvDjRO59vWfwd1Z4qV/l0ACWvlRPqrswvB7mcuOHDCM4UylkA4q0WMiVkBcR25LPPdW0MRT4+
/XNIB5SH+kqZpUrp2ShVksv8kyArObH7iqjiJlkH9C8xy4COqbHdf9xyV2Lcu+f/D2P6Mzphb3FB
PgFrL6mijxfXmrpj4FbxRXqf3rA7BXrLxKYwcVQczQ2SxE82oOnwigjflnx5meUI1gySVSDMTjnG
a+aPOBs/Q1sI5BNjDCBVHckYk3rO94CSg5aUaSXxHXrv9NBLwcJZGl5TBar9+qJcrudur8qlyGDh
cg1avVRjwtVVOlaID/hQT7zBrxcW/AXgbLnFM8zXCyEVTqtEO4ZMCVlTjybtHhzeLKsspKAMbAiV
7L+o9+IiwuJkt1vxFy3hE1cKvD6wQjZzMDGpL/s5Yqg7KMz/EftB4BOlGpk6CzRypg+clESefvLC
WQi3Jd9x5cIG2NgrXWHKplPRyzvG31i2X8uUvAA5COa5qh7fkaiKe7H7RnnvHkyHR3l+tNvleWdy
5n2JlgpwVx0yx86ZjXEa8ksFzl3Td7LGPKpjnjLQqUZXQ5my6MLQZnIgf2PDuj6xvPcV4W2aJlDm
PCS/DeUcRadttUSIcCSBVeeoUsDXu4k4V3V38FTmueJ80jwFkcs6wiyR9hjQY2+yQLwoZnufz1g3
BvvKcbmQpub5iut1zp/DrBJ2VfN/pmJxQ427LACVCpe9qQgTJNNckz/NEzUXHQa7kO8+/pfTq8Fo
9QGsuZKgRGMvJnv4rnvd1InWGUv60d+ehX6mBcQrq7eumyodLrPtMOidgueGe1loJVBV5JAz/YDb
eSaBK3M88h6KlOfXOvI2QmvbroA42aldHcdZ03yfuMTGTkGJkF1OEI5ln0mb7RS4wm+Z8P5KGR2c
kl8RCPqHGMypKuS7vhZ1YyH9CV+uMmTEAuM6lvqU+9JHV8VKmCa0U0/MDMlfVbIwuMoA1CeJBzPB
4RoHY8ayqfoiRBu+mNE75R2C6Nxf/CotkrIHvgAz3Hucrzg/kj1CO2Xa56SCO4Uo1x23iT5dHrZh
KU1PbPCpjkTJOFJ7NxG7zV+pI6QRwSE7KQMpLIAldXUCsehKJF59UNFftaxc/RPrj5OxXEqmkmws
3deGmIloMrSbo2QNdaQGNiBldx4DmMgcO8bQqyL+XOG3NczRYGBTXXc9RKhihiC9pHXsGNGNRC7A
yHP7zarI8ZJaaCcyHkLEQsqB8V7DTxSS9utKqC39vFgvRzvXb+yYfNHPzSfDNj8lf+ShEPsM6266
A/SLux2doPkhbOgk58NTZ3Zgzs92Ne/mcXwZaxjljjSSZpHNsQCFnOEjZO7A2ikuq4Lee3CEZJq4
mDd+EeEeLRenqinu7q8zT40oCOHo56bzdOGU2+ffXm81uZKrjZ/zJSfOSKjlnzrQs4LjR4JK/3Ci
/2PoHzjmV1p3ED8YN/hdw716yT34530/YvJYbh8yyQtqyy8iU3XxeHnXV+u8lDsQHs0lp/Arqkzy
RlRjBMKDcco+re+N/AV6Kx5EXjqC8KmI3xj14h7PwpSgTAJzy2F2JWREjvgYh86qTPZw4ZLn/MNW
KAVpH9CUBfN8DhoL45Y4lQZW6mZzWxghX+8v8UbM24Ql6wXs2cUtlL8boSbxSWhkzoAmOnUu6rj1
5gclAYMLajORQNKCxsq5CbwD5pHduBddEOLPWdv/v7bfQVvrfYz3RH+MoDJ3xsqVOukdaqgz4TIz
IO+LUMxu8K3WbRzKzC3bP7p+cRDc0/fQl0UsIWmhXE8oPOhAhUM6ISzKW7jw/SlpwKpObCcYfpn+
Jl6GZTHhO26RiBRJlOYo/UYRSat6Ou9uPk7WyKpot71MGaJi+PEmhzjj6dhqN/jwCejP+poFF3v7
Huqn749F6NOPbQc2PGicPJPFUQUsms25+2Q6nSttQkXzkVWFDj1/nt9OI2urE3qjlj9rfZQV0d3R
zqZP4HstDR/PASmkYxtmSTFddduPlXJLLYkxBKYsJYPDfKiKNsSae/5BXnLyJEQrfrpNDpyXXCqS
QDF+VaBya8CUz55jC6/yicBh2uvZsl6NfeRfK7ogGnKfSSexzWerd2OGsy6hqqldytFYOsbiUx5w
a3z2hVbB8MRylVzBL96/yoFSsdX8FwZnsWp7EG9M1Dp0tU+0mlLAClDQePo5i6Blfsa2ClaS8xsb
Do5Eu7nmOuJGfiHPUDmfHOf5/Gl/VJ63p5hfY6whXxu1zPhfmeH7NFqU7TFiosP2KvHdZahTGIRd
E3HmgDSMX5VHOY0kDtwhXvshwGrzT/NsHHpIUlofCNZJ6lvo/WbW2xPkYzTETMDwA4HLzLq1efxo
IBiMduewJqmwyPclmquQMd3zRwZdtNG8bgzU8GLjQcW/Is70378MeGtGTTbiYjLY9IiQ2FFKaYrj
LhHxyDowt55y9y5TCqOfDhrWg1r0mN3SMg19XqMhENZyEaPnjHrE9MJQwMrvd8n6tUBPRkSiROOW
CoZP4KWUNVmioeRNEheSxRtUS5VA8QSwfW6saF6VqlY8B6/TAw8eHlMceDQswImGglLIVw6xpbFf
GuO4KFybgHcPkE2YMUsrPfBaL7cgdlbWFAvAghif2Y9l7XGkHjOe7YViBN5XF6QUX8CkjuozxWGd
zrHm+ueXlt/xOxEX1livSrEhu//55G/F5nelLW+I4UiN/kWjfRv3NmBP4hE+PiGoJqQTB5l96XGH
qK9rZYuQg+ons+KS/HesN4xI274l2USPKt0HLxAxs9wf04TLveqeKEnD8ptfkzgeO1kgHHhxNcw9
lV/up/Xndk+NRx/0TQA+Vi8F2ykFlqmciWAj11gJ67XvQldiZUXR9OYiTQGWDzN+Ngby0mxOutTY
N65tSjcTw1jUmPY2ZHmTRSDzbWz/5r66QWqPRNP6ANCmfPggu+x3sihIYmK32QbtPfQmiZDEqnh6
S3NAa1I6QPYBzTxJK4wly3sT8hQA1D0M6/gzG7WglsYfTOp3Yx0YkeVHHL6DxgkTjyXFymS96FwU
SbF4t2AhNYvtbj7SotgFbS7dq7jwPogXs92dduvvC28+u+m2ThPPdAvm0SBT+94uGMGvwkgUqlnj
lRN0MZE/FTOU5gjt7jgTyCaFITWdeuFxuToAVoOwyzU1s5DUfY86T/n6mIaMzOQNvxx+1DWrGB1n
i72yu8xM+cajRQSrLsmxosWJAtAEkz5kQO7qadLhL/eUA1OSPowrICkVXFRuwYxJmoXblbnLSW1v
Fsip/26g6VdmaZ9c01/Ay7XvNBprnU/dX51qyu3+Zq6ewUhHVEXEzTfQmDk3Qegb91uOHpz9+uUk
jZqEoFzkhZOPC6ZC6tXmGQedjYIlB4KeAFdoXi+UzSrghCffFelPDZxDtIKbem0FKqmoUdIDGq+0
9nduQCS6Ouup1Tmdv7rT/eE7y7ttFIwe6PL6cIseShiYbXZQqOsM9zT/aqfef31XAz6okC0A3Ttt
J77qJFVKvItdtaRG8HMspXS5vx7ndxXoSFWkw0XjLQcptO0cepDAc5OcUqDU52cS/X+ULfBXLd17
oFjc+D9iQdzejC2K082zHqRd+7K4J0c6qHjWqopgnscGjighGxGYLYnm6S/qG7cthU5Y2r+di/mj
56GqfPMWY7qf/eLCCsc0CqK7cH8Amd6yxXl5YerN8sQjgUvuFyW06w6se6VcfTEDK3oDqNGjfzLh
624Nz81R2dYkIi6I0YbYWylSN1PmUSwXv2dCmY1hNXGs3EkE2Rq5F2wVSnBqx5RDIyHP++wk3MDm
TUJ2flJCPXOQOQXQnCYt62UBgLSQt6V6Lhr2WVn5Kdctdn8BUJkJvinQk+wltmckQalJ0TP0iI1h
MKOTOLGGdULb4+y5yTQDRsicbXDlNrCMznrloZEjk2uo4q55Hk+dCOCdgwl+JXz/eFwlt8lMv2ad
zBPq5BujlyKK4yoJBr6MNJbHQazySxrQQw3um4wQqmKf8hm/mTVy8ytaE/OZWWOillxpo6Um856i
NsJZQgRCrH4xhhemec6M/gdLNsyqfdQFO0qPaZUNGz30ZFM0G2tExG81vGwBSDO20nDkhZDAxjds
CazhElTuvsQzyHswfDvZzNhEoyoGbjsq0NtNzuavT0LQ7TYsx51mxtKudEWhm5eXvl4TESOQMZ9y
ensQyACwO86tdYu5ZNGPzAGBwNbrIYLvwzCtI9YDif0PE4d7kQB57tk3mkw93nbu/5BKu03w+aSC
/BWvDf3BXQx3S2G1f3CM0dJKNSw/r8dHkbM1mneklL4NZ0QbCWuLT+UMfVuFbwqDXukwErnJHPWv
tAnilBSH0WPa+bP4mU+44FskJHyb9+PnUaUx4Y8Tbm3GISBqIEG88QIbVGGbTzbQSxbDJIeNfIpa
l8AGKLJz695fjnEfDDYcLhaHEjglaVQ3BC88u0/sxLW0CUyfmB/uOe8NR19gvwTGnSKWJHdS6oYG
wRsEOjwy31wtf999ijMe117ljZlvdJ6KGNM0ghgH2hVM2t/Ra+5pAZ2+RtfGNPlpXN42ZHqlK5cT
N9AmiNcysit8CDwVNavGrwJ7XemLjr4r/CYfkzqlYKQXM1c3tiEv+CbdZDkNIHpM28j/rs5vn7PG
y6ep/yCjzGpfKBbvsO+s/vkKMY7txAVlWKbYjooCfm7GMZWPIlbnDnWK992DrBNnlyI+lkvLox0q
HavLtzBA0+Ggcpcyomx/5KWtcU5eIpuzV18HdXIhk/K8VY1sIJiqj+hey4d062XvcVBrRizW79xV
36aRVRjYjCzkooUqRyRUnht1KU/iL4ngCpGXHGd+ekaF6y4abMkByFjqws7LRKh6kVUIr8Fwzps5
Whc1OrO5NMknbFu7QhF9kprfEWF1KakPn46l5zXIDD+6u1epuYfPq7HwofBu89ppYzGtLSwzkHuU
XDEA3lKQYF7OWDQEAldZb5OD5n48a9hDSCdm7rEF/5fH8Pc5I9y4Rcs2zzgFOzM5zPf4iaEDKThR
YeLKavvu/3BUHuc4HlbZwvMhSaweQqt+WgR37bWgsTIY3YbPHbmjRVH6qtpTeWR/qapYx5mJDp+f
fFguQ8HjIWqAHhKAmrjDOTg/e+N0sEF7PqPKUdWalMVKrJ6oMaPHzA5katZZiK/aVZFxQ9AwfKk/
7ETI6jYKA8LMGtKf19vGyzdQtdEzDpcuO+guHxhTyrCIuOqo9qNpJR54HvoEnbhpV95LvJ/kMvik
G+6dvSGtz1l7Ar8b8v8lYqsMDP66R36Vpx3NFR+7TaaevbnnpQMsTQUReap/VmRUjbfo/2Atp9W0
jdeaO5zGZHgsrbprveG3it0/c31bSrJNjptWcOF8exB0qpM4CW9dh2SHR8GuPIpcfLX21XII8Igx
iQ6DUzXdd7ngiD5/LsBvvupCKD8pc4XrtZj+ir6nHj+fA7R/1T+4C8uveNvBgeUmWQfXOW+b0CW0
TXFcNrcenk4J3qDxeL2XIN6wTWJ++o+XOgs3C++kevb76x5vrZoir8dOype/bD9PpbflEnkOFC5l
A/hwPb6XFB14yjO/IxbOAlFzNaI9GJNI0oOskqoG7rqip2JK2W6Mfz791E6GI9QQSV651hsxnkn5
ouHr3pJsr51ozoElyGeMZLIfYAHrKHmiLi17KAg05Iq66fSJjstFPJy0fTqQioAyxoZYB7zsjvgw
MjBSb1xmJPzi54DoJe0LPf5EOj55XuNvn4XG1aZ8CvRcQKQ+p18a70wGIWjf03u1mCk+pPfbXNJB
2qjoSf0qjiXe6St5pRe2TYplbdH7oIGHFkPdS3GIiiAeDRF8WC67jABr6kpkWHV4xkGYn4B7rboO
niWVXd2N81xIWVK6nR5ylFzj1kMd7+fkkNb3yBWf32vivELQaK3etiurC7/T2yT5q9JzBkBjbGNc
P/Nq/irLZRjvTe2yCFum2Qu3NHMr/aXjb2LQLNMr6+Z7W6+qkMzAuUTuDKYaEK3lb0HgLC7LF7v3
JIpgsmp/RcWJU7Q44nHcdeRq4euZTB7HLIvbKGdzZ5pl7F9q5d7wbEJz2MxRN/SwsYgEidIgKOn5
tBmiGRv2X9Yscqj5ys3aAp5K0hfNy9oqr5sg7mHe8z7We6CorBVCVAwkRK0fX9Ku1gNCERPbTr0P
D04GDeRg305ayiW6RshHguXJCRiBU44y7srh/hebm1A0oyxWmk/4CFdulFcJGNktdh9KwMTgA3xZ
I0NbsMucyYNps78I74tV0jdTa2nMNKfFIq/f1BQ2gySWoZmzbOOjCizB6VUU5LU3PfjF+Jk9jtbU
8+iLePMmXgm6S3kNKLDH7gRG8oPX4xvlGUAEIG2AQONJH9dgmifMKWzmqszN8ViPsyD5asEPQSyK
a5oVmbm3N+VXJmaVdgpHNSJFaF3eDcFeCgr5ZVXPLPf8FZp3jtqS0XIYGk9Dtvc++IyCniBgi2MH
TrnGgr2pT61y8zh+ulWJwmOoEYMtYOoiddJXC/OvcX5uFLwcFTfLfZStPuQfNKNapqVJawagulyH
NMbZVtxKcpPU/1W+COffJl9eeS6VaC6ceVxzz2HP1xQwMVHmGli1IF+xBJej/xasu3EuGkxpaNe4
xTplnMibAAJki6GJc09MYG3Lq9JDyW737c4w3aZ4geyw6o/H8WWSVr9bdjXfqJ334wqY7+yq0v3Q
aPRIHvAVmXvZFuqKdPvTnXhDrW8D80DUhD0DKNtuLzRILdXLTNxG1nTCVAvOL5TROy4u8I8GGuSH
MclW12dr+D7/W9FDJyYywhcYaZ1T0IieMcYq9wfCQSfmV24SlJ6myny4QyXnIXOCTGW5lWGzturo
RgJy/eIbs1cdc3BSZck7YZzWm4Bqx9BWRrt9ruzvbw0DAYqEETNy88oxINeNLM04gf5LB4DaCwjd
5QyC3RCGkWMsorMyKqgPqZ02ObT6/VHr7mRHFCH/j5iQe5Z+oE3MGD9PS1KruaWNhDZ7/XFbDmxy
nVCz+qGY9FvJMYJ9wuVgnYu8ZDKC5Jbil+MrAELvsbdM6KMQ4X0OAXLeEppDGe3rTHiR2PIQUqt4
Q5ydnfeENordApCmqvkqRdO2wUz0UCm6H9RDFJYeHx4ubjNvxSSrElkJsBEeGMg19pOtfwiunZWz
9O8iw7YdaZb9WVOj51MpUcBFm+UKuUYxyFZzKy+XHp8iJYz9rWkZJTFfdJ8ek3uA62TO//4lU1zC
CVseSSwDV655RvcU5wtv6zSUoJJFj3Phxbl53TmsiXvY6kAb2UKbexbNAouqfeBmRs05Ga76BB3o
R8rwulsmncYIkVH18bSZJwyo/0IXRCRql+QuhzIyzaY1wTnJP8Y1VBiAkNTUFMm/LEK4LZy3fsOf
nkxpY+oJ+MNLfYzptrqgMB8zdJ1KTchNvriqQ3TQ0AEjSZbhdtzTRUxyhN3LKJ6CJ9wJ+LZlUZOf
0cKZCdiTYBIw6A+HdNZM44oLtyMryti/iEXBkQy8atW/dA7zeZL8R75tdsTQt4KfApaKJgo/GdfK
iydzRseqVK5e1ZehVv5Dmn8i2K1NCIiJ8HGY/wDTYgInZSzs/HLePYziLr+MrYjyjbPfiqvvv1FU
5kgIXCGG1XMZ+vurXRg2i7/M+vgYy/R6o2H29D8Aekm/l2UPT4jlLiicpK/ffgY4E+77Ca85255K
D/FNCb1R2WsoQQd/rpWqdtYfEJwtcITAKlOQ303rUviG9UHtWA3GiZVxl0XZR9BVZ3l/BTMHGs67
8MkeOzCClrVIASGFEOWgdiPcDk+uNnNLr77Vg0ZvoCaba0dMi0swl3ab2BKsOv50EYdCLEaiJvvc
WW45G/tW4Ju5FgqGfhfML5vfIEA6+kqcDEmNAaYN+pbcCU5+xFuocOWUybyqNdA+VTkiCppx1SuP
x0iOnUnA5LyVCt1zOm8AEoWOmPsLe+MutTcW4ry9XD1n1Xm3bF8QKI+JTSLUh/E75/5mZZNn86ao
k9GFExp3Fh7guiCgg5xp8zGaikOa8DPN9V+VCQyNxd5LGpVZfEi3KF3pxxHE4938QBZmI9u4p/hl
WYS5Z9S5dNRNQRypQh6JoB4jpV34Cs9G6EIvl6R/dNudpBH5hf2iGqQLs6gP48KptTiqhwmdBLkO
2aWODTJnjRzZfsRiyAQ1YT/dS4n/0Ctdz/CcSjTE0v6mWgFMGOwfWx1MaLsJ7IKxdlj3zfyg5GGs
BNTNcDyEfWKZneeo+64UaTPLwIRrIaV5MVklunXPWcpMgUyv2RFHhs4a2emtvXHknMr3lHln2HS1
msvYA5ydjiWr1R7T3Di+/8IGhS3aEPEmCZ6cyLrNIvoBxzJxU3kaNWf5KqbjWRdgBzKk+RvGvseQ
1VCnpy9QZbWlpXL/rnnacONR+ua3Wtc+LjkU3mmc03RUofVa0TfjsEDxyFSUd/ZiV8RVmeODLQbr
pu3ztw2AOEYnrN0YSjRLXhvEEGDBycsZaaLFH0MzUbyq1muwkBNIsbXADBHBuZOzcq/t6mwpPo6E
7/mTuzGSZIJMTBtCQsROVqBG8YZ4WQ3hMmQL2wOPGFezMlcQGgCvjNLcniYQqQod2LK9h4jtvZDQ
oC2YKzwY8+Mv3WUt4MI8xaa2+qvzlDbhydwHX9rGICEpZe87jlM6Y/IZKXT1tf82EEQZhb2TA5gm
N7MmlngTZyU0ydzvFk88mmIMHicvuzVnR7gGhFeTk09owffWIhHmwX6c62YZo1PJ+gqDtdY3Cj1/
TtN8IoMzt0qy4ssF+JJs2P2ctomWlqqNJl+kYpcB+dWDfrnweuQFhZu+aEgQhCaGqGNKiW5uG4Sb
sahyWdXyqItlMTIRG7gY5uI/YRykqrsKm1GhsSk3ycKNHYFnvHtXoy6fZ0eEHpFTdqimerv5ZPrE
bt+u5UeAeO/yPT3Wo7K0tvLPnteNtilf5/yyt+dm9AKmmqmS0xbqQqIuanOWDsuTLJkseELKGFVR
BNRynD9WngzmDiUx/HrjaWPZ6qejDarl8INijsg/+nqwgMoW9IFfNVb2v/YSb61PstJQizLx8G/5
c0hx8gyCqjVfKSitiEV9jT8elrisbXDV+2yFUshnDvg119Vy2Ddp3hZjDssU3al8aZXOZLTKDfbb
Tkm1H/n5eYyfMkMeTT7Dj3L/49vtPDTJp628JRA0taXq4wMEBzE1mIpsecLAo43Dc1apULROj8sq
hHoW3lLM8Tug1Tdz1RXXhG7Dgt2vPsfj6nZKgFcKrEiaX8fkn8+gq6SGdJxEBOW9sVGbRaONw08m
ZYppTJ/hc4bueIuVyuJz/ZJvoG9V1OZFBy1Qef/MULY2B9wd9z+32JAk1JKWeLZY/LhK9ku++IFW
JRM826byZ+HAZppofFdeEGnZGlxZM7A2Aaq065ZjnCpcRtaWJSMpsoNMXY5+NVV0MK1kBNAuyec7
KUoTAUvA9kmyhPnB224sXWkizJxD6/lG6AOd/TloVumdy5sOi+WlsLxJYQII76qpEKEpJ1MvaysT
P5BT9TUdv6XcbYIKWQEThcP3htAbczwuKxNBKbC9Aa4boZcMb3fe4oFadCkeLcEhDanfBfLHfG3L
hNaM0tEdMlPPDxwZFsSE2Sh9a7r9hhCdVp+fQxMu83Z39KiJ6uO8HR2reiZI30+mVFa/uVfm+g87
laoPlYMUhU8nZTv/0Bzy7DuDET3HoJqs2Og1+vAloaINbJY43j2pEZNkhxwpruvR6J9jf/T8mbDe
6P6YbmqHA+QIU9Vewg6kXesVnYqa0lszbBxjzncyYbsz5cruyR/+nrm52YaWnrBwKheo9itKtlwq
504EYCEECTD1sRHXTcMV3RlcVYuyJ95DE7lrsCwMWZEPpA0KJbwvVay14az2GKc8k82ZXz65AlN7
q7El0CDIAPa3YqE92vut8x+WbhjEcNc4v0t/Z9C/RNHh66yWmcqZjI/5dfp6aIJUNTku2jHod/T4
Z2qXUDGx+fql/tkQ8HvQ59deNs/lpzqKCv+LCtU7sthvYRr85Brr3mdV8+6W3NUpYhuZD3N9UewB
TJcc0UGIg0p0lICSQcpDLpFAofqBpBhZXGYzIZuDyVgALr/BVkneBylacXj5hMufeSNjN6m7e4H0
5J3JQByc/gVcGwZIEPiCw8RxyqsruOv2ZV/l/AwDMVkUpXGaKaCriSsUQY27H1+gjSKQ/zFrEK8L
sy4KM78Beaenhfe7gr10585gJyCy7v9R4uvJns9qiTCH01Vb5wc0NT5wX8j8blGn182RQzWHzIQA
0gu2h1aAKtTuEgezCxFHtHB3Q0v0Q4S+J2tiIF5GQmIf297HiHJ88bzO6+l3VR2vMP/spgBnq6In
fZ5ecpPpmhjuS+4/Iaiao6ToXat4tVFBJCsu3vTiMU8ge0NrHrV1MDSa9A3bJkxKh77KXkRLFzMs
Oz1FS9A8shoi8n4n4D2YCDo5YGjrArSEY7ncd7hHfNSaTDBcib/JYJDdckKOhOA+eeMaX6M8ZNMP
D9hBcSGK6qL3/yQRfnJrMb14HVJofxkeAzMCdm2IacBHtcXa+LdUiiMvo+ASyCOUmcF8JBJ36ZmI
Z6dCdSMflQtjMEpAUNoMn1H0WBFi25x/G52oZqHzGTpXJvVyjphHdZTOV4u0Ky1RNHZkazJGKodj
2VkRfFxDGeSc9RLwsMUKpisAGuAmZQXo/zOlFSGy5mNTWN/a/NkWWhMrP9U670aw5AYzQEKRS2lW
ggocu5UiNljXu1LcrcDCZlscYs9Ie4IX5i7JvLp+4h6GMwElG1kV6NZInHQ9tFBxCjPyH0BzC576
di7uTZ5ivRQtnr5zIP5038sPZ86k0KxC7g8UDNdRywKKNtbpRycFuyTbq+Qj58GquAKJuDwmi702
S2jcKDrMUkHpZScvDCIKB3o1CAZBP2TCf9JczLB0brsMrNyeq3HMSxwAYSTpq+Mll5vHBXLFh0CL
EsltoixBtx4hdDXoOVSJ8vJoKrj4VUqugixM47v/48z6jb0rKSdclBgd7MaLNpPx2VJjh1Oh32Z1
ddxHUnFD+UjaRRTuhKL9g+x4I9R3r5htYNWkYHHisUbXW7Vn+46e0gezIr4qCl/cie7RpwvChByg
dSFZy373f3HRdEBHp9pvq/BZlNw4PgvBTOfLgNwTo8XGP/WmFZ4vQ11Rccws7qw2E1L+1qpAc6fG
L0ivBf4M3JR8vsU4n1SZsGEAOLnGkIyj31Wq0zfqskvCARy6jUMOQefPtFXX+++jHArV4fT76daz
XxJAOm7EgbA7XBJLnXd8GDhep4DZeKFAy96XkEJm7CWDTrCdztpdtSYpLzPhOP2LWdkSJEmGUBS0
gY7NssnIZuelPfgwlZ0tC9r3rCIKtABAOyusWsvLXpxSxLD2CyK3E9DrBXATvP5VmBRii86xb37z
SW92VXgvA3ogCi1fOrtR5GH0u0sBgv4J3z1AYejX5h4HwFkJH8usEfaVF+1fUOr/HMTsQiu7hJnF
WgVBn+5ddjC9+aHLXwBteLeFjqaoZ5Ru283uuYCE/1o5bWfeCLZt5Fz51DsqtrBcFQMAxSGBEqd5
5D9ap6uI+TfqbwKIPnQePP1JifBWkzkoOmNiGtEcSfyRWaqJuhH/yDDrNu5Ut9FYcveK7BseXxOA
q9Rk271lcvc9RTeRrpv1YetRngmFeCzvFpknUUfaXC7XEXEHE3ELQ51eq2UqtZqcp/kWiBAEcONV
nxb1WD+rs6e3uTB1b+WWtGJkq2YqWVR3umP081XKvQPMUhVvRxTUGhv1Z4vrU1/TRro+rgL1a06S
JetH8zxM0a1uj97+FDx5rLy1CPSdDIAtL/cW+tzFY8TxxGrAgG84nkuXNlqGQP/zdvBiMU3DC5xh
C+ofz/P3my09ygRTI4wIz0+pLfq/iRRl4dUjFlbaSLU14ukqyl7my98XqmlRzWFhJpw21vk5gIHf
fPTG194E2hBJ4R7/neN8btBQ/5eM+sBW2eGj05LyFLW21H4w2+25TtvnLT0U/1bRAh9LfGydYHk4
xy/MHbvVfYV4ZslZCxfzme9SNtcwGzt+5iFmL7lS7Z8WZ1Cg7xbpVtZCsY7IQyltkZukP8auU8gH
lh0KALEtW3RLI5+Q8mE6wRw8MMqEITKaynqtnwTQvahdFgVGVmmApNYqF03IacGa2c8TOFli/K1u
m4trLD1QY71oV8kJhS7YcQlGX/hhOcik1wSbhMoLKblze7jqPvwUjrqDA+Zi5dlVHFAiXcuY5s0/
Gm57xb6vTsT4qjgpUzFL1yzI/My3ATvf/ygd9a7JTuH5iQz8zeSOMQr+X2ZNfWo+ROBmEE/FwUft
jyi76YU/RgcuzfM1EsEEhulpnLsPol2DVbVGXIk7kHUIPqn3sUg5VfoT2BZS8CTMxBcpbnnpezM1
PC0pT2yABTeTAuV+t06UJQVh5ecLYSYghkPjV56YxCAKKf678rAgkT6/ZjtJNB7DK4Q5fTxzHBdM
LcCcC17BYnAmVbLoUj8Q3lRBKUkQDvaUdVyChrXdmzXcigypK07pythQpLDVu49YkHddsWgaGrnx
WI5P6f79iSiXDq28HZFPnqea8iSNuWPL/d1+MtZ6CVm/V+kmDFwezjLHJo/sWEsyYpwDU5miYmvq
sAM3Pdx+lk41gqiBn+DmmFwzf5JZhqtVAXyHPAmKmnSexJ5qtmHDbTAo1DxMvL643+smCjSXLBpl
D88inmTeWrQtz1frDDIOBE5J+52L/X9Zl4mKxeS8i0/JsP4oaJUhV9KoFiS6+ssDNRrZ4UCWws6+
5S2f7seGZ6LV4GROVtlZryUqd9gvICsTLAoJiq7pDFqlAYccs8DAx3L6ELp5VzLlqNCVIqaggbCj
zlNj7DgXDyOurlmk2+58n6X3+gCJ9nVTSizTFvJSs9LVb8LKuxc6d+k4YX8rw6iJEyeIlW1FtRFm
YB9VqbYMwcZN3vp0CvA7bIGA9YzDX+BVeSJqub9d7dzn6luUnYDqkekxWNWidim9IBWO62p/ysWw
vv+HUH/W3eKaHtIX9evmJ6jdErNEoEmjRhriMIQZUFMIMxxIRdeWg95LWBH1cEebbDK5qWDj3F7T
yyN1XQpdiEBHL4/rbAWlxmoyVPM+ArS5QXchQkv6qgJyKd4y2SsnT0Tkz7XfH2RUZ2rvHA0nSKIA
j/gGQ0eJCJ2hg//8TRMsGLKKwGbU3Aa+mpSPvhmwKi9NqBhi6XKKYswbUkU7qHfhy3lATU1GpxkF
9xvQAcBT4xocScjalhY+QUouwTR2WTGEoBZBbL4Og1O56xrClIcyIruT8ibQwj0KtNh6bdGF68xX
X5qIr/VJ0fbjaNyf5P8CN9OPbiw9VWIktvpkv8KyYoNrDg/OaL6wcd8RDy45nQAY/9+eAO7ESiRA
yTSjMhT/ocihr4hFjsc4ue4eWlBTUsGiD6HrlVMDjdsuzC7bkQOdgrcH2gqRK5dSFplEHLC/cqGu
OJpcMstvLGBRSt0LSsU7ydR4q+ELrjB6JmC0g5+hYFmHtVYpctqpSON81BaczUwOgwVocobz9zhM
8EmHJbv+IOHy074WUBJz1UrEIlCsBh1W83BDlkm7sMvg4xEDPu4oXjy7wy8CNnrakKV4I/CUVXfG
m+rVsybqFEIkgZVkpnTw7kqbtoLAOu9DclbcHM+42W3jhtCx7XJ+Z9qj5PiF6WzCA/2Qe5d9fl6v
Au9uhUvhgdIsCuLBED7mAjzptFPeKkCjj3cslwuFQOw2RquPtZyeQ63RswdG1dnBp2so5DF6FnES
Yjdi/4IEyUBSQJicx7XkMIOOVeonukgOY0uPdt0lwsk58kbWdJPE+3P72NZnb7+bZArdc69OQtuH
8JSyXPw2I158HqFBT/Nk7dXrjzUyU1HXD29XLGm4E97zy1d7xo7/2wWXH7tpV1sCUfFPxVTBjUHV
8wBiS2TiaDWVnCw4z5Y9Em9LKRKKO1JoRPoy4stpkx3Hma4CoE+bHAJN0eR+25TnM5ULSBDidibK
hXSteJS1R1UGzVyCQG8WjQZeooHqt0FE8SyvSJFRYnSzxSd8NnNrCNInl7+R6n+g9gbgUaU/6lZ7
RcFjwm+Ir1RxqJse1jeBW6w1BKXh2nK75j4JmvxwXTd02GKvJSA4adRMiegbVOVesvuxHqs2CwAl
7dujCUv0uo+jj0fB/qOKaHAbxJmG+wvtb+xxzOlfF2sDE88VmZTvVLjhmjpTGU3XZHoV9avBaF+m
sKvjzidG6yS6fvHa9tRq+Mp4l6NGY6aZnF1AU4LM2yTbK6cFSVU1PIxw+uAu3YM2SC3GVZqndVeW
BcfJaWzBtEY0vBuROWFF/v6CSE8+OtyqJgVjRC+CeGIsR5MgzK0ptGomSr5fJTnwuc8OJt9Nfxxz
YzX69NMUuszZeoJFsyaxs78qxdWE38XAWnVEg3GkQJtjaKnZJovG4mMZbw5Gfmpse7VHYqZ/s2O0
GjlycN1wIz+MXsqF2u21v8SUOAw+bnjq/ATlFje2ZK0IjNZf46K5VSnW/IRRjJjzyFpDEZJCZj9M
W0PYGOpxCpcnBzTsigdwmVVKyPi76Sj8aVq+Mapx/KD54SxEXmtcyh7XsckWQO3MXDfmQ4sR6CMn
lbwlErHfmgfjGEsodeQwD026SCxNBqDZoq0mK16SsVteKJy9s80RnHd1t9t5Q7UoV7lGHZSiLMV4
gHwh3Wz6RLZYwjsD0aYEKyj4mKnkh8URC8aqQRcIPpjvMAtvVBaJeNFteA3rq4SCoaeYkzfkDzue
FqC30pmCgL9nL7q6rA1NgAwznSDYVRceyaBgpN2iBezX61Fx7LzugGIK3kpPrftGe4GryIk5RJt7
Wo86t+XIwmPv+xWSBJipXNdmv8aUFWdmHsni6AGeKJ7yYtJJ8XfpIv15VYr4zRtcErkVWmYJADZF
54/LhgbXQiPM3eiGCpcs3OPdk6HWVREBBhKXLg1PK60tqZauJURNGInS1WTsInO7zkMFK5/lfPTq
6OLVdlXAH5cFoxwNRujhwDhU8ubBHPn0e3xatEj07OmAFFLClG1dP0QBj4b7HUw755VFniFpgfNY
fj3FhL3TkPVo248awadu/OgtNW6p73BJCB01pbDmEaOThMnFOvckVcVMVvwaadsA6AcX/rvejZUE
xKhzwXMxPqwf87emO7Iop74DU0O621d+zOAeikB7TGTuCFIN2+MClHd8/FTbHjWtW2Ffg5Aa76CA
h3VLwOxpUgH+gCS/bbftupqoBwroe+T2LypYo2W24CmySFpBqEpE/lyGhBJ5gs7Ncuaye6Xqgb7H
Hma0jbNxMtKEYxDZjmjqIj4vLKhC3d+ldbfYcV74YXuDtXvzIJdv/9g/fhFcK1zDtPMNaaal9Q93
quo5/Rz882A/sESBK4vvwM2t3g39LNycuxOZfv7vCX6+30mSv+Wh6rqqnWnWlDetVEcl2Dh76iaZ
ZYSgcoWnTcZx7nbPbc8Szydgj6PcZpcyWrYSI5ic0G6e+VeBSMWWW1Nr2IoIrTLON2bRVPDrBU94
zL25eaoLxJ0CdmapBrjDXaqig0VwyKZMmonghmgcqj9jGXTx4O/xbyj/QxCgaszNBAIqDdqI6rGH
rQEf6QTAKnIViiElaVv7Y3JdJVHRSGFKKYW6Fi/8CjKbOi9iduNhD+Mp1SHHYRpRAh9x8KPJ7u5k
bSHoN/ZfuaBiNqL3cLvZ/D0lgQfdH3IGIsRdRFzPckPnpxURtcdejrtwF2TW6a9ISyx6GjsZViMj
Z36b+XOl67eEjzmdO1esHeeiw4HqVX1BNTVECDzOSC5E3QWbaLKP8YEjLvPM7WKIjHhVdz52NQeG
KA3cfspyAhbnY+jytSks77g6WsHG7wR7abPTDXRt40sI40q3szj0ih5YA9NQJgKnBS+s5cq2DMCi
XgcNx3MPZkw4rNbiRKyffK0MTIgzOI0rF+awCi39NqPqfzrWP0vZk5VuctFJZINNotV/sIXsHRwf
fpN401fOZENN8jmzaaOmC+EN/LLCEbfZiNiKkQglg1G1yP7m19SnR565FCbPzSFhgS72ONPF4QsQ
8YsDMI+hhIA6ETqdhXFb2BClYYtjLTaWbsvAOH0kodc0VwavbeTW9+grEInX7IXYmP+kn6rEQSpX
hSTHzR2TH3X765yyxkznbRnZgRhnWRvb95TO/pZDcdOhVEByFdYo6yH+CF/i74yOcl56HsNtOwiO
N9nkkWqkEwa78f+f2DsAvaI0nYDL2SUr5V83gPwfGUIpbyNgSAkxDihTDKEBg72Ga3q6EgSWq7eg
dg+mECzyIcd87rgzsCVJ2JcI/G/SEXiHPtCqoXxXxcATdeocXTcEquP+JNhYlkyxyfo5BW0log0U
Jfu3WpS5MkujB9tZgQ+55bTimkX0HStc1EkKVKGr9uA29sU9+J/iW7+ouNlsp0UgMXuYlSwiJUEY
lVomUAUpw5zbPd+GQF+wl9jd5122Eg9EmC9Ul1rGNNSOi3hiaXEY7Yn7l5KFwGzy3wIFlqXtcXOV
Eq1AxCpQ/m4pxbwa3xYLud2P7iy2HM8CGbmFVAEAHpWmtGSU+QQsb70d02CIupxX0lgFfoW6JF3C
QvUuqP4ggb58dFZ8uo/8G5b4n079Ouku+Z0S8K9DnEVU30apykuOQY0YBXNot628gLBsrqg7Nqg1
jB+KJGsJfFECrm3I/GqXYqxIDzdHiJvH4mrz8/vPjxge+SapmJsnI/kmZC0gSFF6T8MLPQSbo30y
xTXelK53XfCRC107Aha2y9EW2gtbe4G6iWMWkh1THnrzK8txAdg25LZtInqnlhZsliKAXgxjg7OT
C6fffL+/JQIhKQQC1SEkDjcku6lebFjbUZ/KvIp5cH2m2Nl4D8mr3uNk71kPLRWzOTqNdhxaa3t1
Nm5ZZP0zOpiQSlJKrI+eOyZgT5u4F1Oyl8zaxbm9flUKBvURlrey1mrXnH7d5Bo5D7HqgJ0jTRqe
0NGsaK9sooUpr+xdwp5ZmWyeZjnQDXQqY6LCztdVN9ryhGATEW8gIz0gQo7QGl0UB/erit9whGki
YNzB2AqvdbJQ7hHeDeH5TURbsUxzqYkoanmRbNIJOJ10xnbr6uBa10MGV7llhAjwLWOGwz88qGx3
0vqN4bd/HgXC4cOzSSGuIkXL+3S+GL0z5G/MDPWPjCDXnXsDSRWsJOj45nzIeu2uTY3AZrO2XjCD
k77vXb+3rZFqJHLrQ2q9nq6Q6y9z+wUJO0y31+r6Hc8kDz3XaPBeRAv/c/kRyHav8liGqE8nJ2C+
2IvaWYWe722OLu+XVMdmNF6qqhoobr67L5NZ4c3Tc7bCX81dr2SWCTGlVXGlf4ASAE5q6kcrZfzV
0EpRoiKLE8Nu0NdFCa2zZ9In/7r9GBF8P4uMbq6CrPtwDpU4QCLEVGywkz/OZuqo3bSJJQkhv6Ea
NmnhMJjdqv5Iv9gzsrx8zQZd0TLookYPDRdJLAABU8/px6dBDEPJ5wjyeM9OwPSLN2Fs65pIpQ+s
RgwTgbDfjKPGfsPphlrdQa9BVkvyIziv4ITC56UiKcQxTV8pa9eY1kaWtAq0JEbx4yhBWldFsj4/
KAX0Y/xDiDy5MYU9LYPnbEBc83RQxmJQKasIt8SQYw1744aXElzWzU5l3HiJh4PTqvt/ec8daxPK
8WDPZbF36fckh/w0uzSF/jENhtxII2TrgxrU/ztn3TeY4nkMNFMyoNZjrSZFtNXlO3LKbc2CCIr9
xtnAxUmJ3uE/xUl771k2W+M3OZaQO8B4AxZs/G3u+E4PieaxqyEv14iDVOirdX537fBD0en6aJEx
fMoYMfKKnaWzYqlU/KyASAAp/vsWXLxJp8iLw3O5SxH9JdasrWvHAgCEDfZX7EED4xf7a8uPQQ6+
PPuUmPL4XpaTU5jqZUvX9xV44Oj3x/RT47Of4hFh0xdEkT2dNschUfZuJMl74xK2OnrWCE6tSP+T
hGrLVzyTzZ5EeGWIrfy15X5DrY1iVkN3NPtwFxcoOOYtnYspNhnTGXSGc8TFNmJGTt7BdVJViDKT
yHM0TzKmIa+5tTlwGwLMADOqRYdhYHVsE/3vh33dJa+1R/bZckeXlqSRNdjErERA93Thrz6b0wDR
L2+s9t3Smp2AHgzXCOL44vtVzN0+6LfPBIZrLsxnF1TiHDmtJidNzRgrdeBYK2YqjLQoh7DnynF4
nZzUfbiLIjGs6QDilkoRX0Z+3aYoEsDGNmO+lxiHlywtN7IHwx+D8cCi6dWeFZeuGeBbskVsxX9n
t0f34gJqiX/I8J4hdm4HvM1ZmiTpofkIratWVvNO7docnfhgOcH3fm9SIgscyXB6x8pQ5GnjdHXt
GiLuJo3Wi6rnWy0QumChCfH7FfPryX59f9JQjSQGUHk15zOo+aVcEi2LZ3YcYqaJON9N7oTmq4a+
XqUNUvogHuBXSp3S8RokRxKIpmv1nunsBLXyS+gLV9d9k/VNbAFoNVva3GKRHSLqlW3Pm4sojfSf
L2XOl1/4gkdkQKK5DUd/Evz2UImcV5ESLv/jzTNjKx6Ij/Fa++AyveLFe42TnQvW585p/achxnyw
8XVEmz+cBxr4wljz9ZJQiUZoDs2w7hDrWF2RrQ4nTyP1+WSEhbHLtq92VzhRmfyzpOXrl0kx8TSC
5xl7QTeA0Zc+J9hSXIVd8WCZH7DtXj2X/d3RTblhhIoDIBcA0xLxEw2XAKnrINRewMbQCNwFl6cb
rUj0WcEuWrxvmDTT5ZSGAf9Hu66xXe7DTMD1XId84efBNOad1koiR257bxcMIngFiNGglY1Ghfao
MsNvTyyZfGX9TmehPyrUaGhJr/VS1UT4VjV0hXczV/I4hQL/N6Y8sTSNDVjfJvi6TaZbJqKARgEp
qzYT/W0scEzvac0uT/fS5vVNg4uDnqG7JrDqi7I4nu8DAb0mzW3kq+S7vweGEhrd7N7zgdWK/QXd
0QCF2JOLM6+jwJvL0/gAK+b+e8OnC0fGO9Jkl6g1ZEBFwgwje9sFc3lqNxMGY/1PGgTkYzfOS8ru
fPSlUBpsPW/SDeHIAQq+LritJt7NVBDm3PsBRpoLYca70Rn3dKIfySxEuoO9mfdEb8PqRExbkJxl
gpCQPlll+/lKQTW7AyKMnNCBjITMcOUJXaTDGLuHVF9uQ9d5VCqgF22Y3R+zHN1JNw2xYipklDv9
0hymlUOiu0B04rWb2y3I1/goUqVZ2IRkQJd/QQlyLEBx8Tg9exPRRxuLOriulvWoKnc67lrdA2sx
mbMpPtjO9kXJzSbNxY+U4fCP+bTw9WranCZZzG69prczmbsNoZALFm76k51LWzl9+2tzh7r/4Fcf
/YR0YVtdULE389G+wZ2ZX0i3orhiY2d1x5cfIGubgjbn4ZQpVrblizsthAJqEAvRSKNmzD8ncdQJ
0OAOWm9QtDa4NeCLFIIESWmL4GKznHf+rKpJV9AsmRggGwJCMwiZroOL2PgriOlAhyA7bO6gnF3c
KdHqVGFnS9khXRSd2AM7v+gR3u30/Ox4VMMVoQSXHEp/IeU1AaS0uI9XykAW7sXjlzoNQ3wigtkE
46VByHOF4+1llB1Kk0vfMOJEqAQbbqz4L4zV7GioUC2SC+xW5MziUXLJrKo6o7YE+XKLekGHcQis
h10unM5MDgUjSqbVck/1uNhDuGDmBjvkXY19wEpkLzl23puDt3EtHZvcVIemHUtU4SwdjM+5t34L
vFg+pMb0THezuPlZqCVYJTa5eZx00MMSqdAK7QT75w1ISdHcmRiRr5vmm6NOGcdZSy9OfJMIYhpe
XeF3ubrTKaAlXpigY91P7cBT1OyahKggJkx66JeFhHQwyywpBG/kxexUEvXLlXBchPqgVpdBRHcT
2AYC2OMrEGNYLWQgfeQUwUXGt4iaEyx1uJ8QFGhaMKgTwPipj3GOaSTS8Ml2lBBeb24JAIDDXtCt
+7EZtpf6JWstDXqP8T5fwzJbwCGYEAAxs4ss2CLNLWbnBylicMi/XZwQuKblhGkHv39FRfaIsoIO
OZptZkBsglB0KEau5K7zneScxJv5lkbam5sBYBtNgrpWHKfDknhEmpy0ahxG3buW+9GlaqR5ElM/
TqUCC8OeyqnK6+/m4JKdWInXm8/9u/o1E1ZREtrk1ZHZMY/7zdQRYESr9MJfhSSGyUfNwc2z1OM1
cBFq23syLs0HrriyUzLb94/YwSiLo9OfVWNs6AlqS8nAXmONTtnRhUXY14+Q1NWZr2ge2/bALl9Q
qNpfRuFJycV0ldsI/1dm1z/P5OQFS/ESs6KM0DrhKI+phYnjhPezC1iIuZ3+2yUovoCjAHKhGOzB
8c07kd7DLiu1Qdn1LgwHaErj9Cvzhp+wqZ/RuKNDbV40e1xjdKpONULa7WhphMU6i7aRAcRiK4fy
G4PqjdM1tBZu0d43PynbDEg7g3BZdr/Ug51I7aVjgIZ5GELaAjJbO1vtjByRrHpXsc7LNY4QSJkH
M5fc2y3mB7Ab6hG7K3bFjtFac/YRlyjIu6Z0YXLnABEFBVmWLZWpi/TVAZP6BUxmHysf7T59cfe8
EjsatquzNFU5/1pjGWJmrxBCbWKGuPaSxuwu37YlEGQxHkb6pT41K+M1uhwotWuTn0wyg6vjteae
fOTdkL85UsPORRboKabYcwFFOkAD+CXkjYDMFDBUuuWy86cbriWwPLevEjt9nOFi58KD5ToG2eHI
Y8lGt+DVfyu3zCvsXHKB8UtsVl9hXJv3ZFNlkwBfCh+SxptynNaflIoJtFi4NKHU4zLVfTClF6dM
EW923zIqttoUKPH5QwSMpubNkXQ0q7/9UPhMxGbp2JjJ8jaOoXhYfpJHmMUn1OEdkwXkiJKl4tt0
oxnh/epQ3UbzpKoKmutZSnm4Eqgk6kpSvAyWQ0FxmzmL6co5fl/Mxuh6IK8cXLJ8elq7RzoasIe1
poE4qbY9aBC78+BpBKpwfY2TdzZ0rJmrUBlqb5FCFIGbwqBgjVSxUddeiTdtMI+EGesSLVMntpWb
Ol/ZlGE09vtUe5gwwwz8Ad3wV2sMdWP9suQj3hmN52w/Egos66L7sb/3ZTYXEHO4U8So3zHJQuam
VLnlIVM2UR8/gKh5Vni472BRI7onyJOcKEVuutwEHBsjay8yToS3axbkjtPTL48kvoNm86zrSPVt
tILRfKL3wWpgxfq6Ayfwxk4CBjg6q0GDYFbRc0gt/BlYIlQixzpIa+u4KcL60hIigTxH0fn9aIRf
3SK7XuIZbU2jY87Tm19OM6ZVT/bwBz/8qEN76fZZZcm/VNo3RrapRmoLBukU+7Kgm2Cbb02kItts
pT+e4eP1GZcKrdNpARQpAPjoadspFSeAqz+VxV598boqySJJKK3PuC6qCNcko3H0++e2sTIqCaxO
42gxNf1zZkl+2KcbqkD8IrSWKJuuPpRPWLYaXUjXhq2WagFtm2xXvHoDa3GE2vyYT3dqxe0KS4WI
eMTf923us0BuMKgqj/27suyVR+7xlo79Y6AMGKmqt6I1RM0xX3KSvKIUSjf8T8EtMG5jXpbRBUWV
0TWqpho7WXgb73s5Npbg15UPoMppuzGbi2IgI2ZFknVEMZvybiAskYlnni9t+D3vFSWKmGHAJQgW
vdVB7tSqwAk1P6XZ1ljnmR8m0/KLFDGJEAZ/jZJnAzJ3/Q2jvuGITIbMGf1y1DyNKpHY4+hF3TZH
iPp+gu58zLkrmwK/YY+6yJ/z2wr8DyLF693KVQVc74joSvATZfqjiDPmZlovBr+Ed1k0phVWKSkz
MmNqHGJnmt/vYMwJEaQPk1sz1PBq+7jpPw7hdaH1flInnbYqVZLhOXuB3iC4UyQ3eBaP5CFJgkw0
HrNZ/J6OLtzWTn3uH24eteJXntmNsEv7FrZO2T3jErjNIE30RId6ZWq32diB0Wbb0xlmhvsIJPkr
gbuJA2MdJcPQYF3AR1X6fIvjH6J2WrIhyim05SgM/Iel1ia/Mz3Fpc8YYOfMUY2pT23R2XuPLNtp
O/wxyVqierdESW58zpX/TXABOUcMdvP6BPAZzOfmIYT6EF2fDnWGW2H4ZcsfqmJkU17dWXEecekZ
a4ywLBXwW2lBjVRdpP75T2cmzRcKiHJDgmubJAyLwAOVOQTl8biJ3vCrnZKf2aD5U+JXt+fKbeAj
dYdzQdQbTaIgoscnPGKrDELMwMIKd+fVkw9WHAMhPrWUaonOiWbIbqXtzd4K+6PVBz/FBscgb3hK
wJ+1ErA/Vjh2C0Y9nyHFRct8KAhUbZxAanajpTez2kKvnwSd713BbJypPF8DmsnhnS6gU+MaUaDO
dBzfU3HHjwq2Yo1aP7f2eazEjHXk3ppiCV+PNXAEU6s6VotUMsGPhS7/tWjvvCdLrZHZaQyacs+G
D6+QnJJ3CXp99AtWL1Li0x6JDwzIA5TE1TZqiL+I5vXU8R8fNJGfT1/Czj5Jm07N4YC3/+1KZoVp
72ALlqrGdhvc7co7wkfE8iYTlV2LPNYiJiAnwenQUcg7G/+dVfMjpc8V/j6oRkLmvPupholKWIyE
6STrhW3OA2fJReFglRs50S0HgSQdIwP5IfSMzA3m3Zx5FvG35i6K//PT6k0uDbkOTMYR0DTc/64O
0uIrHR5sIhtNrrcxxeNjSP9ZaqmrbZGACnSGLIX2uPLkJ7+dYtvsaZOOFa6fSYkKdpbLTV7q/1b/
NiUsFUSIvrKbcGrRBibb3xBLyOXxhQ6+XrLVV7vIugjrcgm4qgWwRZrprq0Pf7P8bpazTTBGkYbZ
Sn9496YisedtMkbnREyudTpvfShSmsiBe/kEyRG9Df7FHXsB8t1CNGGmfSlSQxkOVg369TlhHwYi
Ah0FNmPTEp+gUHvtsBPy6p7QB6BRpuIL6M+/QDr5iNvS01Tu9cbtAqv5ihCmrwn30SCp07aUSaI1
YoAZvBUu2CLMs8jB1zJDtmBn4J4F1ZOAikN1AIJLOZB/A79yzduL3PTtyj8dMzE/MiinRsRUCxmq
WrSFVYH9pxsZc1A5b5tSQtCPSvGzqor/SWeJKsdcZb5bTM8FzPVfTsCf0h674pE9DozAbejZVBhs
0H1QegAeuQBCATESbRmVKoI5mj6dmKwyW3Wg1GDKFIoU4aAGJk48i+Z4uR9Cql87shJnfdaUq1SD
XMCQrMxcDXxTld9YYGNDbkLwvy8ZvGWXTksPxhZDwG2d49n8Pq5uaUlda7gDkUtQrWirlDjFybOD
E1hurfaeY9UNDEur0724CLKyIqrCElLlKQ1kIb9sU7kug3BFE1yIRQtJZnHvhXbzUMUE+hF/duaf
5kD56Js04mir/0mxLg9Pf7GGXgOfgeNEdmIru/654Q6wCVtkqs8EdEo6U3VwBK7cppgYvJUdPLG7
Kc/lLq96KsRf2gxsZKCQUs1T+zdvHb8m6EL+ljohS64PxTTI6Fsx9Nbb9VkIUhPwtMFIpDEk+4AN
gjQTTDFLds83zc9T1xsDggS9YXaOoGC8z6OSSqrwY57I1P80Ll/6MSoCCQsmtu7CbL+7OeCnOib7
BlkDr9P8nsSyJruYTeigeDkWnKNv+5H0LPA98Oco3kQS3gFYTrA1Ey+gBGUjaRb2ddSB/kAe+9jg
1r89/TgFXXnPbqbZPt0losMwxxTtK9iEgBpXA1HzMITaU0br2dL4Y94vban14xP9slDDREfawjCT
YEVcHzBs/9U8DYVI4gaE2gYcy/HKNcTPnlXeAik/bcM7I2Io3IMrKWctRn9moMkNSrsugnXHM+Fd
LjRlTpR/714tAMO4DDTYdc4g8JPgh3O8gKHUz9xLgefCJ7vb6j44HkodhVhZAKQwiQGBvwWGAlXq
MHBuddbB6AOBp4ypl0G228yeh1TE1+W9YqIp19NcNv867DKbnNZTbk5WAuia1e2OPYJSIN3kqHVs
l9GhQn6QcKSNrOhCbTUl7mossmY5X95qNABw6ois3JgRAloJkKUNTIbj2G8AfRx9RtrZDjUvMyYu
1WWBWrliafGEGxyPddAZyCbn9Iz9YmM77Cy5AZ4/Ujq+Wy7zQ4KYIWO6w5Qq4QcO8d8qGkPImnR9
pT0muLuguuh6uLKG+yUEm6mEGz5sZGG3RnhpdztAT3OA+feLD5fHKZpY7mBEHfqAgxZRccblNBss
/a75WdnaEGkq7sTcBKt1r8BPLaDqaul6Qpmrwg23r/Io0t81ZCrvJ2wpkMkjI3lDTb01UaUlH8Rd
euwd57LWN/llajvf1dxQnzIB28e1mKnsZU9vsMM0szL3eH54x2eOQ1c3/Mw7tulsOs7KI63lPQEv
Lg9iWXYT4MWbd5gMSSWL8JdC3RTvJXwrgUX5O6xTs/OqTERJf9JjAg9FS4ZFa14f1P0/0I+0JNeZ
YhNdV7XJHRnQiaVhTMg1JwyOFUzPqLPtHAihR7fU6TB351XFm3BN9UrJuR5rQpi9Hz+TJfvQ5gLm
82F3WHg1PnGs2IRRx/ASuHEfkiKVpdQhBgqQzoBdjg/FiEo+8CJ54qyu9180z8xeSTX02a8CMLa5
qwJo/0sYHP4CUJ2nAZ4VumK9rZ3UnUxpbABuMJkSdKBW7WCtqAt4ERyDTlHkD1MdfaOKLV4Ll751
TlPkvOMy1Q21+EmuxhiEq7eAE06WSlhZKAhdI3LglwKl7B8aajL13soXMYi1ZPWbI8wYa++ibDEp
CmOVI40YbFHrv651AWUDaLaFtRKOpL0NDvYCAm7UY0QpVmGD9qB6/bRUyGUsIC0EmMvQMxOpML8P
W3C+4DShgrah2hVmb+oswtTcHhZgfAdAjDiQngI5AyGubzq8Lm9QQwgsiwPuLoYGTZnMSPz4ixH1
9u4YG/yBoNWtogrx+fHpDtZEXc4QB/TuGcJyY/pEv3ImnXagA5awpDPEgwMjlNYa3rxwKb79zvfp
UVz1KzoKLRWUMlPe72uBstCBoFEBgR1KN/Byt8HEsKFgkIIYKNL8PGxI0T8+nEw87JUOL/SYeda8
Y3If7ld0CA2Fvzl8epknhEOWyPdjdbc+HWQgQUIpZXYsRvlO4X11lx3dsDhjGoGyDyCFBlyhnpBF
ezjZDtsXqLQIFm/6sJhojH7BhkpESVBURtUun7VGY+lnHGLYYIJbqLpU3jv8aMfAwLiBUdrJfQPm
yMW6nzp4js/8DH7XokBKnUDBerTq+JFm/Iw1Eaa7H8c4scDKjorVPDBorqaMH/Boyc07lwX6s0/L
ENbmYzUz80VmfYpTxyMaVgzkKt6TxmnHyvIQqiEUGs6IRVrLCM++1jmDdFsQdn6mosNxAlI8/5Mc
AxdF1hHasuSPnWxFMVC8HW7Wi9H1rurkbG4oaKRDtt6peBYfpHC5UOZvgVA+1TQsv2xciZ6JqPqm
k+49GvOppDlPs2iOq1C+XPhTRQfDxpM3OWb0ld7a+pjblcPNh7yzE6sdAhjbGRE8/Hbtflo5jEJ5
3j/KkoCTzaQlaCTsb90jMTOo0m0DsrkoT6DedQY9GrfgVBTJOGtMWOEy5tDbo4K3uUr/WN8IAMvg
R4c+14ePpKhJxSeE2N0rDsA7owiwDgSn0EWz9o3xc14kaSpPvqytrAQeJA/aDBRUzi+IGHSOX0O2
1wkNqUsIxeEDIS4r1HH/qAZcyqVJMN2FqEV40shXm6UtFtn/HhR0tGLOVjm7rE9ZMnskTfxMxSJV
ex9psFdtwIGaDQHrkn1RIw4+oFszeV2qPHG9cHQtushbdKtBal9qSGZltRqfs5FJp4F+VfUgHFuI
Kw1QypnDryZiLT6ngKorfIkiQXwZOKqLfqzo0Hf6+vjFWeXO4NjUZ/pbT+d9Nr1PGES8lDzR2+1h
WQ/F0hMdrt8oa+jwp27tSLGu/yWuMGUClyCXI78HiCshD1hJnwKqIUobHH2GqXuvCkEPYRmGEvJL
Pzb8LMA5T0dMgUW1xgUeyOPBngmEDQVt5jAqbiI//dzTZKc6hoTP7O8bLknBYsqwfH9PE1hnpVpc
nItDaC+kFhxEt/wgPpH3wUb3uVJy06X9YTUJ9Dmmse3AijbJsz4MTZjB41RjGvajSRyktIRJDzGG
yvMJAEMnDjPAUG1rRARlXfNseoXDibhuRidpu9Sz4NNaSoezBHL4/tE97Gzb0gO9+7rlp3IcTr//
YNuhQwe6/g2q2Pli3zBxBTJ3B7Fi5O7yJY3fWCgNoW6vw8oG65+Bi+dtMmNq/sk7oF5802GxiC9H
XTEPHGpQQh+RUGrQDCozEUDUbaZ4/cqMQPn7Lpj0ZYEoOWcXaQRP3ebrgtda7HWOlR9ifBVIUCSm
KVltyqK8qq0t/wnNMrEZ1MTdFF95j+Qo8SdVpgyQN5f0yGOwRlmkdN2b/9GKI1OOSSPzaZdT66Ot
gZNrjRohsgw5/kSQtWyNWR9h5qHciDJbo3R8zbWixzkX2YJzoJQ8oLswR6lGQKdpAV3R0qK8dIDv
FkszjL3G7wnG87NzKxJJ+5kyaXSCoO8VrZq82xK26nx9+FtqOQ4Sz5iEl/PbEahFtbJrv3orSu2t
xB4ZyHPn8zyq5G19XfvbZVm0WGBy3W3yDeW7VShYY6NMFmO+BALbnd3wD4Elk0GPU7GW0rR40W8S
CybSxaHUwl70kQ+R4rGldddFROSh4n/G148amqqmVVmhMTiWUQQqYaRh9lXpEjMVQiYCi4Iz77Kn
2esabvQFhM/tjC32/pDPLsrca9Tq506JydfAnVtyorCzZvMlSZLptt/8baPhmlPElz1vjSA4+6Z8
2McKHEh5TzQRP0jGCIb/t2bd2UXxaZLdHMHhq2Sit3Kco8c0IbBvWWVDdxNDTH9zwTyDWLMq37jC
3boT+K8us1oc7Y19xnz1sLFBpMt0U0kSa0oejKP5qEmKZKWtVZKilInKVCg+pYMl7mgJzcyoaxqB
mw38qKGZwI1y3s7J5ALO8ebH+g9SUmAzAjFrZhrz9suFyF1NVcXa83U9kPSDBP1N2vF8JiE7c2Vh
N2dWOBTIlrjQKeeS2ZEv1z4HKHawjhLVIR8g+uq+tiS71IVc0uGT1ckCH0pFE7mA8hjcTZnmExC6
pLzUtdXr0ZrcYCUrOivC/RJqF0W93RY/FbWJ9SPg/sHwWMkNslSYOUWhVtaP2dcjzGVl+eo7l+u+
leeWStI8dO4Nt6lL575k985emP+8d7EJd6JaMfmPHaC2Kg06L2SbnXKKfILuxOZmix3ZT9mwRKIX
hz1ST7Rt+lNWeDCOGDNIYY2ZTH35QwRTvXzKFicbBSr7+eFVeynjtB4cGohMv6OX01AlhGjSXTqS
8CIc1W+6UNNQiqMr2Ukqvc9bhHzocPxvXqyJ99ndHF0ES7qyCBbAZC6L6IKgFSNTEdJ5aibpgQml
3R4CAfxUZo6ZnjPZOotacp/wCoRox+VimcVE88qi19ArF4NTTeUDIcFrC0Bx4qKCKCvkM3IBp7Yd
Ll9e2vcIrysz5B8kxwaFO5c+34oTbr+5hG/wkz6T46vj5bJhlSGt3+RzbEofIHLZQaZ328VuvcsW
yNsojjMm9Hng12mNoyI+LcqkI87o6bedi7fO8WjUjzzY/5pEv+mStpUS6sDCQm6lXDp3Qm11uAl2
2dNTDc0FgmFSixfWNVmMr6WQsY5uGK+LS0PranDm+MjkeJOZPQuh5QGajzAZ2EvgW6Ia4yhQrzuv
t6XBo12mxv1dcoeYR/RTkuan4NG6m14SBHC9mvYGXDNtZNhACKl8tcngBIjYSBZCbyBvMeO/p6SE
wnlsOAhMmoA/w0WuF8cp/5TlUFrWbWkrFnOyfy7F9ahqJ4nQqZ7xCZ3JVw2D4lnxKWsqF9pGToSl
i+9+9B7vDkkBkQ7wd78GBUQV7Khv0fOUtohar2oHeY0cHb5/tX697pF5yjYr6jSLFvXHHRDudHcN
GTLdU+d4HHQiGRXi+YGmp1r/g8B+SO/LopJi1+sk7t4eUaEEXJC/UjFx+5AwxitdUA824c2gPEHX
ULOt5rnP1lhQQA8NwuO5pPaOvr1ZrMJebgNDMEoe87QctT1SpMHx5AeQqwaKjwOQnFScuLs2eBRh
El45irFsTEtcx2zzypgWDkOIsbC8g+1gN7N4y0DVuMKXjubtSLOMv0VW3+l5MXExziorWYrO9EcH
StkLyw+ROfKv90gVbtqacS/SBwRVtjvTxf2ytEYcUFZj4jvUEmxT8cNqz9g8iyUl8X3X6t0nghzy
/CHRVGW+ZC6k75q60/Nd+er1WVPF30ZB8/83rFM117PhM6zDVUEfC7uU2dGfObqevibKJhy+C5P0
TV0hzEuPpKSOvlImc+/11qiklhK3Pd+e3sFQH4ZS7x+2MmS9kN5nkM+X7wOd7Q+2PifhehxvbDdi
8g9majubBaenAAGnBAitAXSxvkf/m51Srah/aRyGH2gJA+Rc828uMgyTXS4/WzDLDBxsFl+fzls6
j2hbFG2s0ZewqaLcF4HsH8nYc3S4RHJG6jIEF/Rb5hmUiKGud5+MPkbkBBvUoYxwE7wwUpCCfi33
O9+LVaf65ccfjIlnAq9gB1Q5z1XzD/evwuSWhWTAmM00OA5e9Sqp1pCEd/avL/xh+uqxgcIsPhDl
A7z39W1bbqE/xJMI0QLVrKfRfi7PoN45cnVNv3LSB+6K95ZHK35UWnDg02EHPuKOPk2jg2zoXmi0
OjgbTXmErfq+SRcJhp8xOTTL6Ax1Jy+5kjNJiRxBspqerB8wjYCe4KQDjiOymvx459MJmpkxsWGK
GvQqG8Wq5r23o37997A2hAPaSdSpa7uytN+tyTNl9Z3dUyINeMHZl4/Uttq6F4Z41ReQ4/cV+leT
/JZhiiP3BycF4SeB0iLR7tsQpNtKAsRAJDTEcgoR1CVlmgH1qytu62wccnsQuRzCB8MUqc5MmK72
dCTnk9SiUHTO1XEmoE79vwq5AtvR2hQ8RxZ6xDaJVjR1tPKENHtm5TXTy8WNdZIjsUB5/8EUL+vu
Jdfqf5Sz7oXaRJXNaUJnlWziFlwi1wasfmPKXRXMXHa0dHF8RiTXsCyC0GBJVzIXCZZJ/Qm3NYaR
yHAAINpVIeySg4Mf/P/wAs5MfopBZEBl6U3tvF3rW9YSSgyqCxxJdgdPVlz0JZT/RCYhdEXqR3yn
cgTneFbfxWGGC09VsSpCZZjkIEHU2K+Q5RHq42Ca+Sm13h676+ErrOM3RKhiZqkmCVDnEMVmiGuM
cb+Vyj09uQfE9no/7QS+OX59a2Lzcuoi3XsHAtp+BCT16kX2vdMezyiFNJ57sQXQuJ6p+4iEyyIc
r6w1wXU+CY6Z1qipU4oG2on+eyzMmPQBooFk2CNSg2NtX0B6gLsoKCsdy+lAwiUm2XN30o/i67Pm
mZDN9MXEEQOW7LYUX8x49+0z0lO39YJYWwA1MRt80z8DU+W5A8pUe3+K2bvlISZ1oypuM68hIPAB
kWg22LeKNsyeDAnTOJDCcflRu6pO+PZeYBwVXAlpjqCbqx6mPiW8nX8YFqWcubB2lnWPiMoZddac
fUD/4UWMxTCZ3+SQGTL2aP9KyDOu61CE2EzYcd7BBvGGrHtsaAkO24AmJ4FTN5rSNdMBfavVEL3k
rYyF1tL13NXVroCFsopSQxsgd75KCviw6u1Tcwv5nf7yIbo5dc8c/lZy9snCZv4l253HJqrOCdnj
8NnbfzvzF3//t3p4IWUHt4PrYBIpccqkLxm721vssZslmDGZ+wLXEefNRVdtzwU+vFVFkB5+6Amj
X2hFKbsbPBOhTjX69oSa/yqVzhocXfgHpqEavSQkzXb2icAa04sJhGP39htbeJlgZb8UWCLC/ois
PaBsongW/SoyldAS94CE5DTdhC9IJfxScl0Kn3un4xXFaJbr7jS+XCfDAI8586G4HXqTDU6mjZFg
jjGHi0fOWrGPL4D/phC7eg8O/GiPGREtpNWCt/6U4TGiRhG2RYFJ/NwfO3inrBqzM7QgvpQLVkOo
+ojYi/GdvhiYbeBejseq9VgIt6BO+dST6w5LLJHqczZc0F/E88vGC3StIveExYByE1btXaVZmHoz
rTVDtDVP9X+5kf2jdAktKtdOpDxEpLqIAIXtOXWmwCqZEXAxJpx2gSMPmLTi3sj9I8HeuqLWFqY3
78vc/+gZJ34ITzc2mBA1jGD/jRbzVmRWC1CxbylqOd4hq7Plo2tvEQ0mJA4w1wKTfwglaWM+y5Il
YqcHjTbnOBJfbhUc2+LJiAbF6qmjUYA7kFGHjL/omhi8S+YMtFf1GgJZ67kbw3BGi1dpC4Cewq+W
xx4wbsTLSDRg0f3NZoZIHMZ4TZFe2Fi8tQxtq5vgboIKC71uNRqhSb/s2sjS1VBDEQddoPxq6CSi
V5bpml8bqD6GxenNUWF38H7qNmFLCtw2KnciWu2kkF8gH+IfFssUH3cN1gd+ML5iB3NiS2UhtlcY
2sUc0YVNB2KiYiguaMRqpG5QCvj5lXBHzd8iRLMw/u4NNhEx6B1TyvJ5oJK6tr9U8Qjak8wxclRx
Y4Vio5wGug3iAOxcAJ4LDJJ5+kxNwha3byaFzyu69vlc68hNp7agu+zbwEKz8Dcqoaxjd6ZFLaaH
0gyqZlc6KkvPe4kLBqL5bpidXAGC9ycVlbtBVTfLgPeIev9izIRBQ9+HjWB6WKbSITDn9LFjdkH+
gxdIELPoqzYknUMxFH+OXkklxIUEipkSkHEqfjTKrDPo6+hIrPuJixITuxePJ6J5vb03qzFfT/yN
8JaoVZQPkQCWRhG9Ihl+ojzqO6rl2CxHmNZJGqzRcW50hJSxKiV5GHpQMDyj5xsbz6CfgaasRdku
s2wjDMvSdVL567tTBP5sb0VOKi+7O1WK+ZRp5RbVuUxZNslYMo706Jou/2+5ub3+B1YTIydtzrKo
rpiN+OBm2ryzDaOOf57sde23+uLBYWUhfG2ZQP1E2vbx1U0toHY3nDn9wWITg1gTOKKHEJ/cc53c
Y7+I/+KS2eFGJy8G7Hn41W1tIbYZD/N0iccgZGIvZOTaRJ7yV8dB4BmUbjIbzfUx22OYYHA0XX3q
XFeix5L8rOZmWEj7aB9SDnI/NzNAJrrw1rnRLb/VhS5xzrxCJYCEtC/A/3s1x/FHsA8pRi2xEq/F
GnPAtC4LZ8tCpt+e74IW874Uzc1/11Qh5YXZ9rESfT3Njjf0Y8xi677mtpqD+iWal1j9adhfJbar
1W2NFze/I+kn1/M79bWrzm4D81FK5avkcvGt+tEMLQb8EVY4Y4bAdXCP2zOzU+xabpx+KL5WIZ7L
psVFZykmS/rdX6jNlle1mqGFpcHXmCxMgbu1oSfflzAIm3728RFfadUNE0uApZu5sWYQtvWGZJjf
LRmae36iyH5emCw5PSLsfYGf3jMcl2HNPc58tXeAoZuGdi+xQZo4NJBM2aN+wd5YhXlIJkoBAbCM
oI9eJ+wXYDpjzcGO2C8yb9X1LVrxqrbKddGnJjyCW/0UCT0baYv0fZQOXLiMDsEozjtVPk3Ipyez
XxLug77c+sBrxJBJGqnEUCOY7Zcy6GnymRYj5NZjIOqELGeGi1mTgWT1RKh7iYq/QkEHl9phyBAN
Ug9w81I0TZGbFIn+7w9wd0J9csvO2Qk2l9hk83ZaIZdnh7vAt2+zqIRQrirIYjRZ32hKt89aTyvJ
/rVze2EJ9qAOeHMF1S7F7tycd8iZbrYj49kItLq8YU6xDLIYuGoR7xSnK2Gi8jKGfCkt+MPu55Z+
1UnNmydmyDBnEfPDXk18GTyZaVap03RjQkBUbgGaWFFnrJN7wysPF7R4GdB9yU5Dil27TweDd5tS
N04LSHEWoCI6zpRWzuPFyLdINUeGnamf6easZIRv+UJDI3SI01sS8Vd4QNmsbN3/aWmtsEMzUBzM
a6L0p0qqJBoebNMCfsZRLbG8H4gcXyEEjgOmQYk+cCN1NiI3gP3eI1LujsFdwFQ8eKaKZf8qC+ZG
wTgVutlATONUwGxRD1tvuhbrJs1WcFdPAJyK87/l6ZFD71o9SwGvazUqBne+qIuyjcduxmjuk/Mm
Gf7m6xl2GoO6Hycgbz2EcIHQQmGnlHOmCj+3BiKYLApKt8aHEQ402lYJN6NYJPPBumwZEWHyePjX
c7GolUEH2n+r8PkySmL8blYABHIE6HMhN/xUr/UKs1rRGMX9roPgnLiMVrojsenWyrKmHjsSewBb
wFkZq9BY/ZslyDMKvTgFOSpXX6MtMdkHVKHZJINkVj5vqAwkocYlzEAiXaUQpzGpXJFny4X86twi
0+CjnsyTIy3+5FgpT/Hrgs3NwYqbQGZB9wPjgQdcQRjgqEmVZPyN7eOdREDlnrhWrJcwP5gpSSlC
lKvbSIfu29/t6dXO/0RgfB+zhrvEymY8xFYrHTK7us1LPEPXa6WlS12zXXwniSmkIZKv1+1aHAi+
fRWozHLAinbAHPJo4CC9zaFxj41kW3X7f3InQ2g5Erflb7nO2J4KHVx/9XExE6Y3yjUqj4MFYOB7
Qc1UrMDCaJuDOy7aJaZr8c28RLQkyKQdXLJ28esdQqYWsEcEeg9svK/P5bm+rJbXLKvX4FZ/S43/
AHhw4wsNsU3tBMQsSz2favSCyhhApGeIiM43Mc5QAVxRiNzGt3/MBBKmn7N92AKTAZj2IR0THAVI
LFUJxsx2DFvx6WDMoCOHjVABR4JRW9Pzar4WZJCK9w99xm1Uyh2IORP+68LHnOGU3b0ZoC5ygZmS
NeBUqsnB8xwJxDllMG6k9Zt15mD7LdmnkWWujQM8zV/23D5X+/mzVWYbcnln1Wz/FZULGqfu/fh5
T5spLqAmkzwvUMdNHJvZKljW+YFc4IfnzAxrlGSr89nZ8tx5NqUCka03KPBAu8zerpfwJDePInZK
B3tPKFM/fbKcmJWJuEZ1IYBvBDeTNkustgms+q8ojujYEfgKcb1W2iOZeOrBv6JObBTUx13RdmV4
qOZYxfcq9yoxKgzaBEahuQxZ9p4fEY7gH/sG2IsenpwDwBqGtg4oD00at8b1oTmaSEbFVd2Upm6G
91XMWDANrPvi0uh+yYfgW4kugNOV3xk9tQ5PbunvZM21gZpgW9S1ilMBCWlxiQl9wSTd29E2ipzR
DZim4FY45VTv1YeKB3fm20On6Ex/LGvo4QKiWqA2BaXdb0ohzQyG4eNREJ8EBzvLBwA7C1mj7rnv
9AJ268pBwXH6vpEK41X5R2NgT5GrAhRb59Ojb5WYE9t09//fUQC0NmmvoFBcim6JzJmmjMDlKT6m
GgpAE/qHXAV89s/eGoH/xmtRY8RjIFB+623ou+MHLOv9sbFmw+5Lp+E+sLLUtI/0MnVkLL0WYj6c
PVe1WlpscOW/c8p5zURmH5c7riZ5snKmYOta1Hj4OHjRpxpJOGPw97EocQwVXv5HQj0f0lhQF5PB
e/pYC/L2D1J1/u/+FWtUtmvexvhnfnzVxEnETOfSMWCqAuDZRZq1kEm09trAoS1o0g5ksXBfJvL0
wNLvKqga3+GZAB/FVcthLAtfL8Mz1iySDfRL+PNkn6lTmjF2JTmJn6J/KxqzzE5vO7z5W2/t6+UQ
j6mQEioe6EyCKtptE74qN+v41MVBHnt6tpGlxUeNPAf91tLg7Ug94UqJzc1aEbx6boMLkg/YLCOn
nqMoEe5OqlRIBa2gHWx5GNG8q6ZZc7CocAbAcKdql2yWC/y1lFV2rfCfbdxD5mcdon0a37ZdkNyj
utTjIm3SvhBmLuKoXDHYAVDzqA67nvS2vBjhkxHGQI5ng1ueoUzdTo7D6KlCm84GR+v8sVnk1a3E
ynRpIGkdjUgFhz25mds8Q+jnlYVey0vOGSQEFrzGFfvB39lW1MgyAarVtmgJ6i2cm913FEaU9Aui
/CJSrehNcR7oRv/DNT1N8wE40fKi5/VZcvyJnJ5NHULb/XTAHL17/wpvZp8vzPgQ8F0ia38K8JA8
GmRCv0acOwo4GdIaoSWLgRURSvFRwsU8AmtUKc+XK3nSvsV1768+thm9ncIoyYVKOb1Y3W+EL4T/
JwRHg3s9CcKSoDDVBrAN4ioVd3PVqsHznyNKcB5Lau0qPSX6o1SwalEsbH4SXF/7rTzFvw2KPc/y
6rAjD9jPiFKPMpRP+j62U1PjamNq7c1FDUdMBzq62uDW46krhvaSg1ky48E0PxIktp2YsVGX0HCc
ME6kpC5A7yP0zVDoI9nJOQCrK9ixdCMLKqJ6ehm6/k61l9gTBHPBL6qToHLFn+E/NCdPG4Cqi88I
jfhE/mVvIpsk5qCMijbBySYDSsWgGxjJWwbN0Qb52vKvfHn9WuV9oVw30BdbxSx5cpgBmmqY+BkS
ZCyAaZsvUFhVNoEl2/NmGhnHU3ywAEMu7XLuF8rN2bKpB0R4hdDyCpn3lf3XBrQHqpVziI+xed3K
UPBm3UynzmN6Kebe5PVZzI0KN4cB5vJCE6WkGwvv0mNPuP+k7gKPmQ1XoJifMRTK6serNYsJyc4l
iYlWkKJVNrnpqsS1QdLUS5lcQbF0CZksmLxXPHs6mV0u/+UNWxsNEeowObS3SBw/0D9mHRaTvzHD
fYcqDGmxJIjKAhseGwLRsE7S+e5Lii/4ffkqr2flgychnr4aIORKoM0WpIq4yRdi3REI0D9G2Ofr
DQCQZskFcw+9B0b6ImUrwrmy+VC2W0KVaNVKLudRbwPFvQdVyY6iAogJn12WNWt+Kk8OEs511Df4
imIlSuaUAqlSqfdLa5NrgSdV0RtVuQt054no8BIMem/MoFDSUhNpG2bDa8a0u9bcSHbv1jGB0ivJ
YKO1lMUigJgQzmTTmPkkzjM18CCdfdSZLkkupHGDGj8mUi+ckns9zFhxNTBmIUSePYddluToaNju
3Z8i57+rpXbS1TiBmk19slMxFVkRBg/MZ/pNuDXx8AIO36wb1b8mU2Ap1HN878mrwUkX8sKjIFHj
srJIZVVOGfHjBXgEi5qBQvPwmnvTbP3vvVK6jgRWM8XHuhAK1c8zRQjU4v7YuasvYAzPZ4HIy9m5
JF+CbZfgo+rOhRTf2YeMYlFxfcq8EyOQU2kyTl6HZCxxjTNK0A9jg+nMINXUmDx4yPP6zSJK/hrU
RVW4APJQEvowy8XQC2QSfXAfk2OW6U8TODX+DtuSKJUGj7xg7deTdOGoTlM3DGqJFFT0TUiwzvqe
3YoHatLMdJBWSAM0uZdSqnRBhHgpSQqBNXdTrGxwBJ7oNAZ+Jdb65Anzo6A5dsi12nZOPLENlXMH
c3KYKmiq+HRKneRNMeh79SAQpYWRf5ISYmbnr+gJA1kQCTgh9/oLmrHj/d5kY+a0ZzcM7RWroH6M
sWUqg8VnL54bgQr3E66ZClp23hJy0nxOHFyKJQi7o2TPjBEk1JIL+1tElfrrHvPeLNHfiryC01Mz
UI3aD6owlgDN0+/v8RV9Kh4uW+f0Q8/PKhmMWI6GE9e+igDDmgh9VcuB5G9XoRsuQW3fo4FlMrWX
yKf41Yo6u9RAyVg+FJaDzhJ/R9TsOR5/yEPRA2KB1EyZ9jZE9MfR+JscMy5/9ERXfw2TgXfv3T8P
OkzFbRHNJhngxc4fKjwofgXyttVbhRGWc6IBRibbngVOBZSqreUdiPX+/nCqKxKV4IdNL1FNhhvj
MG657R0OkCf5GgjvDJ6GbWI7dpxQ/nX22XcUpFhCwGJUaU4zcU4rdOIexfDSxa3Orxy9/cboDMxe
+PW5CfJo6oztKE6W0N0j2esHi8V+D7Rh622eUWOtt8+48S1heiCFnMq/lNvsHSBebCKaRLzLejIv
hN/e42zAH/Y6GYckc0hby0HNEHA4l8iymMTbAoUc7LZ5MtLrfg7ajpT4S20tH41niyCatiArFq+N
nB0lOj1YvhrXGoz3I2YCyuzt9NXhy3DMSJGgaIDvjRfqYmfDsL32UoCVyqO9GrFpEaeBjxrUMPgC
hkGfKKdM0jz/hcoxRltuShHZNq9zR6AAmgui4CHehW3XAZE/YS9CPykIqs4whMej5g6D8y8eUazD
Yiw3TsY1w/FjKunoMXtafzCFX6GIWwU3BHLsBkvD5ldvF66f2ka7Sh+koqeLuHiWGh+Ug0MpBxjQ
+D//a27TVTSfJS7DxIUufjdMpyevxwDFP7y0lQg24B8q42Zof57KMlotr/kV2G5H2GFZMz/FYTgA
EuRghY9GnC4xrs2b2Zxv6vGT2x3hQIWQ9H3uZMHeiT5SWRKwbqz263hHge/Kt/wZkolhiEtt7vmk
uF4TEfH5lAC1HyFZ+jFQ+hjp4YfFdUJII+jsg0Si7UxRQpi+ZB+k2V3ceWI9uMGmAnIk3pdMfR6K
12r4UzE+W739/fsK6NZCq3dUeeY7O/bU1djt+IjFdoYFuP1C1C1X9FcDG7DcM6lJ0dT5eVY86EAv
ACyzEHp5jwB22bjszOcNmM1rdW42fIvqWHd1D65qI98LXf4ljFWdQzdea8Jjjj55xm3BZf2q2LJd
B3qxMyQFR4HpbHp5Je/rrtbcPnEx5XPcn5PWa14L6dQSa5F+1ANwYJ/eSSreVbNKuYQjxIke/gUe
RhOztJYzM0kxYH9oIyGmMUNX1zZnPMsBEk26s6PsxtNPgLTRcy1tz9zgEcQNZBoptJ+VTZvvNzZa
t8/hQoEmve1DxNDANQDUbIGuP2n83lK5cURxMl+UlcYXD7XgiN2IovZvOSTgKuw7orHM7A2GNSxl
nbNW4yXslEHiN/rTcpgoTWJoaeXMFR227HW7VrJtW4ZITCK24BbcNrruXgfEHUb8uzs+PsdQDuZ1
BPHWPmW7Pw+wjc3rXEcrIjz/iHd4OJYiXuoQexnDTgdsfW/RtEz4EJKSeFZKn05bdlhkdrkUO+5A
IGg5+zZceBDq5ej9JGOtJ+qFrHewd1WQsWnIZDuXPxv6c27uSVvoeHunqgfEGuKpVETOxC76Q9QC
0zwO3hLDJdZcFxgsSRaaUz2DLw5hbfHXu/8Mt9+OCOZ8CIQbUuwppEv5lmj2LucGz0YzgP8L4Cug
/5VHn0RWAFeQ1XtRU+jtHHA6J2GbAR4aBBoJvpts3+oV5K6+QV+rKpnoicHgLigByCPB7KwAQmEX
goxSuV0+8kZfVIMDRok/sFtQd3L1gtaulEUhWLVIVLInDBRsA049iQRcvPdxKC3h+Sf/OPzQVnBu
YWvYFgn2LvazprPNmCmj0tfTlH2T+5UhSNCj0xWir96que4eQ8IrJ0+pxh5eBa9+kcX/CZbAcABO
iZ9xd70TGBNW9dRxihw7jDyGcl6XTssh6KVp6KnYD6jfVs+PT5/gcX/D0/3R/qfsk5Ny/XAbCWT1
lP/e+b4vhpekmPsU92Mf/x1tB+CJuyD0J3kY34RlfZ1gNIbGsm86r+hA8dzS5YhQM6oDZ2eMRWbi
3UuxDJ3GuIflPy2X14wPM3fUhiYa+q2wK77LoB1Zkb4sA23a0PRqjHqahEyu/5xjkjPBcGFviLOd
Lm/4As7BOFvXAzjw4f6IZZqW7OFXWQ4ondU6SFnes9jgPSBmIIynn3EHICXs5Zjvt6LBpJvISvp1
Fk/46J7ZpmlYA+fRJJuieXlD3cixvtJcbWQ/i/kGVX7e2Z35t50B6a+zB4U+nqGM5EybsaolrUxX
6pckU3javoJKXwflJLNFIMfLuq4J1LErVbZjnlhccpmDZHCxutW1zHcQoDpe/6h1d2NjW6xU0u8Y
b+Mbp8Q00PnsEwvof4kryAAFNVOoy52QDRAC+B8kOPoAN4HOJSA4DtAfaVO9JAsBldbseF7dGBiy
hQf3+UA2mBxENbPYCW/OlBr8j7egtd4oJUFpfVPX8kPsgtaw2qZ3kNao4S/pIJaf7etXo+qJ9gy5
sqCbqiOWPNi9REzXi/BvxSWKSZaN01xYOFYrvAm/5SZdy649mcgdyeoSCb0tFqne6VydsgXATJTU
rIvVy/K9bXxCKgM4Tcbh/wEiYdDO6llfV/DcDt48XrwH5zFj8Bw4JvwomEib9XsmDAnjjoQO8AO+
H8FW3nCJyB4A19SpVvkN7YP/3jfyVS5ZBs+c++i2lGn+ttZDFSyZikXy0w2pTsBEYMG+LdxRgVii
WsTmqZ+MZ/1NorOw21ZZfFza5aNfZsjJhDNIKnnbJ5gG46Gh1BnSKoh8iB/MkMddY15MDXNE4yM4
bQIp3ggOLSquYz7BgvCTw4txWF1/SUDE/5/rURXh6laUV/5m/y/0awNcIIIYIe0AxM6fnFfyxHce
6LCO2K7L+LftbPM1WESb/otw3HVIQTXgWOAUgO2yIOaNKGp0isUno3ZQ8brAt8T58FlxOUU/s69B
4rXoV2R2j4uaUlC7sVHxfmwth7LOZQE5ZDjHowe2Ke+fs5XXrBua0tpqk02tg9m9mGGETtXnhHp5
i19FBrZp3QZqQqfcynTVbCUUw+ZLMsCZVDR76UX3NG/pav8vGb0L1m0vVDPZh6Q4EP+skd7KQTHZ
gg7nGN0gC43DFASqt2yCPQ5JeTpwu1TgnK2xUoXSJivHQ1F4VIrGRynqLi+nzCxkJWkVS/0Mj3dt
q3S9U5TOO2z/2lZy7Q7lpak86z2E/JJyS+zZIlglcvh34+3QWaHsYX4Yu3JRTxtY8JUQ3LiH3wi2
x7YaV83omXyxDhIwjHbzO1X5uXRAlGJITuH4ZiTYqOi0VoXXig7vdVDH73iPAsfA/cKeDyC6Li0a
Xl/rlNPAxzT49ADaHmrtcmkc+WMKgIXxYeu96S7o+py0qMFkiNJvomcskqcqyYb2n2ZFU6Ty4OdB
N/mo0f0pE0H906YRPXanSSoiL0++QCL+X869aTW4y+ssX/HO1a7CS175q1Ws21FX4EtCm1DP2snV
sH+d9PoTh7Ksh24uhUarAkj3s943Hwv2rAUwdnC0nyGz19NWQ7E49zo+bPtFjw+ccvGdK2X5sj8M
cVabvVvCYHnF3HLfNSdVyK0JxzNjjrAtB7erFQ08Mvt4dRftcOjS8YINQnKzWpmioMsmRLXUn2Ty
w37ijhBRAiwK84jEZxtsIOp0BtRgE/BG1aCIE7CQCAr4BNTCznc6z0DmBqyT13NTMU550TdKQUGf
vy9cMTtUzJfkXtoJNzXLvO0aBhWSR3kcAlUN/cGFKH5XB1nzd7azyMl7F5mxaKYu8soe+bHC31dT
EN5BywBTYzKK+l9HQ8XP+XkLNcQR9DdO/FBOxsvai9QxbZjux5kCdr9vRdfMeEoMdGDwPVv6c7au
FlfNMXaFFldbD0dwg3Ia3r80LD87MJOBLS0A0fY1RxsAwPIMhhtdhlP50mtlnlfefU9oRgAxXc9d
ITMuPKzz5Iqd/l/zR8pYfjw+cTuFd1b15/fOm/UtTXtCCzkPzMN6wtG+nJKBkZ1CTKg3ZOBcKWK/
sxYqhhKo40gVhhG3l/BK9bF2CG/sfgtA0oH02Ik4dQmljtrIOPDeWo+hjXlsnUIO+1RsqQH2h0vR
HJuJGNAPbrCH8a6pfqXwergkaDCbDSfjwyfMneIglLYkL4uY7jhBsAJBA0LQyoRv6DwnrRAkUrKx
PewlsWEZSUzrN+yNkyXCowiLxTWst8haPph4vdnQHjtdwD/fSv8jjomPq1WWHURUeGlp789GohSy
nFG4THANsH7n2Brw1IAsZp+ZDf5HskAF/jKPw2m5/XFDE4lOUO+B3b8loxKP/TwZxVNSZa3EzB7t
0jHzhL6eUeaJKy9TDDKQUFCr6XaZx/+HNv+Cq1S+HJXCVXo6whoAJb8YRSYfY1gBZ9b/wwcaG5AI
QymxcP9uIAktQ1d06iZnfHQdB3xNrJyeSJd+HM5m5TDRq2Tz/8LVw4DZAaV6aNrltL14gS1BzE2w
7dQ3czVW7innK/+GfEDcE98dEfWvi57z/+tvKUK4farmUHJVhMUIrm1fQUKB4NK5wo6gWFAeUssc
E1vnVlNVsLe9YA4eA2SCNx2DUPuX6TlKA5Ywb40V+FupOCUAseIjRQYNqZECUC3Ddx3kAvHwIjd4
TVUfTSrq+jDDA3jG/X7ircLvxBFpk0uw6h1s7Gda0n4+n1IyexUynEY+nJZQEH9rJfaYd7epLTxh
TSJvL0/ekG8bt5ofFofbV2gZay0+F6x7qZsEecI6OZBc2FFcbgR97rUm/IR6kItsmHSroUUXZ0vJ
bEgIujRdpTXpUZHuBZEwH09KCt4w6yZ+FBxvx9r2/dePmKLfAyGmeOaiZxrNb2Lv7pi2C/8/wUVh
3rLkIsbAs3WE7kJ25OX7DvNUugAbkT7BVIxttsOsODhonSHgb6p1ku85WufRY5LvsWdnqaSDp6yV
dl+6ZEHevk/KcfcDwABXpgZlk0l5F3TCnDMErK8Y6s+iObBKye2H/aF+n3whn+gOtcpEGV38kuAO
2JNeCbicBtObsN55DhYuL+GxFkIthDCaLLiH5bS3DCz+pjej5vb3j7fwDrcuc4/ARPZOykmNWxGL
teq+NvZCDbTi8ueaNFu1ST5WuJN4BYYVNOV2tUxq6QWL0Xjmle6E9OVH+IXhJ5Ztn5skR48ZnYgz
tTEmUuTbZYPS0iM3FT/j3FVboGF5iZi+Ew5WDJZMCsDr4PJ1g7aqvXM2Kiwi+Qj3qij36pb6CMiN
UufikigKRgaymNy92jIrDRyyF7Jz1cyKYvuKhX1IYkUUmXgIdPjGQseA7NAReY40gsLFkF9bWa7u
8SjO29/LqKQn9q53lV/+e9tBkUBD7HRtOkcSBd5n5xbN4O9LV+ckGCPexlL96WKalDD/xhjNsZLv
CLrDDELaCK8QxIU7ZDU7aL0yklaXG233ec18o7m80hh8ci7U6RjjaShSoj8Asp7Gi2y7ijzsNan+
RE68/qbtU9CBK6EVnqu/lmYZCsMKinrKYRKixcqBXyElY5r21o4W1+Iz4syTDKcf40f0GYwuqzZk
H0MUFgRfSlR8K8YuHEXLeVNHb905BUXg0QTHxgt5SgFWdT8a4wrGbcFpx2GNYhW6nz/M1uYJUUuY
S9f71BrmP2aVnQDl5Ztv0tDecXabY68/T/jRkIYQQiJG/198zB6iCd/B0VTmTSxRJCWPZZqYtSeF
bbgApgWLGhYPBMVMDJOaap3bHF4QtapXkrkHJR9rYJhJv+AIicon0HucumUlbWf4+8AF32fjgb96
mlZ79rJHRTA4UCfAYLumyl4jTNd8jHGD0rIZVyeH1aFQYEBLKtxkooe32yhTm12MzgaW0B27N8gu
Z1oD7R59A1XOfY9Z+PqF2uGUKk+AFDGPDCNsehYt0s06svcuT/03e/rfmAU+MiX3/3SbRogRy4rk
cusVpcbUl1ci2JeXcIo/Em/RsVBQ3fAY/99KBcu31DprHF4KtB9Cq453Q/HxKjJe8Ks/meqhfFKh
/6oZHbbB3kEUUgUJYuibTNgDAhukvEHHOUcFUjnDCwXavo6jitI7SJrlTStfZLS2RcJc2pSFp+w1
0mmNVZ70XylrygLD8gyrL6SgQDRpo+DbR7QJJxDbhnsPZmtlNt+K7gSuEWyhdja18OnAtPm/liyX
IqzS4CYknixeRuqj+O3vqkYcnzuXAbm931N1e/QJMtCwdngOt4kWuqHYNxNNcHBPPN7dbENNK9/E
8U5QX0WAjS7+GRBA3Aj7QIfpiYmuU/xbozARf0p70EWzPR3UmdPiDkaag2xnrhqJZrVDzF9aIrEI
Fe4tidmAto6IyyEB0lZtXgxf+lrijKQU/cpI5Ker9CkavBEwHaBN81EE4kcu/O9CZvEFUf1dAqP2
/PALmSIDrHb/WUEkK43D/0p5f+2I2rS/G6mgOz2dKuvISBmMZsBWTFeKXOv7xBNJuIAFx7rFvAST
6homtV0tPwIGqJxZ21RafWZfeA4GHC3QJl8XBpzm9s8yZ+kdSbSiiBf5mnm/kXfWORxZgA9m6r8J
xY8oOAlC5R2fDh9GaFMYjbN99+9jupb3Qz/yci++SaKS/rKoYkOq3x1jU2yyWSAaB3N+5udcrNCj
Jn09M/z5tGCUOZGo4uLOu0z9j3x3lQRPiqC+MdmeewUti4M9t6LSlyxJz8cGUab+b3BYxz+hOdq5
NB41SEPHPH8zpe3mfV+BwWAqNmXXpl31Rxl+B3vtwoa7Zbw/Ho+ee6LpBFAyIn8O1tX+8DsMxFDZ
cX6SHU7HxTZFGZGmOGvd9sFhr4iH36nYl66O9qjLepMOsUnjShHjlXEiCHCcZ6WUkpj/oupYEewk
AVJOwZu7Of3j8+I+P72J9LUhQ4I9xIYdDmPoOz5c5z86jxUO1vrdejLgymlaOyxBr4HoZ0cCs7ht
46I06ifZ9d7m1T9rWdNfB2NkB1V4XzZsLR2RDlIfwqLLEgQm2mxb8iHrwk8LRL16UP4U0A4ABWWg
xqFEwn3E2AfmHB65GQN/MGu69JpoZeTb4kiTSTfwmgQQ/E/ArTsa/LC/hUvwkHkedADbThfaNujx
V2vrqWvDNeEmeNpJtxRWWh+gxC8Mk4KCMQeiV2GU1RV48+fbkv/FJ8kESqfJiwCCm3qH4gwuee9i
9ZumAxzHq0Z6sM3/aRBuNzR7q2OLoMtCy9Oj/X/pT0yV0X1faVvetZZO6GHoJwUA7FyV40cqupI4
y6pP1XsSrakD/RXCBmrN78ZM/9aTADWGInuumZOwoDK48PZHZ3nzBKx6Run9Nzc+1wx3lGJ6Tlpy
l5tINrBmG5dWG/D5hK6ssaBVIn9cIWmEmiqlgCTSS/uE+lGatQ5cL84c2q+ZeISIJt8aX7QOSgUs
MlXfJ6Y/KvZiycprtmDhgPG0mWqA939RSPhFs4abMOGVI9XvVn3YvS49mhzj8G3jLMRcwc6TUClN
TPw43717o2ca4J76Bls0rT01pxOs+snVIFDEkiY4hfR+HU5n6GoHQiDnk+sQknunD7oZ5UDX/NAe
IwtmrUpzDM6/uWNkgbo1eEEI3UUc53WO/1ev4jACKdeZwFeZ5kj1BDHSb8axEouJ+Q+x9uFa9kjX
kRo7z+NrcbEy0DkK4l/uHzlpvwicV30B74A5jziU/RvUsqmgG3gbu2xAPjjUKBEpajQagl+N8EpB
HZGHH6ebd8Kc8vwcLY8QqXkTg6HRoZn3JcVch9UiRcAJcPDF4/MN/MBzqtF1wL6i5oOpjGEPbED4
tZPq4/ahQP8mK9BMYfuJceqE8H040oQ/BbEzM/xAYilpHXWxpZ9TPOLFuKVj7wC96zyKjZPm+/S1
ehDSKpHaE04Ea+EbXrfuA2lMdbiXU/AfBcRy1eBTMH4gwm3ae/DaRR+ygvET+UUTuexQmiKz/vMw
FzSl9okqigP5h+Rvtx2No2UPEvglfPfh2np2AXb4uhZPSNDne/r7hiYbJhckvMGNIPY2WxUZB+Kz
EhQsziAcAlZWIO7ZpenyK/8X6xLUriQ3TbBhPEBlM8CQJ3+9wj7hkMkOGpIJ3Rx34HccceZ+Id5F
oDsVITZd0uro1SmOGlCjJHiG1Kswa4vXR3i1lR+EXXESO/cHLI2RdhuUnv+mrJLLvpgw3mN2Kf+K
p4JmHHMqtgtuBrAHYOpDlmyQweED0xprixLvSdXv2CHonAYpLBQ3A5pKvxUm0vbY5VEADcJGSWlZ
OpGY07Ojnz9qCC+JeOOHWvy3qTsFZJytxK3WMnfRS8YM+h33/LL5Xf3Lxd5D8cmVbtZM/2oh2Wbf
4L69lVjw+RANWNtDdzfkEB21QGC6MC58Hx50fiT5Ed2zGINoDupVUITr9i4pVuK/BOxoumPtdOl3
M8OYh3s7BzaRlDpjLSbsTSsspws4J/QtSLXM70ounITGCQVxuTlVktHUWxHfIb/ZR/kRYkANaRgQ
cjE73IDor/OPoDFg+DMfoImyIHwPOhoU9JL6ixBPL5vZ68JfjkMrwuI/naJln6dIcL7Rzsx97zFs
2KTX+gAOkdql9v1BR+Ds2CJn3Uj41DvPxclVsyhDvgPxhxCKlssCWGk724F+IcWlAkAE9yVWK13z
qto7YfUzEZ+GNN8DbeY3xiPSaa6cQ68Q3vzoPzAhSv+v23f9gYW5lOIxPTRM5D31HyYQxFYor+cv
reh01AA2+zfZZCz9mSjwRTcs0NdrchiDLz3rIWPeI3E20rLwjHt7niSZfPN1TGyg6pRrpka0fzvB
e2nPhLev+zrisuHBKNPlsV0f10sJjeXHfWdhone8jK0UKBiw3vX4tH1xYA6KQsazOimwLyMIBkuL
+0ps2V+4EzzM3x38R17J7ZPm1kO+AnDOZlyY9V+wjMTBFu7Zt3f1b75Y4JOZIGskfRCWGf/WPBh6
w/x4FzJI1Z6cbrIE1hd1vSXBxO1brjVXuGcvytd30+mBg26aQhe1ScZKapT68UIZBFcMuIKcLCy/
cjqAbAVe1q2znpVA3YjjuEQSmEPzywmSMDMya2j6glBU1y8g2e5GpGlwystl3JZXy/7Pbaq3lpaU
iVAR10ueyNcm8w3kSAsuBBIT8W5HofMp4Obf07/yxMcRRu4HAl2QJqp5QCy21tQEEP2yq2U9nrYz
ONrAT1giLuflHm8s/tVS+hhLPP5ldLxVfD8AogmzpSt8Dqd8pEsjYxz2fwlB4cN+cx5wSIzP3a3d
AJy+2BxbbOjX6e5wQy5rWQl8LJidsKUkXa8HkBqPw9OuT8WkE3ZIQhDdRDq3Z6y09b2tDJkfE1fB
hZG73NqD/120lUjqoI4jHfGQeDIaWexTHz9+U2eSa4iyd7piIQ1oJathBULBLET2HF9Md+774Kzi
K9dNat2cORf/vO7/Z486eht8x7CsVEYhHtUQCBgOJYQaOfMa+br5GmT83L1H16XepMUb5M+b4Yw/
b5S33vbSpJy409RgUDuA2M6Qj46asoGj1ht5YrgZnzsHwx2L0kC9WerlnCoYfcOibQJ0PxVNj1Rp
xSEmu+/5teqFs3ECQN7yVMBRpYjhQ9z7m/WEpZZqptstZi/SLHosx8M37gDBqiTTNcciRdoPsd6O
/AR+nNw07g+xw5AuPDDKfauKn/ketGMoAebQ6h1PolGWbpn25XVlthPx98A3gbSzCJbSMamaSEID
HLDwzOKwi2Py7EEPk8do8TYcOrlSGBROQpjLWDecaGNg+KCbZhC2ZcGH2pKgNTluZn3uo7jp6clX
h3wFtBkcRtNxzv/y8NR2M96i9ZsnjtPlcDVeEgHnh2qZFuOxT7ei81dwUrzP2RcG8jRIvv9CHaYv
tCbxzF9eCCNdSMOR2IpkXrRWQMU4tX41sFFBicAFCKrh3GfW9CKAFDK/lsW8OrRxFui6gTtoN3+X
9KKO4MOi8fHTJfgu/7EwBVdrjGa96XvZ0VJ9SSHxZuHKZx9fZzuEeKsrMj4gibs0Ut2rfSrJ5dxQ
f+SdZmtoZJdTJ7mkkXHSy7SIh3HisDQItMBxYYStQ6xkUgRGQ+WKgGJi21el+8UfZfVe3Mpum8m8
g+tKSrx7FGSg7luR7/zfpQyZamcod1V7EYPBMK5oWQWft8/x+baMy7BFwUlq+wQIMF568xguBCEr
vlbT+pXzAELUvlHEagKVsccvzdbTBUT3vl1MwdZjgj99Q+OX/TaNsRcv34Bpa4xauhFlH2899y9K
3y0/aNlP8PiizANZzJHe2G++zr6ghRfoOlyVagdB5oY1+8eaXJsE9furDQBChdzhf/PNf5O/euqi
rnqTum9VkSLUFK1DFBrVpOErZjYXerHk9pTSzQrz5EvvRhkrxJ0j9pHXw8obzXUT0w/bwgXd0w0m
tWMC+h68rD/1Fu+8sSFzir5B5nb8pmN32rptLrWtBLw6TnC29DcK3VmXMlQacw3lPwm1eEepdtRk
6jQ9KOQHAwuLsHRsRdrqWTyZAXMFse2Y1yUV/YA2YgRlgvzgSBjbj78if+uaxh1w3yPjHJgfbdVF
JKV2zC5jAw1aIwXAuhex8vqpvSuDayCGX3qn1KUcdSxbSTzkeLA2DC3MKJgzuvhGHJ1pRxev4eDp
DcV2+Dlj3a07LL32xeLzl+3kWZQdJi7NTnSMT8SBHJj9mQRW4EouDp74VUhF643GkDHeAVx+y6LD
XEKT5+QZ4vgsoTO0W6fr/xeHJh2WifXXi7wbmjck1ykSPeJK6/kz2qS5fJBPBNhXdDt6fSl9H6Yw
nqYNEBnFwBqpGq1hN0lIaIi+uSDLH6FHzCVC9EIBM9oswaRMth4qpE+/f4VsiH7uhEJLNpiX4mxo
IFJHRoSUJMtoTX9T/QVTxxdodTdDM3tJHsmaWLxTjhj4SvtC6m67CbyhdjOHWYOrt8tAdTL9j6pl
kpU76vyBZm5dvbbWIfmrnYqVryqgOjuqgCcJHb/zdjq+TMroydPMWFXLnpkPzv7D+E0w/yB3ixwH
3UUl91rmJFBAZ2r8REjNqK5bqEaaA8hoAxpjUjGhg/a/+lSEflxzmLwsk4GEmGLhZl4bHp90wcgM
WlE9bTxd2IrVTG1I1KjPrB2oiyzvGruuf4TjzZo8OGUJai+6LDHaPRi+hdzEX+UZ/eVYNyL1L9ew
Gx7Qzk6mByXZwUPJGTHtSZvcrIAYMlEkvAmDkh3mss+GPVoVoybCpMF2YQ5N5tgvtkLfYaeW/Tfd
YYJA2F+qOch/O2ct9CkOQZbx/Oswfd2XCGIq/t7YC3ji85IzJCTZrvRpDAL9RpOqPU6F8bFikONM
YasjJb/KnqphGlpN9aSPe6qO9EM6LVzq4sgIu3zf1VuOotzEpttiBpaigjGsehzqpnxfdZjY0YT0
qUNJtNxu4RnzXrUmdT2FEvYXDbHYhS0As0XdnLhLlKz/cjhUBuLs5Op7bBW+S2foj2IBr0e8YMl4
hJNKF0kuDpIjKF+hCnzdQByfISuwoj4982uM6CHPILUEzFlNL2fKPXBke1r6DbDVybvN9LyAFeqc
5eVsYcvRwqEmBle7AFGlI2FUUqO4LiR3HVwXC/VbOSLVWYt3RihGuoNDaTzY3qQI/FjlSpxC/jl5
+JczZ6CTTwQ4++PY1Hrxu7OCQlZWY3r/xphYD7GkJkE6AMxOzhrng8G3ASSCoMSm52pE6W+nI1df
A3QqSN5JeCQOlDcRrD3+cogppJMetVTRSvQcWqBN+23sfipuKPzCLNnaAsJZX9TYP1ndRhEtqTTv
a9ubauM+FAJJPrZAq4lNN6sDKvBvnZIlPmPdutH4bFzjqY9oV7F1beV5LHipXnSd3kRTOcUCNfmo
zhcovVWJ5N1LQAmFxq20znigZLYqscW5/+2GA/+UYNZAg+ZJF/HNc3IJNbkPxt09j+CrZ3JWNiWG
v6/DZMtyg5X59d2Oc4R1+ZO1Afswo0ZhIq5Ts7BCWxdbFGYL/B5Zh90VX6BpyR/FpLHcaWzKLXWO
DEmlR55lUMTl01M/idlATcvbFcyHuaYEXTkwcxBGkD8fzxYKAUQAsKyPUPW/syXXA9D3BZu4tOkP
SX+k7dHe/j6m9D1uyrXp1RH3/qY+sKNpAKcLrntja+bOQM1oBrmMPToapY+rPzmt8ChSEJMZOYcR
XxlS1ldSFNfYU3Aa0m0eaEzh7EvLg1Yt5vzUBLYXRMojQJEfY/mNgpQDidqB2A827EyRLlpz4ykC
CfKp0o66+mGtxUaEdB6pjTt5470M5CbCmb06ooOEcnCaAawuvDp/PQf9yKJRZvbTMcRNr1oaUK8w
9Z0+NSiXtrVd/svABciYwO2RRvYWAr2ToZTqP7+0RwG53SkhwGwOn86MZudBotLjkLY/CKqILA6z
tz/LFttlJlBiMPIzH555DgT1jzZ9sO4Q6ufisAm4U/o3m3W62vZQ/xWS8+V0eYgccL1T8KVKapCp
GCT2M6a42pP58eX9WseKApv98w66X3d5TACU7Fh/kibBrz15/XWcwwh+M4G2BhA04jvGlZnJ2xHX
nZzNQSSS1cfQ40OabBuzVxo/HFbPbmZtOO426PRKV2Jp68JeRfd9QQgsGtQ5qqn/xe01OKJrAXKc
TwIEWaamelRmzU762qkMKAIky+Kq/1/60oThSEZkoqFOqZkiFtcLyfDHD/xn5OIR4Ig8qOZsyHer
wzl8N5TyjzLEQsJXLOcrYrkaP5mLPF+bgtx8l4Y6/KVnG4NPLNS9HunhENL8iURS4RA6SNRJFShW
0ooVxfk5LNM46AkerjY8MynasWplN1AlJBDM6WYSpbFU+sUvUyd5FsJmpoNCelEN0KzwB8MZqFcY
SDWep85lLGj9YSQWIkBo9m1r1dGfEKdT8hHNL08D07t09g4zpWJmPAZxvs+3r7PAWGdNH93Jgk53
VueNRKO4F9h8DtU33xPgCc01QvjQ+1zdHYNxWohVc/XkRLjipr96iwh70MI2lGDZYBZmCcPqHU7g
h/E0JFK7RXU8EijIskL+VTCpa57Fz2RNEB4JIZVYvBPujqeySSPdd8xRhSnpK/5lulvYi005yjyy
EgATY7Kdm6RMSuRMbL1aPwbrmBLO9u6/a7ZZa6XBxZmoyXsrKbHYrPWLIN77SXUuIzIEswh1B+/8
VYxX/9L3JrM/VSM5JzFILp/jAxKsitMH2+eO/kg+MxSOaCBd93rRPAwd1ILfVcpPLhB1BXH7ga+a
wxBFzHzEF8QeLSBvI4y4isHImAkzQMW6EHCeQaEBhTUSYy5mZXWcwuiXjsMjVxgjr4bjyGfu5MU6
33EwwC/iI4EIlwkp+D0bYWiIISD5H+XO3l4Y5ieGLQmDG9X0gqy09/Kg33W6BUyWtmqyIwzkMIZE
jWdWUtTUK+BbHV4LM/OIFwaHZgsndzleZprCdprb++g1rssbHjhZMeyFtMK7GJ8WN1b+yLJ2XASu
SPfI0SXSgXxanQjI5y+F+BpmwzM/g5SvSd8gPIO9vnu/CfZfZT44t+n3kshtP2T5nY7d4uVnTTFT
5O0HoYk8jcm0f3WbThNIZIgXRv6rhuickciEfAOmNJ0ZrisTrvfSandMkYuzwnCAGORegHmVdM6d
zdaQppeA6H5xzkTEyd8k8G41ClDHSopfBDjiF7uqIGDRE2Q/XkaH4wRilqsf25AUBv9vJNsaAadc
IHIHlaq9gJdM64xWIBUPEzs3bBFNnyKM6sdpMdIvmpcFYi3z5A1J97ONSf9SI90pacBuTkL9aGHR
ya/AUt4sL3sefR2RQDQviSqphLgG+sS4SOuzz5VPfkS4yfsZECXQgHPo948m1eOLq7vxxSAODHlw
Rt1PseogIuB4O7FyDY44uymduGKCHE9b4EvgpWz5hvHqbBcGNIk+PZhDYfzAxlw4tBNLMuy/BWGX
J7A0wbNuZ9ILRHn1vynmR2FzQFBbpxAJ+34qn75pRy/vO8C4wGIAel72bZ79dsGIPjhTCjdKpkXX
BatsfngZSC72xLfZIQ2SyzO0L84I9eNdnbozC9iN6syS8ZWGROH9PfHauFyoCkjg8Yi7srQgEqWc
PhLhtcfAOoJQfqF4ISct89VxXh0lj4zysH/PnNGrG8HrLxCyzJhb+Fp6PSWEDxTNce9tNgpwPn8b
gMskY9oOWc8y23NTuLZCSw7V+BQRodd6eTNkwx2ivZ3dYdHYc0HwCln6NFlR0Yoys+/KlShyxc7X
YmNKD//LKmaVrrtqv5qy2Xun0jsC/WTSrBlSD3B1D+h5UFRy8UlfwkiUnUvMFDoDu/r1uEy9xGg8
GMKQKLsJSuhl+3cy6SE3Drc3DQU+GpRArzuIdnLCNNLVQ8NdkgTT5tGqnwr+Sw++68k9dzuSqKjI
tVW7JHmbaR+uiRfSU0SudRD9/WRX4yELq1xSw7xPHgRhAOonh/nYQvT4DllnMk8ON0Jnuy6IN5jv
gLKE2U25+Xwe4eKUK+VSRCToz+jmnJKe+VNOWV9RPed4uUgGm5keRXNMiEqY+HBIhOe0JZ95gO6G
TGBNDBwzNUt6cDJlsk/GRhBvX7UsnLm80N+RiX+WgCjT1jiLwuBwExC24tnV/lQYcPITrp6EDBSm
YkjFee4mHg9yWO23/LQroelS8bGMYob79bHl9raYwjeJEG+zopoq+32z35IuBlgDZGl3P/GxIelL
2pnyPgVIMDrJZ4jrKBsBfBbjFw40I2UpW1ySqjk6CCnSe2b9TIuID/ux24VUyuvv5mSkf2rKAn+G
i033bH0ntyFNdR7VGRSyJ5Gdr2KoU9j/VDS6jDvXyEUS1H/exikiU/ERwYLRuB3/BcKjUwIABJr5
NnsK6R5U2RaTgR3e93cMD1xwvurQ0r7FsDuFxNC9c6uhVOBFNW4lYCshdy3f2yvbqNvd+xb24zno
d4IjN+MIFihuztXoWSgr8U6Ez/b7uhOOzgu4nxWhMpX0ZusuBtF3T0HJZjJZ0iB1dDjWFMNgMeZx
Nik6uJAk+Mto+yqNq5g4dsS7eQWlC7qVIR80f8Ah375OqfQloLX4NxU8Pyc/cFxZoaEoL59SgclJ
4TGMXrSv3Eh+PcHrRafHYBrxJiNwbIpCC+X9jBgUZmNiB4MZkZx5uqZUkOusobPQMzn3D8brFWAj
6cp+41CR6iGCqR+sFr5iScUAvP23RJRtdme4pajI7fBPE2Ehp28/AMvUIGZmGNGxaKP2XUgV7ij2
kAZsaAbZMBanxfMJGDah3C1tO0IIZtt/CG+oeEhKwl71gH/Lf63ncz6DcARtWk6pH6p4A+p4mTLI
FpqzlZz3MVm9aJIbS+wGbq1jacPpnaGsF0G4U6VEdQ0e8Ty78BSqabb1lF8r31wKixVlxJXFe9jm
cgygkoU8uzoaR4Wey1Sc3Ry6xLu2Fp1nh+GKEYI83zqunwWUPIk8CsVC1TBQ2wkCnt2rybY2C0kL
L1cl/fqMMuxaFQpnH1LOMHZF4XoIixuOthNWf6HQhL4s6LKBMlnRK6Au394czLVN/+Cuua1glX3j
TMoer0OrBMYbUufMcKIoRr9oz7ZTuMA49u+U/wEI/d8ddA5x40n+aKdG65ZRdgjAiOEJe2g0ww45
XVvnGVNKqqjeoXaQbgkQr6GJ30HUWEND8xVlGPhBuMNBWQvhmfY6vchkn1AzcFHG4v8AhP0/Q+ic
1wuiwhnMK+yDMkZPGgccD/BZZ00Ew1oP7MzZAaYwRiMVSf4bYlIz+VeV557Fe5tYXWwmM7ygFmBb
h/5zGsKns2lDr8oIQCX7BE2MfWwPmB3Za8J8AF7CMnR0uCM7LEvogEJ1VM1wuSYsNwUIe/qBwWuQ
gndIQqQuHR8R/RzVA9NQsyAPsPA2GMo0/djnt5mvAxA0LYA0b+4jcqXt8i57kbGr/FKo9PXjVl44
s9D8u6OZ6SbrVZL5u6ClOyANmj87quq14Uok/ZQ+LuP/fNgGRu6/CQ0WBaET5T74LAhj0rE0LAJ8
mydLH0sfgweYgcEXjq8zaLCa3GCbOemjflPZLbjvoCYmd7IhzEmF/sSoOL9K4glzBP2QV7DQ0ebT
fGm2KV3KZsoum/9X4/7EcoZzs+cSk16+Pd+jNqP29u4pirgJjXA/4SkoVh1I4t4iljW4tIXFmqrp
DN7DDhxowuDNWLJMBQm+qhgkgNqYSjM0NBAPCXpWnojB57DwF9xFaRPiABoLsUlAIPEh3FnwV7Mp
14DEIanuQ0NATz6kLLlyJoN6sX5egOPjUJenUqrgewpDJwvJhNk7EUVwzDxWwAW19f/NKiauKaGP
7aHHF4Vk9ClRr81jOws7eszcL1n8t4o4+fFibzf+tpZPHSrGdzdo6E8g4n89AhHznDbkceADftex
Nl5aMJdMUS0QOp2CVU7KRBFaHxzolXuSl6lXcQW8u8f3+lSk7licanPoz5LgtNzjyMQ1O5EidQgi
Vhp0z1ikuP297pQGs2l6Z9VzEqbeZhQa99yYLzVwOrvLfcN9yrbkwqwnLtUVp1J87j/57dNvr7tD
oozvzNfLPxbAId2rh3nCG/QY0aP4uyF4AVJ0AnyOPKt3VisEWqdtMCVlHW5QT6ajyzUw24sxwHJp
rowuLq3rcfz2mWqLpLlT2W5EeeQvkWNYQe63QoRZ/VNaKZwZNcW4bt8n4PFMJxvxhk92MWwdP93a
ao0r22qaBsPo04yduPLQcdWILxkDNWQgGw0YM6zfu1Gfpl6IriooHU0q1Q69bo3GF/+snIcROmen
OZ0pZemN74UPmg/e+7Xqi10mH1T/NnUedJiqksE1SxId+ofuP8E/zZ6hEB14RlR7BGkORXlbUHyh
PWUrgnCT7uDrUQbD/UW6ZWutlPQTmmMPUJ5MXgtfcZ0rP7CMGz3yDQk2SLJ8SB0fPydy+H+Jolps
jjnkuHZeJwpMgF/jx9nwcz7nd7H6mtQNX4fQ4Br12nGZ9K+n1irUm9LggbrQYJOGhsQWTJITV2AH
/FVicC9qX6XkAc/huWF7hpY5LQSp3k28F+dVnDJ02DEbOMrUeJWbg8iMX1XsT37443z8WjCnvgUi
sdX5FJR/7W2d6fVB6nyoN0Z+ticWy+wAc8GTmMgXLXiDXqlJDqC/V72pWc6hxXIS22tgZ+c6+pUZ
gMUF5k771AIloBDDpQs1/zSDIWXgaoszQ2N7TrSMkn5SFOvWespY9wfExXYOQXb0Y7Mb4xFTQcGq
zZWTELlkFmjA7VwxVB7VmwJ8ZfCEFqG9of+gknAyCeOgct8KtQa7TYl7jvbRRrLJN3xO4sJnfOQ/
32HdnkAy4BmfQrMuO+VyMIyPSqLKhBX+GbjG13HRPDx+WXsXFOxadcTM5nsAYq3m1bvIcuyNDmAz
sHXGH5zITDoN3xbxm+4+XGZTIM9736sL49j2LoFfaRTc5bPbTugvFv5rnuMn9DYJIEUdFuMbxoDh
GQMo4rGNHl3bNhfPi+Ma5zNVqFXGjq/3Vz2FN6tdTPEKYZUUxDM7Y40l00Cb8Qr1A8JiNash6mb0
5MHyzYKcXrjn0q/UZI3PWlGuXZn3bIQXygHG7QSvuKbCkwyqUJfvacv7KXjA8+0IV5VyAV8ud6Pk
r8J9z8loSC4TCyfnOXzzILPAQZgSdC+iO8sT0MI7x0S8DzmdYv+/lFuvu+SVN8Ayc3tjSD9kAqXR
37azAdp2Wpk874LSCqSoOYmhnM3FmHYpR2T9gNHnU7nUnkUeZsnS6/jz8+zvr42zFsOdpq8u7n6L
k6yLy9MDglZaX/CMwkTBWLFG+a+L7VajVd4bqldRxNPTV+ex4p70/DfB/57m154/4UCLllbOe28K
/rtE7/fyPxGOvRnepFOIeZi9nP0+ZQ7Lbn3wOr2JGiZzPHxUJHJ+hTS5Mb6yZNlJvZrq35GuSxaN
TNyaoSHiDmFi+03ZThkyWyBzoSczRnbNq0NYHkM98zWjWPPUo9vt733VAoTuc97PWhqKeq0DhZzW
p7gYQ8KvhRU20ApwJE7jFF/rMuzn+g9kOllsTZ4cRZJTd5sBc6sHLXJbTDAvKL4xDHTrCmKxNAcF
+YdJlEqhw1fnLlqKrw9SnVj2xJ+80M/jdX2YfdpcHO4KevZV7bbWPWOA2JWb7Af77qQkMUFfJJgA
a89DKaDR/ybKGHQaJ78ZIrHGbR4aX6cV2Bj2PANNSbDuLF6jeLaF4lOTOVoxdNlp4zYUK41gRzcR
NVswZW7qrKq0TeiSs3DJcNI0pmAWxXJixy+v10BeRZfavw1E0py6u0d0nIl9KURNfoNfJDvEl4hH
zsY7tSoQ4AG+DqJhsLiZMhro97RjhHBx2/3K/N3w9XZrni6/8q7IrxnxvM/Yr3kf/pW6CZyKQiYd
vZbLACZqRL93fR98jduGIXvP4JPv9dgmQs3CK12gdClhfhHuBudgG2eRv46OzTs+1zmsLrMero8t
CLrO7nvzv1fliu+ziPJg3gQRwLEREkc+u7aCcaWzPVJEJi4kGiaRQRgdpstHu9dZ/GR1C7vKL2h7
l2BocxZZO9B/YLNR85nDkDomUtZL8V3J74DFAvXrW7rGPJ/LX+4ZILveW/1cLr3BA6RiKF+veNGY
zGU8957yM6l+8rF8Rud8cO7uWBvRynKws2yZ9rWJg6ynXBugjet8EKa4FV5FnUJH9U13Yd7MPBVQ
yntnwRVLPkdKMDUlusbOoVuey4Oi0wx0i9Ti8wtKswPwePCWHC2Hgbb2PUKq2Zwm4Z50A3mbaFcZ
gQYC+CoMBdksoM8DXcMzSgnwfRsHJg8lwEo8uyA6bfyOhr00MF7P6ZhqluqkEaqIF/PFEUC7KzCI
Mrct6seh5fhyYhy/8IjJ8ah0Rq9U3VwVXw4jKIN2UhOpCKK9vUZcTJqI7C99IEURVWOXsIfoPEWV
qfGwoFdzyQS2XAVY4iZ8viXSf0IIqXdTez85A4bCfsuy05iDieDEKtpetVZ8dIf9ORQJhkQEbO5J
n3pRA0rBX/Sa2tRKWoUxNF1ZSZyr6J3NcexYZEW01EBafl3Sc5NbG+XG3PgjUp0enAWD0gIN7gjG
ACU7duLJCxiRi5lsHzbWRf7Hypuq9e9CXWKT2XUX9NZFO35zuaq6mRaeLX9/LoJrfC0FUYO0ns18
63JtF4eOC5NXO3qq/JUnIM0y0aPI98L88cOssqCXx3VC+qRJj9mEKhj8PurtnLniS2GrGkvMJiao
Sj9+lHkJDmAv34yyDcZWNZS76+qZQu72ge7K0Jm8x0TMj4J7X8V9YnATYckgZs+sO1kHepHkhsKw
FKn/whtDcfSogn90meCvqNp2Hvo30NLSzngpEcDxpAV+RarXjD0soEXYvaPZxCMuWnCveNcDuJPP
8M+SN3173G/hKhaj92NyQys51y5BqGTVFkB+YDJgJpaLkJSSBN1kMEmjrhxMl59yRnUaCO3KyFVw
qGoID5YWXGIEnPjFunHtyD4x/yi/LHkfs5TTr+lNf3+pZHhamMxZcCSbgO4QEdV/7vlM9mL0qF3Z
QdHilkhnaQhzz2bOTD3qkQKFZ/Pmm9lbDAWbKL0q825Mct1ZX8V+mycozMctCdNNy7cr0pNkk2Mf
OmhGto6nWnKI79KgwTQeTR44NMrT4uZqyKiAqB69ccseZK9iTP/9ghYo6zW5bQhJ1pPMHL6V20Jf
ZHXZW+aS0rRTrlGsq4hEw8q0KK05Fq2u+Oald6AQhCMjt1oE01XIRKeVGhmXYYVv7TOb3qOtGHGX
JC3pV9NM3ay2cmsq24RzvUaGxcJSml9RpeaaPTwN5PZxLuX0jMA/RYu+TLsvna84NWFmT0fAjN3j
yf6wrHgvKmHvFov0SQ10fHOIj9mG6clD4uvLOPfRc1xgxCiAOX2Qa/QEuZ0U4jQfYxsD42FoxJoT
T28KhSnAx+LOAthI/o2JLRhAe2OAEsC21TVeO1uBSuQ7irkmcqxv5ORTKQeOuXqbdkkoq2gRCp66
hWWm7mIKVa+yk14wLU3UWSZqJWrSamlR3xuA9q8n8uUwr0n/ceW+7b51Rc3VqS4kSFlF60bWzi2w
et5d2IY4ySSu0oCtUqcN+20TQoaO1FweIpy1uouWXLz2d3pvUy1DqON0lLXfO0sAcHLa1YbpdN36
2czMfz7/s4LhcmMSIYJCsmbqncmfBOn277vwYUAp7KIJPB6fWnkSSmczdvx341TGZ3OPfVYGB3FV
tG7eRNZ/U01e9AZ/N3WLE0ZzYfstQqA1L1VV3jd75VRYpmqtPj5Miq3j2VsR9AMt3zkkACxLh22I
IpzamWMCSSLqpPaWuOz9CJHACUC8wY7MZLZgTkHkpzC3sH8+ZpvHNANWuLejpVxkkJxATsy9BW1E
epCOhZtmRo2dYhrMb0Kv7q9lcsGote/3+2ShGfyqcECrvuVEnV1HWnlPBi6ARn66fHvLzrU0BSW8
jlSE1McIJeOxjfWDc9SoVxlFG11ox8NVjcHFFPrSyhBE9EVWLPkoPqHnR8xXxCBaM0BBiZ2gNOcA
KQtw+bN47f/+L6Ma6cyuWiK+B84mqo3bkrjcaF2pTVWPousDN0zG+ZeWVXHjtrAk8kIAQImjNoHM
gqpp7QsJsCOVuIyAXcYtyl3x0AJ6CpTL+rEZx/WIg5UTADPQ2c6ETrAH++LZmBODojlv6ui/4d6q
rMpamfJrgPYe+rtU93rkoYMRzB2Q5Ssi8j3Rso/7/pzXNOxosN24RgbfQV2Nij5R15QtURoHIzLU
PlxnKdx1evvww9B04FAXBmHAC6uFGoJTjsijPUkxxYxbns9jUF//mojrzfn1R5udMhDZlOW+PMCV
66+gjq20mJ0luB1sASi6+hNJbCHjSSgMT6jzOsDIf67gzUWn+hFa1sM1mqaG94hWX01lPed64PRL
bapTJBc5vqHSyykz6ADrhbF+EzMzlgNqUnugGWB3Y3Fjb1QoDeezr6Ya1NkVyeqNqXD/06Vz2ox6
t0O+9LTPlIMTiXKGSrR7kOFL9NuPzx0MdffteAoM51ciytLLDq/wYEl0QUYwPJeqxSx4wI52CgT5
lgpyqzgBR1+0jbrPi5PBO7SnR5+Jh5X60jnToAQ/A5xwIB+ntCYB9ks5t4g+5GOyLYWWWJqvGROg
9UFiIleBIxmTcBWhw+GkLAsJj66RqG9GE8U7YthXTA/vDm7fUJkQgKLco4UKAl9BNaoD6OZi+9X8
gT0b2UOWAvQ93DcoN8UgHpKsytqYeC4URwstELTaKeMDJ8twkO3k7kFeU1fp8b6LPqNy123X+IIX
zzb37lLss67tKteEO/4q7TgS5hWVBulM5t8EH3XfebKv+oKYZptMcBRTL4Xuy4j485z3q/Etg9LT
iJHPM+NKka0ADb/phF9kZhip2f5JRKPnrC6N3sUn7JD1JLXh5hl+FQL3aqDnhgZZY56zKT4VZGSF
VJQFRe5sQc00YvSa1hOdPImWUpXKbm5QR60ppwLuk3DJEKSk5FYzZrwEtCXeWTjB2rd7rZR0SiVX
5a3njMnQA0so1l2ROmJVUq/nt77bEES0zQt5MEG1mjOvUW6fVrTNjRUlvgM2rJqavQuDHK1Bj8b2
7KXTAeCfZvoklvPcq4oHKNnWKa0yD0cMq3chvgYn8PCvj5IY3Lo4ELkSV5yFvuyXIja90Zyy+20/
tkdPiogWLrMP1d6NOZGP7Vp6aGZNQWm431BqAK3M9yJuwnsqoMSdevZYKmJ0SEoqPRBO88yx/SYE
lkxyYrRAgJe10gC9l16hQwiIBlu5GjManoWhg8X/j2QmstOz6seNm74PRrXGtL24UbXpv7t0xd8s
YsQKTCqPABXpJgbyaz1bIk3wrkRgEMvLYqydgu2QWvJ1IFe+Im7Oc2whS6C/HPB9f5rLcC96XNHC
imbFqXyivG3tDmDzlQBBZYDrEQ6DKnt0l03c8H0OaNLn9XuF2ZtQv6hMDSozg2CKMpqtVNQqXLdT
NNx5txz2DU+N95OkIupV7SHpGSPGBV1Z1NxbhaoIbc/PyqqXeXyzl6UfUEnWs8ZWw57ukDnmHc4S
yUxIvZCy4DqKeZ77fv7NcvHqn1se5pqEm3wSUjkL5+iSOP8q9FkljgmmC6dHt5YA/WleJAL1PSUH
OBGP/8X8uWrZHHZ0O4rci84okzf4pAG9DtoIfY3PvJk3azS6CwYVlukAZRvHxX/hs6pkVs/q87cL
L19wV97PTWgPMkNj81BY2bjyfDEZfzG5P2DTAD1MCKWfOC+IX6QyqYrrwK8XMl0B6nCr7ku0IL3y
m7bK3qdnIwNZuNFOAszGpWxEG9dZdyi9GE4r0u3R/b/q9moi9dNVGFhX5vyyKJiqIfLctEgTe/gl
i0Kx0jVOpTmBK5R8XXK4htwBg7+8IsX0LHHLEAZi3KYXXE7KGNZV1ATEXwWOKcNHhh35Y/xK2nCk
neSFlgxJv5KIDBmlYOVPzV+wNy1gtA8widltn3TAfvbMHKSF+y1tdrnuaG1VzvaFsFe8RBvNZFWb
LL0iLaOVfcVlgz9ac4m/qE1xlnojZLp4YMqYMluP3ugxCVvlh5yYRhQVdIwdCdTgesFKGvS9yrqM
ooTqXC9Fe3zLpFN8xAMAqVEmxlbt1mp4lGnnAAkhd+usxHHqPcNyqRQSBteU1ca/ld2m08P/IaSJ
SYfRYYtQN+kzJHWFVV2fZt3RQPPQZQlFz8iWR791+C2+M0ysxsCDuD/QKrGxgqs63TbqK894jZ8L
5rRGSpKuCFkVjjAOgNl5Rd32zjPCddMh3FMYdcsBNfajMHIXzhxshtkovYVD9Ej2m+xJVqJC1+ZE
WGOiSnhmspZ58Alh8H57Coi7FrUgozbu9T5vphL5swyiHWWh452FgX1gE4hzulcZptFvjqpyroO3
eN43XUe5x0CEMMZs1q8wtRXzcGQwFtRwu6Utp1vWr1prASGYhcJDKlVfLGuLza/ccy12PYyQ1BVL
lYQiRwcflnX1rOsTqd45tv3Pgl3tE4FMEYKLBM24Ta4gh3ePID6JHqxvTKTlV3mmJVw0KT/CQnhO
QnmuBF/vi0LBNz3PIVO/+Zx9PibFo55aQj1e0cCyav30tbcF0DktRl+q5veFPA0UjhpXF5ikK0in
X4njkuh2xvuQxw375Rt44ib59NjlkVSbDzj1W3Y5hczXYjk81KErJZ08cQ/niZX6cCajaPS4eMfv
I0UUlC0ECxfzq14WxZZ81gfsfWwhaarMuSRA8Kh5eqIy//i0vfGrRSHj+cTYjMWmWPQPM3iH5APq
fJpmN2qLE6R5Zj7krS+cMkxnqMJwJzwb1qbSfuq6AeahtmVddBk66u+UyMG7MHRsowMIAu6Eg8FF
hcQsvkGGFcg1UpwMVmVG9o9djyI/LdipVdmTC0T4Q+fFN/AFXcCxeCVIQPh4BRBz3q647GaIdRCw
yu2FCOyk87U/PcP/8J4CVz//ck9l5GGgSfMv9GZMgDg8Nk6krB7oAkaidqFU4VH+LGll0+Zbo0lX
2n22nD2u0Y/4CkNd5I+Wi4h2fdXNyjQjmLo4XAd+ebnXDB2fP6RPNc5eO+nbmcLwuVKdzmUeptUx
dl15HB7nyKl7+rw7SuAjU9TNOgssSjhvcxibfR1ws5/s+kS7WJyKUMrHgpnfN9pWomE9sU7VGlg/
3zmwLkVPoy+aPnH7q7olw57X2nLy+6pMKtEbg+v/KHW3/0z6SQviyGOmtefsaBImKZSd+jlefkhx
Zu1ZJrdOyV4XM8E3REfpacmELP2IKK5F5C+aEhjGIr19BzGqTmR1D57Tpk4wnlRTkGdnGQwqKO+G
fUHzkAQOQe+0yIv5TBxADvPM70DgvwQkLYlB+hTdJ7YT4shJOk2DQdvqQMzQ6XQfkaN/w8qTQDm3
YXGgRmpiKPCgm+vExRjsmCJL3zIkTft88UGwRJjNI9TJn4j53KXaw+Hp77cfBllGqzJEP6sVK3jw
LmN+GtxeIyLdO7sogDk9c3faAMcX4S0BMy8AMpkHe6l5BgKCv+u00vGxVGxxrpwjErp0I+fZbMPP
jWxfl3ayfoqUwPFeMaeCcQL76SV2zrFn2lfQAFfm9N2kR1cEWeMpHdWMl2yI1MgRqAnTI1CNcOFV
rVZsEYJJl9IN7yobasqIqklQyhoePpDKVqacirgybulUQqZ2VZ9C9YMvtb5zK9hpXmIrb3Ti2qC0
CPk0Dxl7ek/h/VoPvQlS+7iYOcN6e6LdSqjOBry14bdFockBW2UogylwbBiSGm/oKS4bN8vL3jp9
anvKQCvHhaKC4rASRuJn/xEDe10seB62XxvEVwnWLKf/Vny08LNM8LBmeeLkzcWvIp6eS2VnfNhT
PLoNAOSUxYK+3AqAIVk2ZD+YkWbD58tHRLuMWW+6h4XrYf5PrHUwwqWEVrnHwxpui/TeyqX4onm2
inJHEiI7M7vIB6Kjw+lUJSci4PcLYwtnfLsCgAMUwASiqiJseRgHD618h0hj4rJJ1MD1CfPvk2vt
9Vl0K4gZ+HJubCnbkdqPH+PnpwPnPp3wqBKj96IawPjbLsVcJGoLftX9OL4ZakrQZjj9sd4Er/j4
jS+XwhVm0VIulK2gDQY/fk7aQab8D8uFLEJ5Y1Ti6PKQVkcTccqUwgHp20tkXacyMzi4uvuRalr/
4uR/IBaugzDUMGpmBqubGqoO/cA8ERwZRv4ZmarYSYLLFE1hjquGteAfaRCHTE2c9HA1HI9dHbbF
uVZLcZS6lCbImY9U8B3D+X+aiIgG9Wbo4F/bLqDQPRK3BmgUYhFH5fu+Q6x+EMGkm2KnqRF6roD5
jhfF8b7gKR5ZZBVcw809dhX/iOU/AxYx1yAzZO2a6XUiUdzY4cWoIJMENxiiwlHswdY73AGs6HnI
KLH2OO4p2x0TNT3bwu4E/yiMGWb+SZr2TW4CVhfCZq7hU04SZQMNpmN24hRfDL7HSrvzrrDvbUAe
t5o5fDkWlVgm9x9I1NnRC53ve6U2HjNNCx11LKvyWoLwwh2MksQmLOSJIUTn9/88CarQLbRYoTYI
NQlKUkgGkGpq9wUSgo66o7gz+dQfr8JVu6NfHwGuBiUfsi1qUYXlNpT3nLMVEKNqaKJR/OgtEIDp
R7JERzcO5ulfliZNPtb19ctftvn58CgShQfu98bmOaS71wh8uQjeXh9J5QyN747ANemjp5YkeI4T
o6gkCbsx37Dwpnpjlqm2RfI2f7RXMZZuhrsqgO3yHvO+yJtqjMpYGXV9Zo6zym+axFUCyoxI61Uh
8mEDaLWHikHRrwMIVMAc92kqbkUdxZOR2k8NpCT8S9KbPovO6hq7XTy8Ms53OXkCGXnm1PbPjNCl
LWhqAamPtsLYDvS+pCe9LCgPbJguSu+9hf0UgYRHpk7S2vd/V345SQ0Ak3do60i1l6wEFVWjpVFn
UFqJVzK3XL2GLrbwLkZQHRGNMgM9U+Vccjui/+4gbbnm0619Tazl3TGFNMIX3nxuSTYQ/3hUd0/U
EEZB4dD9mo6IsXIJxrUtQwz7gQdj3/q498w7ykA9x4nmLyqWJS0UMmyehkRfuwIWSrEgijeiQcJU
yy+wgWoBCTM8VpxvTcmryl0qYSobqDhy5yo9NriW8jbHD5fKX41Ck+vWGov6f6wAcaIpAWmxAUkW
uNxcXKTT5pWJzV/thVBgNtylLHNBFZrOr0kciCBZeZ0dPM7u3NB9IzT6t3bmg9aV4WtpYgb7hwHP
xnn/XOReX2pWyyXF9qPNhpRTPZTjB5J7iN5c04u5lraUdh5/a/HnoQxg6a0z5LVsF0DLIvI9aqwZ
vmXVQjE0WOOoG+aghI9sIb5NjUDsOJaokrJkxh2y9YAEYHdDe+zwO4Ns66FJt6YfMUpLWtFC4BDQ
LwAj/czCFqoriYG+0O9F2x5oLUwMTe5rNmPfJS3bMZEVI4kOPCwGou0qvtYcseuC3lEvxCTYWJXn
wWNEpcWXewgix1c7MGSEKCOlYlEaFgPdIY1J+/1mYuWvEL75QksJrBWyT0ecCQaVPFLl48oP9h0d
Y5APWbILFPrR2qfEKoUuDDOThniAFWYDK7jLw1I1KadPRcjgdiqGoaMKZaxcXLEZb0CoEy50ESsC
izEF5Zu3prltnKz5qhMkHaELzLSkXofLw1nxXMAS0ADSHXEVYDI0YujyLwG6kJVFBSH2wVz9meoE
L5L/4YFw6JvEt4FSmvJ3raBxwH8Y4bA8/uf5HbIjRYVT8pBKJQO7/hyadR2A+mbNk6OMzMe059cc
ax8QYOU+0oUgSQGQ1qNdV53XpydZZ2XsGIroEdB8vezTHiaI8fO8+UskT1e464dKOsjY/XY6zk5I
//XT7AqYnkTAWy+buDtSv1aJI6Kiusrn1YEp/oH96cOo3mThqmh72/qof+cbD1tn2RRn0MbCcmo2
02zLmQlWaoAn2x/cdYtfimFV55wZC0lXzLxcrSe+h3f6zJiGEXJlD3IKtWvKkqK3RXtU4ATAsaMF
aSBKbmloDONJD7S53KXcreEe7XGjb+irQIag8HL0MhEKOPkGZ3ufzfc32WZza0I9njzU0wkttXzS
Xlwtp4Oqpg9a+lOiuQSmazc4IA0lwBVRPopBbVgan4WRdyk9Fm7RUpc5PxDZ6xB825LX1W8WPk6F
BGeprRwDrj/u/+YBoFIhTaXW5/Xgx/IwTr7VQbvoojUK1gc+wOquEgs8NxoT4AA2k1TiUALGo260
SlQ6CT2YWxwn6z7pXn99FP0qD4GruwoILZZL28Y/Nop5TcQeaFbvxL2zJ1UJJ3hpzN1Wy/D3ih7g
YVspEkjk+g0CFgOPHv+UPmnznhR7MBpCK0Axj9BIEopCjs9UKG0Ztxhsn56jtwOkcHm0Ku48Pa48
X4NQS/WQ6I3aokeQBXRzFdz0INTkt6RvlcjdZ91xALv3WZSp18GhYnneFKk8+CRiF1Q9GIH9DpYr
05+RwJZLvPwsvipyImXICJkoWxDGfmo/J3YHx0GVdtPx4Wj9dIFC9DAwFl3nZLkrb8mYGLJZcTeT
pKrtWLr9hcCv7kU/PTkYydnpjaLSxWdU0t+wfmsEJZ6Qell7j7OYuu+hXZjRFMFxmi4vXPmqAfcY
h93ysOUzNwy+n9lvTB4hR6Ibc6RuY/dah2HjPTYvkkxjrGr+JzmkIuoevijPUbn65j4vnuzAuX2l
si8g3zEicFExKZw69ffXyTPoD5/w4Sj/VwBYu5ee0t/8Yc4GDjjB/SYFex3SX+SyUoa3lL2D9uHC
imFm8jwBHtg8DhGqKlUs/jTXx2nJ3QbVDzZlWXa54neIB/aLoB1Jqja1yUHFamfdG2ooSizB5llE
WlOmlC53WkN+guNcjut2n+p2Fn8IfJyfam5C+5MdzCyUTmOKDfE7v3hUmNLyxoXbxSUfpsmsD1wD
Sln4M0UsOfWDxfQ6KqCPekhOXPgabOwMg2FeHkJuyUEYWHZWiQkldqWHvzGRjC+7fufzKS0Yg3x4
lxhIysMBpjLut0e/2wO+16fjGXOnPiQVtYzxDep6gFX3zbLnB22h9FrIo/8HzZ07gTkpCBAMcdoU
7OnqqLQzuP3vBFyR5YlgWfMQeO0oRHgu/NzMRJAGgyza6Mgf5xUKkBzUPE6gKdMFvZ7Y+75aBRl8
0pp96b99x2VnlpQ8VlAClVj3uAOG+Q197URsUKGoYRumcnKJOD5n0gRiCI/qKxugaeU1k66zj+p+
BsE//RWtOv294YV9UY+MrWipXu/KEzmmo1n397bYkpbmPymlkRCiH3Hpsa9ABWi3dhiv1lCOQFdt
hpjl7KrGNZonUSi50ba/pMu+5di+Q73E/u/xdpeO5tbMtGWwwjVRixAb+G/JLBvqgmgPSDdQ5z0w
skWRxvaAPXtvqyZegMVoF24cTXilU4xub34mNuVSu4QJ8skUBBvlBdtfVv7LbcwqA3w/B0iUUPH/
oMJp1kDKJXnEtf3cFkOZJlUny7/VTX9HixrYkUNwYeO0BWN4LFCOQqYSQpDzfitHACAcN85Qcrz9
F0P691P1/iGMcDTIF3j5gwo2RZVVVJv1AMnltrhV5+snUhaDMa6EpOkZQMryJdQb4PeuBb+hW3PG
WXCl7Ymzysd8cg6wgmbuPMikIqxWoXGGBFUceHJVMtRTRR/D/4gsVnxwhkeCSBkmgIT/pNqhUxVA
j/+ry9fFhrolXapkjN0o/jKplDzwUmnvIoTcrR+IgNEMsyKkPZru/dRejvwIT1WBE1B8l7ww2YxH
V4lk7BEA+b9Hz2g2v/FhsQsrvVwso7ClHFKDmrNrg8MMXY3myJ1b00xqBNTlT/xNUEREt3du1d0/
nkx4dgU3tC5Sp735/7gq3SQQcRXAYGMwKf5u9cgLajRat38nP0MXOvbt5BLuqQwX59CPnbjqsOEh
6NW1KbAQmmvDkslgjguMR0xMvI5Nl380+iNigE21+a7H6B8OKlyY1DMI32BWLaq1zaXdrGn8TEWF
z2BFIb5DOT398qBTfghSgTVEIjDphQqrt7ymuX/d4Z5bnik3wPQKeyjLkgp3J2L2QzMmv7KIOg8J
/NpEhWVMsvHs/mILd643P8/hDq4RCZ4REizrh4Rzuua5gAEokjbHSwCHoyjuSP+FPNalsCNYJnKk
02pdfOSoh+4kQ9cVBgeNTw7n1YnxXuwzeUlrvpw/H5Evn4IHU6PbUy7E0MkEDdxr4do/OehcuKxR
imWnS/f5Cr3zDq98v5gwU5mDQ8ucjtKbBXXEh4Ic3OI/G0aSCwVbDhBrbXyw/ebb43pZZCNemPM5
2fux99z4+JaKsbdcwHpRWDdpLoTyKp0BFiyE3J8mqmts1gJU2lGYu5QRvIAp/zJ58wNudRQfVAt1
EQQIY2YZm/o+C0tvKviDuyk4pVgdQdYb9lszmmSNFAYINvnQj66uWSkCL80AVUM8ktdPUJfl+L7o
faAEvCmgwFT+NWb+A1ln+HBk7zLcsORLgl8mFHdtKGUC/4qG1K58jqh7572rVqcJ1LwZCbjLUX1f
6PlI40fSHRGo+w2viDcEltRc67LBiDvVeeEUXXHdg3WTvr4BQTHBndF+eAgqAlpKIBtxZO+lbDZG
dn505UYKJFQamwzT/6eDmTuPpqrfioN9FU9C8m48j4d1YU1T/1VCbg/qED4mCr7dxSAasNWpuBqX
F12ieTlaDZgoIwjFd6NSmyGsFg8XAQIddyfCyLHDRvsiulBEImWtpLGVSeEALS2kv5xPWLH+go5W
Y7kVDGqp+ngDc5WVhMIJA6yiufwT4WFfomC6vWjeXCt7tp97NNPf10Qc3ZD9PQs9sU7FgYGFbWND
NtDmbgiTUOQsSL8Wr5fp2qnRDvpYuG0GfZd1zMf4+21ve/2kNVnpoOFUnQ8+wKLh0WuVDSni7H2D
/dSNcDsNG7qvU0h+b8WhReZg+nJLFTyClaq1w8z0Vvvai+/7fkp9i11HwBx8NPTbqiGEdye3koYH
uuc//sPlGkOdJ3mtLqYazt768kfxlGZqsCyVB+cn2+fksr6Zbu3J5vK36800UOfrBB5VhWmiGu8F
QP68dFTqSq6lRj8z7tGMtoEGV2onMjM54fXInxCH7v0aAR5itvoWJyAfAjtNpEQL5e21/TQHXhn6
vEF9owUam8zYbRCJdVLBaKZJHoXdXUXg9+kf5TWP4J36Os9da0ObVnWjyysQvCf94XH/lUkQS5js
pUMra4VhMfC6+/PqriRd9zOcSn711EBt1iWw5FVEw3beG1p+RA63UpCvCwAWfYKnjdXb6aH1Ogd0
HJgBme3jGPcuNvEccH+9vbc5iQvBzgX+bydZc3Hf9GOsGwxLItCv1HB6fO3OjeQNzl64JKarmuPg
MAjm+H9lZq2T6uBWf70Ab//TIOGpodksdQgfVgcul5gY2hNxPP2r9EeFMm2PalqesP4rt8T7NXA0
5bzzJOam686+wFhmZIS5qjo/+xcqoidwRr7L/d/6Xt1MX+yldKsS+CbwhE06IVtkNV+/7RgUomIB
ByPX4jMPSD69T14oHrnMAgICuwwoEsh5q3Bq4NgdZkOrVAs9/Z+AO+F/NjARRN7ZpiUwyLwoshiM
tgvbwbXQ4aNeXe4d+FTrrOP4WTk5ygjLOiUr22zCbNqe353Qv77laRJsgfIFfWfI+dyAQwjbEkBn
ZzqXfnoL60f+S5BlavHeTPixILpWajcdbN9Kn2f7PbDom6eJQQT+uqHtl6CPd7X4BK9x03X0cGqE
qEswcCCCWIQeHVo4UhBnO8rQtT+o79NPvgIEw9B2FqT2aTpDTfCJicmEqrzNczH9gU2RDfcT4Sww
AGdM4NZ5TFGEJg0SPa3V6NGP42SBdOZZgESoAoWFprZKH8NTBeMWA2mWjziw1vWpX9vjG0wyRJxC
UPDYI7ggFEvXpJr5Hi9y6+h4i57e/glB5P4SSXPBpNuAgJFBFcyIfHK0jLY0Feqj7rHRpd5303j0
FRCs4tvDV492OPC0o1Q0uPKpNUx5S95KB7BO0sMmb57zjXie/SwNOe77x3AHq3VOacymj0G+VJkN
kmDRSgQhXUFEJeTYn2wo33wfR5NZ8ap8+XkIA/1OYNovwkc3cJE5Jg27AT5hAcNNOxiQt2es3qYI
bJZnbGAbk7OQ3rAwcJXuPyuxXCeIgIB45Tgu7p1bI0kGPoPHRlh8npj75aImGcfgfsg8H5MD9MEy
p61FZnSp3WCh/lMaYtEONZ2AQeg3HDR6dmOJSXb0rWQ8m7++OGR9qTurZqs3q0hRJhHMNG4l2pF3
at3rGoJKkKg0MgHDSOmbTfhkbuaL7AQ+wI91nz0H+/r/QrRPRBJFbDKOyPRmz1M4xsnjL+NCQ6ml
bIOVnZNYpyKkZEgBaasy0KFBmcOc1ZZcj9HykU/HwVBs1sfe0KkjzdKeFjiizTR4MurPa6Flvky2
6XJQp/zrRwCmiDsxiPdSjVvGtH/owJ9XFMhE5Gm2NL/U/sgUw0/fOX84ElxwhjZFQ9Ad75qI+M1w
akFVUrCiO/+NG6PqeH31o59J+v+N5toHcjXRHBEVQ8F5IaBOw4SrDR5lqKhRG657zXEgHsor9LU2
L4yeTXfdOsqa/FZiu1sYUKaR8Xej90Ticu0z5Y+MhsU2zpTOAVlm+P6duFS6rgCubQcrjM65nFVM
yyCrDmLz4SwmRnBa+NbLSvRKqnVHQmlBX+evrk7FjiU+aQ/uOHFjsq9sblJtlkCae8m+vvOzt+zB
jYjOV8WNeYwc1h5tADQXTg32IgcafOxcVYCicO93H4/IDKlNvhVgiMabjrJoRHDAWBQdrnqF5B7I
Lv68ds6RIkCTYzQ5K0SdYNE/EBpd2r16//i2wiE+FhgzSzS774xHUjyRjqzuAn06ta+yVOg0L5ba
kH4D3rAR4ugCc3+xPCPLmktxGKeoKjxGWZvrdnpnkA4wDTs28g2KmRdn0ZH3IxtUjR1W6W6d82Li
SUz/60+A/pxulovaGi6KemZtgAGqoOBbko0YlEOI5JVoOdNx+XkikKd/fldtPqw2M9VIz6Y2yXqj
7ptTq8u4d+w/GTL2EWpFB2d5UCUxhMZ634qH/0FZeYPMMVQAz//pT2tQuEnblqMxnz3KNYeTqQ/z
ZyWpamofhCRMhxSKCUHsHHtANQPNHjyPWIKVb8y1t8bpKEVwifPYb/yCbiQ3OA64rF5Axjm3Wh6m
T7CURdRk4o1bDTo+b2kqEzrLJncw6gHVaOls+rEZ776iZOouNWU7+TSeZwJu2rH+LaJkq3f7eF4i
SDZtWMYfQ1AAplkHs8EjXBWHCd/Vu3n+8YGo543vzic5W3muy13eMnNBUH/l7CiiXSpwJcFo/TRv
5neL6zJePuCRPMN7g/g8QA+s8zU3weS5ePkMoDpMc5hRA2N77v2uV3EJpnvH8i2ExaLZgb5Lme9J
Ru3u2jlDMR6SavqBDduSGZZ2cMKjWTR0f/cNpeBu84tgjPkYnqTJdOSa84BtUNkGgz68txbbad1i
xVwYWD+3oqQ7FyQx0veEQSOVkE68cRxAYyI7viWZteBxIdsiRFmlltUaloNGbFzdJQuhHqlsB7l0
45fdjAin3gLfy4knxXYc75T7lKDre2bls8yxskqNm4UzPYLrQ8E9ux87ug6CTgiTy1e3KqIZW//d
aW+fmX33ixcgsMrR+aaS8UsKyq0aQYS/FeIb5uPJdtxbw7f3Y43Sc2CUGGUTO4HJ4AZ6U5CbWI4g
N/F/DlQKwB5lvc1RaFAPYjhiI1CAKMkAptF7+uU6Rs8zyn/F/s/3smB6UUVbmK+2aZQ83GR9Azou
EW2rInk7quMtNhbYJ7M+6GEP80R8bMgEAFT7mdpN6fKuUY3SfJzCvClOPqpBk0/DqdsNiTIpC0MG
oi8KiJgOZwAi5bruEfF4ofHkiAnwGyn/ejYvr5HPcI5xOzXH1HvfTgXpv9p8y0jqQZA+31mR7Fd9
J8BgRvCrWxim3lRbOkV0Z+HEfpkHv9XJMNQIwOL6SexYjVAunuB7r9npEvrCFOMRNq/aR5V4RCnB
S+BxaLBEkCbqiXpseATatB7jK2/whmsIYe0tkKoHeIz1GnRQ/W7Ipj+4iIcitEcecQtrzUdApbQN
sBqjrxMzqiKka7CnYNyn6k349SOUjx8XX40652ArTJTXdNmI1O1SYAoGxz1qGanFvW+BrzrNj2dw
fnlebDcx5bVyXCBygPDqgvtm3Fn4uwZp1Xgm1pekmq0IUCqAiplDdxSAMYvf9VzwqRnhGamQlqaK
G5PZmycdxNrMdulmzv67gC9rWSffJh0iiDB2SwdsOEZTQfM//+/foEYVoZPf+H5jJWNtNU3p2lgM
xoCXfHMWeIQBWlJa+9v3bS63XRWMt9vfqIH7AjCIYAeF9UNLOnJ9wdQOMkGqrV31rqwZo4R4EMTL
On1VMLK0A6GZpINf+fngGvuY8IWTIl7o9MgFfBb3DiTL4sOSI4NeoDMsE7IpNph04aiouLLcHUjZ
R/7Sqbcudci4fCjjXkRj16VGVNFinco6n1tSZLCtsZdgbOivqQcIc/9rCMAkJs4IeVHpvPg0tI9O
JB+IuwBawzGyUhc1/H6ik8dB+AmwxU6kWjmsQwPPdKhjJdincTL8Wie8mpa1ufVgNxCJm+eCJMsK
22URJUlAb1ijbpnM/1PU6OQ0Z7qBeaqnk15d0BHkIbMYO0FpwdWGY9zx4lopvNE3JMazRvNtoPBt
zjii1WhUFIFsjaX3CqNUTWX3K1eAC309PliAo6BDhQPrcJ/0d2VffBiE0SaeCJPyOoKNd84BWA13
S07LfYclMMAuvTHZ8oQM+gpI4GJ9/x1afSZTZWFyhOKTOg2xdpbbdfLEUj77MTJJTDDzUs3/ne/H
eve7XHUKmjv2s7895JTsNX3DLiQpAYjdeNejJOpObNJDpU46yCMc0MH1aQLpaKmRAB4IHymvAxQ/
+bx7vnEWgb8Y9AutP4nCmIPoR3KCX4FOzZBpmgPn6xssBa3UjrfCQ5O9PMbIz0LexhHHOJg+3bQx
szLezZM1Mw+A8eSQWXVn/cyeyvIHHFqLd6/FVqdKuTyeYYEHqk6CUq/DA8LLGJaVcbZqP1waPFzl
ewwcaGigM2V4NFuhgDmi5PO1s5vqWnHczpkyxfJMbZh0rfBUbsBoY5PB7852xO1MrEWipz53X/om
/58RYcK0MDLI2Ba8Iy/0EOooMs+8v38oKQEx0/GqAYG+PAhmwMwCmO7pNt4szdOym+yLqaX5FTN1
Scyx5K/QaEw9L1J/f2rDr3jUo47CmdLJ1rryiSmPjHUcQc19K5nrFVD8KjHywYGV2hDxxvgEFBz6
rGk7vSx37vbHkoIAs9IGgyPzWcX6dynWEufvrww4Uf5NkzUSS/0fah9kSXxa8dp/YgY7ChQPpRjV
SFoSjtKMMOZGfJ8Qt3fqP8r/c8/HJRDgPLXpbk7AewWg6frEgNpDEPiEQpGgblbsqTsTM9ZNpi2H
xf80V3SXpMNzK2D+AQ9Hv90gjx2Cq+0HmLAMiTddKaZuR/nYQCcP6dXUxNrRCeurr/wccVSyg8Gs
03/9fED4RmxVnyEk+ii22gTIsuy0onaL5jAxILO8h6gZahKJsv64I0gcguQfZGcz/TJj8Z0JgMu7
vvywk4gdFLFOpCsoQgngV85VPjop9RVwiWchRqz0/7fDex29lyUq5z7UoVV3FCnAHJ2g+IXPmDv+
pjuf9PQkDhHzMc0oxXuDxyEG4P2EwAG0zVCfbPPCzYK3RZl1a9rxiYmzk3r6TxIqDUCF4XVeoWc8
bi76zooYad4OjSx7j00SzPRjHQjTqzV91yynjharjrMHZj5dErWDyo/K/YMKTd4i9JG1UK+wORx3
aLPGYoXTxjele9io+ZHZb7OEiFgBeBSZTXdWVFm5VXsLo+7vvBLclnNqxEHjx3iZ9Uw8hDLKftJK
4aCvDOMcStC/4iRn7aMS67iCq+a9wMySB1/7mpxxp6/R4zeXLb4y4DBOk2yJuRQVntZot+3JS2iq
zUZn+J9t3s5FCIwrIoik3rzfoXzZknmXvRXNpnhHuylCf4PE7dFG3iR72wP4rhHon1n0f8vfSxqz
SWsJKaRTozJZZMQCDDJiHrBM2ekEx4EiTocExU1QfsL/4DOnoKRi9pcR2Hx9G4j4GDg9qZ23d8Kh
OZEPEe7dz6/Eqzpav2cZc/8shPIZmXvamtwxnzyTI1t0LiRqWQo37TZcvbnaUkrgkdvbrHAh/PI/
WMBVQ/dynP71cIVewJxXzi4NezLO4tvbqiidJvWknbl9HjFEdu8PrFgfYgwDyWfA7bJG1ACQ6MV4
uy0/wOozSdFwfC0zThqxlhEzKCIYFufdLI+UCoJ2tRuDUByfM1Addrw5DWsgKCcJhANP2bRC1J8g
S9wwMxYJ/kx1/9Unyvtz+HUvXWKJ47IttvkXuKmE7NqNi+ZavNlQpnyyRDqy3rWSo9QjcespyL8D
1ly3o1dP7yG07iPhrwELq2CPqqf6DrHIml3/9FnzfzqLgGRqBVksQZoghUl+pzEZt7SVINjRHp2F
wHUfWhY0p9CBOSdDnwDIG7HfUfx8LpWipZRZYPUhNQ3YHDCsQ+rRgLHQZ//ApbLW09/WIDghNt/Z
d1Aq+UOZ0V0cyiv8gYMgRCvidBBTvgUKOSoktpc61V9W5AILpLN4L8GuixZ3kx+c5Xh3ThaEv8NH
jkyihIsqQfEy03k+AQIVyepWLOWC28xrDUFNFzdCLh5cqDqbm+EBC+wU/ZWusiLEy/fM3IhlO/0b
wmgzFuTWjIZAixgQ/THlmAEcpSnbHtc/txRwTi2mRgTY8mJ6uuY76yJVp5o1a4LL6iCkatOGUhCh
wlzpai75oF8aWbvcV8tK2YZeOr8261MX6S+QIjHd7U9SwyyL0Y9IUcfod/ttB2ruBSV5R1RKkjyX
3hnsHtcqH5mdr1tF6PmlogjiKnzUTW95pFFFUw8WS8rZtJZkfdsmzGVny/ghwMHP9LHs36+qOWUX
TLLI3gfTOJzIyc6FO88Qa4on8UKeWxBEyIZsPDZcHmVsITno/BDnCoflQzwUohfsRJxovCtui8yP
aPuHtaAp4kkaHfkZ87jP40R4nK+oNPqxAabgicV9xxkNrpolKq889Cq8Sy9AVJyu7zbCGIDsUEn/
hOFweB5u8NJnejb87oagdrJyjRHSrI2q8iR1FmtxaShsVs5hL41YVEwhCANsSZeHMtrk+5bHQ1zr
rJUZiUCryega14A97JrlEMU9dNsNTL1pbdJoRh+clWjtj33m/if7x9NKQ6xei5uE3OYAIa+WCkab
lFdVK96ETMygZ7QPHt/6KA5MXHlZ6DwdWVxesffoSN7Gt2Jpte4DyBlH+jnKMMSKSGSwSbPgSlS0
GYDABHw9I9H6AyCNhU0HNfseBa40Pnv4rV71OMwXfLjtKFQQiGFxi6g3uyRqlf+4nVN0d9EEafoY
7VS7hhvJ/2Eq8FIDI4Mr1osgyWMHHmobuRq92DW/CIkbDE+kYMdfcDZdw0w7refytRZLqZxTPLS9
KvBZNP821w8ymmPfhz4jCnOXjaYY5Gnu7P11T2Xd4j1seEhxrD/f89da1gpQIGgamn1RsuOIPMdU
L+QBRsyHzaSR5Obe4Zw/aMy40DxZXYOA6DtbirI1lgA4UsYRecHBEMjzf3hTzAMUb3+sJMcMtc6o
ny5YV4w+G/eL49uh9D9NhUD5VXvL7VlhHXcWhh5/o5BjRmWd14/HC/fRlg98jCREUkKHuEAtIZPz
npb+rxa2YjYS8qErVaOUfi8pE20OcV2XhA5iP2M49pyeYtN200izUfecHuwh293oAdvhmRIuUPtv
LYSY80rlCBqt0+isG7iBTHgr7r3iZ8UOPfFfz8AT24KLrOw2pNLux0DcS9+sGhKNHwvhQTWtWBdd
ZknCRhkfpMvLR3jOnvSK+JmZAW6xuxgqrIffP/EqWJ2pypg5cP6ietFAmPY44gBvu4slrf/VhqsL
LbXcyfX7hmpkV0F0tP+YRbgrJO+MhY3F6uWYohsvsAkRbgYej+r/YoAPKLGXKE/70LeZLICX9SFC
tdvQSUg4ePdJEvDxkp5hw2s2XjdTRqbqU0Ot1R5ku1IjxDWG32lxsFYsIMheNqw87L6jV/MG3uc7
4VZhUdS3AdpxcN10/+xik9Balb9ZSYICt/pBoJQiYG3iMSK7GbGNdChDzNiXaKBx3SS4w7gBWM7O
no6pB6AJjA3ICBPlaGxRWaE593FnYLsrrvDsPYdL8VfXfvkMZXaGpGBg6UcVR+NCG+5FeNJnGCEP
CLyJ2KbW7vB1UXLMfUDv43DkqKGGrp4/bXj+EakWmRoUytFCsGiXhsbiO4EKBbBTlIAzGxEDPFa5
Z8YQMDprdTFOuWnyVoxXH6TpWRLUNzRGU0SNgd7gI6RSvXd02oeRMIPNv8IOEWCRRPJmOhIV+f3/
esJJ26w1UU3EIQN5Amz0UoLS8kFrMdy0s/72L5m4ut7gSpj1Mw2t4LwD3O1OXdhLmLljVemjYzRP
ATgIiCZ0CxqjuK7SVw+GaCNTloIHg2Zjud6KxShXMVJFWC9b44P7Ozd0PMuwjecbFsrLeRgAVCL8
FqsW434hAniEDapVJxdPx2GcB/re/kdrKj6FtxVCSq/E7rXDI+MC6qbyXtB2LahrTXoXXmAQtyF6
MtRapACOcMPPvcpTlX94q3u937hLaXNTbUHFcl8M64gQSqihQ6Mh9m/1oILJyhM3Pf6Q6fQ+qK97
eMpKraF7YnxHcrqSAvN8LvccsglEzMr+GlBlTD5c1TiuYvfhc237+Adbj7PXS5J7Qlo/Yltwqgp+
VlGWNWhCnXfD4NxLqjkxWha+sAE88Bt1A3P4J43n0IyQSNMb0vORtlX+9b7+Tq/R/6NyiVWSujVh
2zxCa56Ejsh/0D31K4JLP3wBdlfO1nm8bZP5yaZDOn+uhiJzyFZWHlhv+jyWifCIPQ6Qg5r7nZRb
61BsbsItf31gqiVAt9LxHIYlRw6pDNeKT/l6toppQZYHimo5NweKE4DZknk4A0TwsRQWSKe3nJpw
6Qa2prnmSVTnJZxHZpL8fCmFlXuLoS7iaMgWoNnvYodJiZMJpAa9HFZ9tVTCiUV0sLJtC0yiXv/j
YSkiolDN0Q/6mQ6l3s0iKxJmn8eYVh0ehxGdym53BC3F5hfAMyBHI7cNrh115bedJMWv+/4kShbO
T1M/0nzrDl1BRfibyForWIRr4ceJHWLv0o5wQbY0BXjKdIlxmz/MOh6lAP2iW572oVhH3LixCveB
ZQX//zJEgY02DVEqr3AFu1cAEvGQmrgaSkq0MrdNAAB8GdNSpY6p8BsFcpannPgV2vp8DoC3GC8A
5FvUxamIzkR7qx1JzjAXprLlTEF/wl42pc7lThyGDYxL1lNmzqxK7+KSpVPG4sRs7LHuS1ladPaa
4fIseVFjHLbL5xPVp2yOew3WEYmNsHs0UFfwzvcWM8jXKHgEpSI/3qNnr8KMPItBnepDADbfEc6c
CFcOi8AuWl5ZSCE7IUZzDrL5fNdHcfQlKq69BIivn2d+puk1N0w51oiKPteFLOn5S85P9nK7KFnp
gCvlgKgFBci4IuguwVR7eyikiWvYBMMzX8feU4tlf4GHDYc5k28n0CrpifFmcRGtm5Ss+k9vN61z
RHId3O8fYIcuqZtX/rYW/zVpW0uN0MvsTWYT89E90o8S78WTLhKI+O4zEG70Kl9GDZ7FJbRD/YEu
ZfmhijNaMuXX2N9rkR2bHHh/I2IY1+zJcnAUdyCXwGNoRiPYdtD8it8n1Tn1K+ivof2SKZekGiZD
CShiCQgnLw92xsPmn5cfPwk/uYMxYpyj2AmKm5wPRtPimGivWJr5HFH3LEyvnhJFECOSc7quuqFw
H089yCptgvvx7DczJdNrCfFoFdPIT9HfjsQlVQUlN3ux5PQ5+iS3TMsAZLP7ZTNT+AH/jMFr9waL
uZUvMTSZlMWYTktbR20zuRedhQsV5Bn0biqB4vLZr5zepAz7eo00iA375/WcG/H+8PvR0B9HkjGq
frTNIuScWH5hq1TrdVcYmHgWktdPi03Tk6xPUjYCRPdnKIGLJeQp9Jd/hpbRl1qqA3BXgwImDGUQ
kyWABN0PUtzVZtCAq59FzUCz0Jeia9WznNbKK9LABENCxPmYX6EsuykPyORRKC6NlmrGmytHCIy+
4gFJDeiwoOwioQ67HlhX179Gdp1WweRM5ggvKJN+WG8OKoJJzIjJkGiUCZJ9poWeLv40xvLET40K
x2+o4bjDCUsq9hy3ATOdHKlANAtvEqdsxRwJ6rIrjzcyb7GNhzEmZOsSrFv/+exDcSmtIBc9HDzT
1K8ac/ipzMy+YKdbQkJ+rc/gd6SG94Y38HVZptMMRD9quhcuilxNbpq6RytEyyjetK3KtQdFXEch
pSuYDPMwE76IceMYwnrEZNrefyDkwCaRvqnZnYUM+J2pD0hFdeBGjRIrXHQQI5hFu8DIrXVySKbB
qLjinzoxScFzgHOMv1g1PRzFwshWGlpj0431ShJY3ocpa2kA9oZe2jNLF6IE0yyhYOtAqlUXoP6s
yUIOTX6BPQ5hWPTyl4xzXXOW9poIXEp3kpm0xCXkzRFRRnP7zNFR/sYXgJDt/GX2YCtOPuvkReTa
9CR36HYn5ALkkKdnRFTfv+tZh9NhEEdpuFnhTM1jixma/w74TJwpujCZk6BOIaCDl8DF8iN+0NGL
TNLwCFiV4V7JJxDqbmHV9+zaZ/grT4NiS2Qu7YwUe3S1/svHr46n732Jyas9pVNiHvBNXEqhaBUa
ljkO4hnvsmCgSZTS1/zWD60v79y24Wt15BwSwdnF9BuEZQZx/kLDadlR1++gtJCxWNetfmBtGKZq
Lr1nmhv9ysEarJ0R+o5eE4evA6F/1JWH28A98tcUzpvVepBBb+rHpuZTPPDc+IC0GAXe0pY9jjX9
Da2ithcZNYO1N5LayHTG+90Fbd/EtPQA7aR0n3zTV+HgoqFqBMqGvoH9z7TXRomgmQfudJduSwba
IOt8GrPzJNkzTHFwizy4UCjw+BCK/S/ZjmeOOOFzSrWGzZwmmNtR4hGBJdJzAExiynfKWXu0ueWJ
gI8w7z/KUEQV1g2fh4x5k4HrW//yngw/BcXHXI6accKszKAJqPyjFX2JfbEXFCidPink3WyMs5nv
nEsyeEIgnfSrRtRIg6GZ+TRlu9R0hRu09XHe8CNtyy2F34/MkV/C+2DsngvbHgE4/ybWrahV+g7V
rzmBrkJvmdfIkidaqWUFxiR1EHfPbuEOtkcb9puV2K0FTcLREyaFmIjolKgQBMGFAO0gffI01fca
gaAKLNVfDRWiHBV9tQJ8VrG86tv5wlXHNrIIVLFgsOjvbpBFs+zvgdRcyQ30LEIYBZ8xeF1MKPx6
/ywjEtdxjK/oNJ9XtuPhFoAMzEPcUqkHxPHiLhsEPZm8g7Bds9YYN5pplxMrw4/6BEQO/7rBKJK9
GR5CHVHWJl22t682JEz3muVy8/PqUf1tVrfdSHWePmlSobTTuWNjPZlZxndiyz+l1xHL3CoBWpfv
jSIgmVp7/DeXHVS29pHNFFywYKTp8wVsSIJRRbtVNKXR5ee3MEODSY90Bcf1PJAeJ5xRkA4oaxx4
7wGZsR0ItkY2MFDbUSyu8OqaA6YMIn2qtLkB2IZkJNvhv1mC2z8ljXxMLBZYPnQNGDTTqqe9wTD1
5CUTCwIzgZsK4k/JKCO9GE4ySLMnHz7cwuW08KGmnReNZvYhHdHgs+RvFGwioi2Vix8PaTMOIQs+
XYWL8DGKwoKKUfLT0fYUy9wEyfiiOPV7dBmL8V3Bk0Xoe3CyH7i73yJ0bsEss05tFUlJ0eiNEK1V
UtfV5Ezlnks3K1B0TYq/dCUxuxMzdgft9bST2OxKe/qOw71bujoQz7HOWZB1YlEWxvMkZMeTFM5x
E60uWDz1ZrqhY4p1iN9WNtUQ0EWmFv0eLde5tzZn5uS6FHuWAItTWPqMlD2CKTgUCwvXWpwXQNzo
TxQICqLjOA1uB5pyzI5+4g2ebe8d9nfdamOMY+dVVll/GpiAoYjhovz7GqQ0fl9FnRE9SJxaNlTP
EPiHa2zpyDj56oR1YLmwjKQaWrQD3c0hzRwFEpHqgAe7kbZEBOxo7aZWBZ419SC19svYbuieQBri
9ccNtvBgyvnIJIFHs6dsdRpEfbgkKY7u07GkeLoQWxzYJ6SCcAie3Hk0yqJzQDLY1nzOmlUvxvS9
lQ3UhGxFm3iqmKEEETlCr1sQjWxktjuI6Ykw9ec0VokYhrpbrp8KbKtYuqUf7aadO5kg4+3DmwPD
vprotKji7wG3MGlJGN0CYTYqv1/UPwxQnxKmd092qYDHkDy07jNzfXwI934nxHn+rVIRJxXmZrUX
L69b75jzVWrjHMaBW+1b/ZGFCpK2D5HHZ6oO0yVCumUOXFw8Dw3HqMNfzbmZkqLVAH0AUOee324I
wqfYMby/Ol9YPMhx4daNnx8jbDQOjwvNviPWA8KbC0nCE9VpuMdslP3Qvb2NMt5UKEpZxAx8Vrr4
aQIQKHMEU39WcX7QtoAkVlCpAZmKtc6hQ+w1OnDZSIhSVrw1Kq4xPHceW3yyhdy6tTQRr+Hx9Ht5
PRdIfURp5qY4n+WEs/SnOsktjkon2w7wfgWhIcIA2T/JHfh6DPmzJyw5HU5li4+261s8jNpV6+fO
IxFtRNMdgYQ+DC8PbsQW788t6ZP1CCPNpveVqoypdCplA0NRjNxOay2r6UQlBS0Fp5Vfdj+4E7el
UdJbJRGWIc9xybGKIISrRieOuve60V3e+ZypKg4Bu2L+1u7gMIWIvkB5rsBl45V1wUCqaTCP7UUf
OuNAYl4+8qS14vjMckA494szAVq7VbKo6/zKMAf5k8sujnEbDaB8AHqo2lmY0kj6SuirpgY9cp1C
xhJQEbRkKngllaWosOLGuXtjmU8KBxDRX8Rf/cx6ezLB5j6AwkhnODgac19uZs1cD2UcBUeyeW+z
oUv5izH+tZfbC0ClWr2+6GtddP9eB1R6/OMCPHqMsx6Rv+RHomOgnmyDRH834m1zcmcxH+F7wnsr
mPUpt0m8L2P6xmfcAKUc1SeKcW8YN18wLUG/Nr/VS9dOIFnZwkKGmjZeWZxlUXk+CmoctemHueyI
WbWqeQRjdntNNSp9N0ItBmB2/8Bf2JfXbOEY1as0WGDgO61OQhXA5gH5rmqHe45rGGl0G1CLj45w
1uPjnRl8uXMIKB3wmrAACnF1X7Tv3+ag/xBfurmukt3K4Id/H52HrtW4X/AgjBwnOjjI/p3/iiXD
mJQKj+kZtC3k9GqC/tk0FaARCJa6cX+kz8Y4DzpIHW7bmfERd64Uq5BnKII/rXYFIXL/b0zlkXWB
KGYnF/h5MQDSocG/S4jwxqnxH18Kpm35xvoPAw8w0pEO+OC/lUbIkgCu3h+NsVrsMjwHv83IpvrL
gQj4BFXqVC0Eeb9aKi+77pvLrONRckhXNKCLYcm3FJwKMZYVBwUrE8L2VNENpoFHF3yGpKLWy65h
pNsO6CLRq3nwmI/hKnsPfRDvoxVS7AOKD22ilemr0KRpQYsoh+miX8iyBOWqFvnV1dSm9a4Fk942
T8puEvzBDx9/ROSDkdCy5qmhRSPkhNWC/afpmK+GZLE1iv8CDjL1I6DdnoKWkD1xJjUxYdKtEQ2n
GXDv5SZBHfI8HqXXGpMlklmuBLf++1WjYNTVYhv9oQWs6sV7q7dMZ6vfUHu6LD2vTHmfSSSbPKUs
U5FKn6Th3oyOjVsw9KyRlI4hlMWmI05TV5+kZByaqcGbNRjgT7GGSq/g1DfwLJmx3rMbBiZA+s72
JZI/i8kTwTrH7PEGDJSWRMCixG/VutwFa2Ye5AqFGCOZ48RCILgiayoOXtw+Bwz5EzfjgUlnBVRh
5xKHZ+aldaiUXo2qE5CSJ/O1zEDJH/VpfsbK69xuPHHtb3J3iLfjQNRU+/YcocFKvzZr52OQwvlj
tQS5Wv5psuoRCaqXGBKBRiYtdA4XAQgxsX5G4Wg+bzxlfrIsTTxlnI+uUhdFZIkkr65v6q0FsFsl
Q4quCIORAn2lPsh9MJdaVkZ5n0gzDk8ooEosVWMxyiqO/6I2rUkh2ZLlGFZL2am0dpkTs6S/ZaXT
r5pUi6RhgYBTFHvQhvgE2gYJbMSmHNARg1ZnXxVZn8VvArZxykgGqKfg4b2fiYoHSVwAlOgFZbUL
IRZYsO/h1zdlMB0YIGdenVLVB4xvORjuWBKVNup1tu+17x+MVFzTPw8oTgPqzb+ZphAAkJggbvs7
WodHK6uZchSjEtWlHypn6S/m+28UyrQgP1bdSVSWIComRI2qRIcdiGDNUaDulyFvCZW/1Dmqpg6A
qnT0Vnx3+3If3iEhAU4LddvyVGZ7xiDahuPZ2fSBmBLb5Hcserwpci3Ktu/jZYj0/iFT7y8u/RNM
EAasBxrdaNsCmFVWS20BVtCiMPsZYy87JQeZAqEVPzKc2eTR3k+3pS06zjAuE89zobc6UNrz7N6e
Vvpr8xlxU2ReHRxVvxFv7vsMX530t2NAiFwLsUloKMLG/JR1jPBxVlC5LuDHhOsyzPr8VP3Cr3Rp
lS4LPv7PQlxjzBW3/3xKGGQ9I8ijBGMT/WM36W7MdLKUc9WK37bnM/APX3+hYr+SgyzARqkChMrh
9Js90zjrNs3h+o9BbQDheLKrjuiocfOPP8wqUCQz5uxcs2umjxN6lo5TkWBgxAqk8+iw5D6SgiW/
xFDrkt4TC7Zh6F6Jwn4X9vj9q4NlTBkUHKkwE7rrDDYrqFGPXJ1we2ODZvihMp1hCeenlGBlaAXx
+vRMHWAsiXhdAk22kGyHJkmk8pYllQIfdSqXBp1Q80eN6avbizeOqTsazn9K5uOdacbHXh3SOY+4
pPR5HO/8gUdUuPl4as9SF1rW67wARgtdGFCiXUE6U90xtNfO5gBPjJTlxDfTaytA1LOk5Z1EgDvR
+aNc1GdY9foQLdmLT4eSsEzRKP2LZdmD8/fuWFaGq3aCc7HeX1hy2nB7aQCmtEOcYw1lgMFkMRJF
HDlWH5TVf5R/n8i4mwqq7i3uiv5oifZMAgdRV70Jx3/8U4rKV5nt1BvcVwLVVjqWAb+N+DjyLfte
qd5tsuuo1yhuXuEPCtnt1OViGZ2Ghqa0wkRHgHo6kzmY1v8lBhIBQTDFetLjliNQQB5UIKhzu0lQ
IuQK4lV2wXINO8YT7ruTyyAX48b4lzkkABHrYaNLNk4MSIttmWShBgyxSBa51oQ74mRjq0JF1QFp
/7pt8JCCnH+BOHSElo8QAG27Cayn5VTBVQEVB6krzDeGu7SJzdxGlOnP49OzuvICI+LyafRjyD6V
EZF0yU+U8Y/pOcWVlPS+CJ0ngg29xTpsUxS0aPr8ZFdxLtDmzMWwgKCDy+thIc8bnLzdWz9EfEQw
Fh7KV+XaSCevpA+qoAdgIG5fKlXmG+u2C3nHtOu/mJIWzMs0HEqDUF/KP9vyn/6kZIsGXGyHRLUu
mP/Ola9bF3X/H/rI3eG6LCpUVY+Dg5/WsvfNrcIcLmlu3zm7trB+MkIzOpblg9XP+ZO/I19Gt/O1
tNttVvWfozd7/ofLzYP6IvESDhvuaLCCaFbmksptu8x6D6ygwbe6xp9B3/R2wcmUeLVWvnfrIMqR
Ht5ropyG85i585/Agt05b/p9LcxD+tstKaxhcot9TG8XiV6D7aJJU+fPkRODG5QP4QoLz5qvbyca
jLn+hQYVIbdnlf+V1JdmQ1dCG2/AAqAfdNTT9FxIq6vsUKw9jb+KDTdpeJjmV1vEFAsgQMi0VffB
8bf23UDmM+YzFKghvz8EjBgY3woTOmGBKcRoapZd2wmMa0mwotLzp/v3Tw8gYEJmIukI5gusPy8d
pXhISXFpHi335kDnk2Sx6hyXWEcSO6Aqd8rGDy18n4aflHstobVD1ICnVbdnbm4dYG1WyaVrV8F0
X9dAgAuCnRpH8K0Xs87ZeJqjOIZPAXVzgcRVxulSQwTvT5IkWpjf99EkO/XdGpkeplruKtIN8KJR
gtUtgZa2Jzp84v78uUXvjtQnaSe5JM/w8MAqp/k0WuFDS+dBEfDL9ZbfAEuq1mKNln41xD7SWClv
sL5lLPlk8CLy7mW4wiaILN57cJgD+kZLSc2KCsEzNdTszgDaip5hx+5I9qFW7L3wk00ytdZbVeww
GbTFr4i08PgPBNc1ktJURRjBisInh7XCh/wwf/KjDEEJZ4UptZXRDpG4WyDSdUWylfp3QpR49nux
cmPNNMyv6iBUJkapsp1sI2EiXkXpaOmkFfeyeeARVeac7srjNJtqCfMeTLm1axMEMo1/iCWl1AeS
yW7SrR+Dq1YI/GSVgeY6VE/M3bnBRH7FiKM08gvRt8TMoD8YsEZMKZ9sVmbjn2Zkev6TnEoRM5eB
gAXK7+R15ksG7fHP2qeizXSCAoeyNXey8oKa1u1K4m1p8Weq850mkTyhp0O+AK+I3ytV3Vh7KrXt
/U+0RD8ag9RbLCQKzUB3etvfDS0Nm4OKm8yjOO+B0q38BRHoYbn1LJrb/ysEGOOKwXAskPnUOqLL
de8kiEx1z/0DX+0834s8C72sD6bhFgPDhNE8CRSCKoQ9SDPD4h6fInEy3Yeki2IsolDxG1LE6neE
T842JSvo+L5dteDIVEOSdhIaT2kBZBlJ+7wpYq5RBkDNDAEgtMfDUp5y2fuqoRSgBuyEwnQct7TP
PkHGbUZAEYzKtKjS2DzYn5hlaIST2c55igQCBO2PEj8FA2wZ3RFosM1iOAVE8U6mRvU9Gc0SkyWK
3ACCsnP0LxduDRPVv7+N04ytM8TQ+Ai9qyejmJmxdjBCpIbQX5638SSDaPUC+YdJdaSy1/cUDq4u
rpGZgmLb0xgkbHKOrzfr4p0T7tr2D7aEml19odttBP8eg6N7Db4IWClFGtRiwyeObetEelv7piqy
ekLe2o0mVvu2QGHSvVJf4z1NiGhf8qUrLFpWsisOm4uGnxeyyXz5t1bL8r4PaZd3vrkiTWP/wxPg
HV3+YwCnHtjy1c/nV30iHnOsBmgkLCbgRQLAz9sty2tHWQFz6cBqzZFX11LEc2pLAyvlDgSkI1f7
rEm0WXQhBcmYzHTUyY7j7HpNAUAwkrULBlL34oc3uhTTdIoTKjYlcTFVt+KuTXXY53HCtex+Yhrq
AwEpaSn6cSGG02uYc1iRu4+fRJKUzEwy0mvmaI0zeO6lkmcE4HRgmA/OOoY8XRdr6pBRO+xwOuUF
caDzeR5RdYjXFYKaYS3N8w1B4eTBohfhHbuMYwdutbdd9j1N+7KMYor3zRps0z1UW19f6fDN3Rnc
MH59VbmGVD4r2EA3bs38o2bjBJf0WC9Glg8WtAGDylLeWbct6AwaAtPMVfyNl8sfqVouxV2OXkQt
I7qRksE4Ol9dPSSLuyDmZ1LNK2eA4efsRLNhDvbV5i2UB5EHJ7MYfGnrqUjB9PrykMTyNSkUy8oj
TbKHJGBGFYZUT0wWAYqzkcqZmYvTjZPmuXUVbK/G7I50Uf4HplXfk3AkzvTJX/iqPP2wi/ZHeUOS
dtOq3nl6kWZD+vr/VNO1jKu00KI3H7/2S82apte4ruAeDSELcirYLtUw278S5HPXXpPLsTJUJPGO
YOPJF1HjN6rExohn9IYtjiUmM37z9yS+I20ieRQ6Aio7kW2eZ4EiqDGMBs5nn6PRKIRwSwaqW0Ri
Te1w3vR8L8U5SJBy5Au2ZgkCQF7ljU/PF10GIoeiqZ/q/A5gttW03wyDDTPMYGB/vGQ1PcpXnYxh
Atdxw3/09NkTuMonr/0csfqh+odGyjbbo95lKs8CM9Z2mRpYvBOHutYRueTXq0ULUREArVBJI5Ho
CGo6eajHcnwUZtGRSG50Vd4MEFIfOsR8dJ0udYP93v/hABrOaAT/YoAMYTbH/2RCR8NY50mMcLAH
iL0qeMn/o/I+S9Z7bW3y1tJP5roki93/3EaeHbhxw5WAm+95DARrWd6//TdVilnxfvEkISvNFv3Z
CPpztjtRHgyqNEklmpWOD6ziX/jxs6M69299DTYFg+1MB1/vUOQrRgmZ9lMnnt7NJL4HNBaiaNqA
5xoHcFRjKNs21Q8UWJZSPzkCT8YU6/u2BH6IGQmhcJ3R6XgmYo6XF8jAzb0y8HRFjt+XmjFnvpq+
FAXiFZBEaUGn4WvHfP8RB+hevbH891N0VQcEoaLNpUbgGaBs8GRZ2NHxIquTRIr41s11SIGiMOaB
/kzNJVuASeb2eazl3/X73Ivu2Denz4VASmSbjVZaKkcn9wdXWZrPhWjehgmMsLiGNXb8OwtaR09W
KR3pYDPcLdvEgypQWSsa2gYxeLfmLUQaOJjGkhAcV4kFNWoTRJDVkpxc6oZE0lq6NyUceaRn6Rse
LdcUHHk8atWhXu9CwOLJzL6068m/UvaUsbg8/J78FlDKHdXhEF4ORqVt5vDCPH/wShxDkcTVBzzi
jNReTUgnM2dDp3vjL+njjt3CAef1Lm+5KnZ00pB89aIlyMGKBmlKYptJnwocCeGMcUfm6Vf86Lc2
hCx3V3981FtPUST4QJAF6CdGvGYF+fUG1Jqj4azOhvxXDHK5T1i/U13VlTsvdpjtUcZIheJZJ8XR
57+tUoEe889dTnQ2vFgmTPwO+TL2+03eFYasK2EQMbmN8vxYLW4OpYvE17HsnOzpR8qjgifHdGnK
jy/2ahkdeajqyTAWkhy9EtMG8qwz6HUD8NQiAqn6F9NwvSj7EbZx+9TJBIJAIzbcRhWnExO5fnym
ZFySJ6OPuiWGauB4t96rN88+Z8RIwBdBRIhF1eLCHVZexIuxNeQXocx7qLYlTpJnsM2D0REjOnzn
wAZPdQzFyARWpPWGThXM+E1Ry5gBdIs6UiQoqb8VI+6kXPpoPT7ESjzaWcMpWTV27kkV4mfEDoPc
CoBYG7i0mnLFLFUujH6ak/VCVVnPZiMjHsD+O1+iBdcizP2jppjceIkLbSCv5Py/Ab0g0mOT9MAE
qG55hx/N5gHn0cDRLAE2WfttYDz1+8XTQkm/EywKemcqErLN6UZGu6m1CgdsCllkIU5EI82N3lPb
OiOvVlUZRy7OMIodj2wtWavrNbfKwYNMPAvRabki6HpIcjS4OkyhY5urG8m8TBYAyObP/UObK8yC
4/bCegJ9kBWTERnG/OydnpCVct/sXaWUCz9k6g7UHBs35Micg0Aw/tqoQalkV2Iyjd7DewyENgtl
1MFUN838GE4jBCLMKltIXysKkgkI2WV8Vv6STr4X9NOaWe7xDTD6vYRwaEQ9xpEhn3lVpHogR6fj
YOdarQ768YJlzo8aCOF9O1bfZc50Y5UxtfIwUu5pRjc8sBNz3HpdCApiUyXNWY82yFWvlxrI20n6
WEHhN35C6E8p5K/X4LBV8UFGnVmKW4hbik6kg8t5QTYLcEQDoPk1ewZ7yAFclcwfPyh/bQAO247c
8GkX7y5CJxdmeuLZdkvCgJ7pR+YHjcK0nOn80qQMg/CgYPkkWHVLksuoa+isg6qZVGnYGxJpme0e
6g/NUyVYFphUxaRpWfLPShN07FGDwthbt4T5VFu5mr21j5aSjnWxseRQpS4rrzCoXiunHLZs4uyz
CHsYP/5a3hd4/238vesqongDnsA1E4dt+9Jo8xOfuJR7Lhr37MPGqMH4rGExrS9kHFIMEcBGEvoS
EpKZTfEbhnFzm6H+0sh+pvconwgcqpYmv7xrP0a6U0wiWOGgpZcNkXf9AumBWAWl/lKYi1gFptXW
oGSGFtNNY3frELFU+W+AguQM4JQZC2OULrsyytyNQzxqrgR2O62wEHMjDOeGVYB5CGL8J4YBUUA0
14Zf0zVgp2709xxwvyC2bIZUCeOTfkSJgcKlW6naVbLH1J1PioCqS2079RFusGeYly22C/2G5S8g
f1SPi+iA7bAQrxhjqWm8NrKAOpRqtaQLUh2kUv+oOrRf+bTB3j18nooWqPxgUcZxcTcoYOzS6psF
kV0eFHaRuWi+cdWIi3ENKX26Q56DkTSobuQlwg9sZmctF8FIJmSv6jGYOeAM1kqE0O1muOQC183C
XmpAuv/RHx4eKXIA4bNJzmq8GDsXtd5BYT3Aa29MlXGYz8koMovT9UOMFEJjT7mJOhG2NAs1xPEx
U2bVXuDboxyffi0zAQsHG+I9NA5A4Z8qJ9VkbOSvOxNhMmLhL6qDGFGYiz3NKNxxfgIuTupx7s76
0pY6oBPhRx5JTSWR/mv+NUbMH8B6YfLvmRJotbk/rwuoBvL/NOzz0AFzhSjoewGzhxcfFC2toBv8
t84XmTRUO/6l4n6PSIJhFSvegO4vybcSCgOxCuHu+xO4J4ykbVzgzJ122jYkZkqePpleqbuSffJd
jvE/AYB8fb2AN8FGfDOReHoZjOEkmDgbVuqAxY9FLqc9ooV9q6S5CowKfpMXz5dFeR4nMWB1iZHP
5AukBH/SgUnTOOLAKVjloc5dZOKVsGXGH0Hiy7kLj1/i6LlwDdQPfJWiJgv0rc1agK9sBVaOT9aQ
o8HCr6mYZgzSJtt2uGVCLrJlN4kpYk8NyX9KFe+vE2zI4GcAZH5vdsbbJigljif+d90y3AlP4gcZ
elxJetXsq5OKci1wfvduQsuWKpiR9nVlO3IWOXyJ7IrhLRS3wMn6XyJS+OmujwJ3Upj84oB248V+
uQGhYXhczzRGNCKE575OE2KlKK6uI7rtUY/2vh43z3dbzogpxxqYF+12yijB7FN7vXY02PIcHFFT
tS940jpysMjLeSAk4Yz6BENZVFO352HMc+B9rkOkSpEeswbA4CZh5cyNrYpb5aOAIvQg1GM1nKRq
r1xghsf3sqStLXeiXIz4A0rt6tvsbGRLtEL2Vv2hmHE96Z6lTt2QUbNGutOVVCK+r+vXRui/4+ux
uba9zeUlVj/5EtV7oZcBjdnIX2BMzfqYFn0+9sUw95xYptBBx5ys9H8E9yrh8V4zbyITUiKbNdhe
dh617wPknIaN0wxKoZJIzXFBFn80pVLYgAuXPiydq0ljzJBPhS1ZMDteApVO5UQn6nSJnOgVONQq
i17hNkQQEvNNjjn2uC0u/p91pGo77AT1NawgrIAOHBb4+YYrvP/jKG0YUa6PB9qcSLsC32Q+SNuQ
/71cwgC4hZcf5EGkT1maYTWeNBDk2q3B7pNij0QRAVogOX8J4m4fAfL8VzqlMrGTg5XMp5TdNqJv
i6vwsMj3W1NPuHQQHqUpbdHzFgKc8rABTMd08YAAUi5/QZi2DyuAbqnkrAQUnAlcWev57S4W3Lgw
nji1zStBtusqyWLKf88YLqhfya8LWJl1FUL60l6F4phFO/MamPbS4hdOWjQUQZ4Wysc7RWBX7YbY
0YfdncliaIMlOFQ4y3UqJmNk1eXOo8YN7TsHV7/vJhXRqaeFa6EDKV/XHew6DvBvR3bQw4p5cPJ+
QaC59lHjEDPhjrD6o88tNmXqTHPFp5VVo5gZ33lThVpq3zhiHN7lTkJP06zARUtryysq/51qRCmH
/Nvu1xwHrZPEgTDuMZY//1F4eCB+ij2acELpKjIn61jbtL4rZqV28c0adEh6nc4bGY/wACwnpuua
h4TnJ48oeNFGA6ikvYDeRaJsLV3bXo/iOYVjJUZMAqE3NICuw+/2jl9Xf46B6efgWOHsDKdD0Vdr
HgG0FR3iyFWgEQwphEqM4xm1HoEYw9JoKX4XwiEZ87HZJl+CbAornbbpbpXPyFkpWDDjigpVGNMY
JUdMRE6MYAxuDHBSUQQvnCsfD1NfHo9F7OiTuKQ1xRuU2QsWws8W2CWdx8TPxTRoigWeCNO2xpul
f0wzgdDWKWLdm6BgsprDnPkELJrtZO7oxnDtdhIKTTnU5ke5/e70bU6iWD1rlG5VwkMfFojD+5wQ
i6ydQAFAH54k6auheb8/8cf/mrcpQS9WSdWR2DiTRVZbN2yGJQDJgBq4oRd0m5ftstPGcSaj/NXx
WmX2GAVf0gRkSKjZ292WXTqCaUPuQ0oO3u0O/gwd+qTUbMrn46fsR6e0Al4+OMnFT8j19EWdLHQ6
EiU5h/gCanPBZDF1fZK1s/BUXwCYR9S6N3L27DByEnkSwSRam8UZl7pMHCWUOF8/7C/tROhiv//2
evEWf+qca6SXH4nckkpRsI+e9uX98Y5vn8fxRje2tEc5yvMfZ33y3AYRY0j9/bbNQYqc1Qh1E8PN
usGeuxg4oacO3BaQLjcHQEKlBNtKFlAsG18rlhvLO4UxWNsGhJ5hrUcqh093HzKNf+sFczMaIZjv
oB0LoXqYnawoZZGRiq8QfFQRINrn9qBFjpmRDEqwnVC+Kl7jQhKNNo5IbhdgHx1KtB09Jwmnm2V5
7cxGks0HpGV/5i8Ds0zz0LaVoRi3vIswjQfJv6mRHQGEgDS90qkk69ieWn4m49MQEsFrakqi1WCn
WrytxPJVRAIZjPEGfpn4knPXYcfJE1+6MNzlOd9rJVUz+/sI4rLCk5uDHmOYXPs5joqwqIsMyy6J
YChpGPiDu7rf63kBJmZ1uhNncRAITJQpAYJ1+AgXXP7uFbXvp5knvAYP0SwobktCGABnq7doEBTR
EzNh7VK4Vggx8PU9CUqoQ5n7nBYsGwFIVeI/OpWjuGZUuzMPsgMsMb2wGwO5ymz6+UZHZ0/oMcqd
Z7gfDEw6x5C+ESWe2J9b2mUX6dNHSajRS7XxBtyyGuGlrBvntcIdFviT4OOnV8Ya4wGsHXKq7ttv
8Tc+0yi1McjBAtvCYegLcFUwuYT/hxAinMm2dgsU0cYbgdMiMuN1qO66UjiCyKKP7XyDkpmZIFpx
kGI1cFhcKkMpiJA0H9A/m1yv/VpsjG3L8RDgx/M1OC6PR7asLqNIjdBqXPFjcGx+GOB91ts/qpdz
MVB59b9L1H6TTT+UfzwLs9VtybePe99UfIlBBcT5QYvTE5qYm7Kzql1XVTJ5gQhyTW7TW0xjQc5i
fTTIPHvymVey0dkulE0wVzD65iEa/WwxsX6WfNXoCxS/kCSgYBlk4bwiad3ziUq1m141uR27zHeQ
q84701WUti/YZmAyurDFqd3aiUUIP+Cm9m9EBz/O+wFT3vIe5TcPaMyAiSVDg7bLESPUkR1+YNv8
J490ZCleLV7LHnI+yWpc7HAkQcmaw/eKQFzAK9F916O4DxExJ0TEyL/mxXCiBUQwV3+BjiyqzoGr
4U0b0v1FX3yjD/5GSbibQK4bJ+nocbuG6T1uPfufHXoHRKqMzE/NFBu6m0dnjy3vd90ErTFxEE2f
b6SGOgLg35gmSY0Txz3Kr9EQlG+IqFt164f7Fb5Nw/um0pEidKHqoEHZA6YWcbRakZPafDp6QTJk
TdGS98EWtO/UBo8j7f7coGSpn4ZD7So5Ym2Lo7aajbAv+wmXK0c95Xl5HyG53ZgLfvb7ylt8cbzn
91b3vBkJaCd+dYuwwXhONDA1DdtOoeqVSsbwZNSBJvx77a0B1DfdGWUJspuzKbobuRYRwJn9YRTj
UonRn0KuBO528MjSyGYcCmvDoX9kEGU0+c9JEdB5VBfD50wnx5qznzQxWTc46PQCoBCNLGvBkeFE
0L84Q73fD9lBik75z5T8q0c+9oCmelNXqWLXSEs5lSXMvYPG3urqbj55oX6ln3DmBvnZny+88qXn
toLP7jPugaqaT2bP9Syd75Wfb9Cr3didYyhCau3836maYcFstRAvPM1lyZyVpgdgb2pRK8XfxR7c
zKJFtdWXmXQya2M2tq6iaeQyy1nLs6lGuqn8Ne+iplNA5/GVmkN9N8ywV0W0u+8Jlg2Td02QT/69
39DZs77bxhgeyZBj6wYy/h/GAn7nwnQFKr870XBSCPNlE/crzBh/ua+uNKGV5csolECH49Okr5j4
apO7SkUZltQynsTNw1HdSmHS2rEn0ZmWdeelaRRuvwpHGEXhhs1PcEYDy8wm2owcYRwNWNU6XjBl
t09c1cCuHymKHeN+A+ovIRwPq5pSjbye3s55w7qxaQoZ61s4g/IjY2+AcdrieChtS2rvtpAXqXOo
5N7NDaLlkfoROFKk17qpW2D0s3dgW5YHb0g0L11yhhZABJZEGrLTheAjCrbZ8kVYHj/voQx+ZT7q
YrsVtrpW81zVMf3ye2qBGujFMleFFtOmuPvDWtN+WYDO32sgylm27oR1q9cZDoRsPuXSK0dXSpFo
2IEsjyTDwaHT54edk+9fb+hxg2agymQCsE4AQigSI76IwC/cMbd2rP3pg/BbJV+BB0BQQ8bCvH4r
eWB4yb5NDA5wbbDa6xBggnGQwvpzSCZEvjLivc5/CJ+AgAyVJPIPgjwfyaUMHBFmlnUg3WP1c+KT
f1afcBmDOE7mvN4hUdYzIPYNZSbne7CKkr5MHlinzMGfSAwq5/i85CshDG93Fjph49JEqb2zmwWC
EhZ3nDVChcodwklzPk/vG0AQkYm96+ZdWRCX+yB6QBJciHhTZFyMUsUybdNSs6iKJJIww8V36p/a
IgdMgg3/NhxjYd/mIjU+3VTxFcOENbWE1Df7PlYxn5nA0reJXp0Z9bK3WRG3snl6zu6CtXXz4fA/
3KGQC8HLhoOTY8KCF+t8pG092egK+y/571vloUz/QTQK0N7BKNlLtiNk1DsbGqHeqkI79Qz8XBDm
s8ll03I8q7jBSNML6NhEgPlQMaxHDmJtcO+4YPW4bamwNUXAO6zv2bxat6Kv4D25ueEKtWZ/qnVP
/7+ev61ipTk3iBXxIdeDyHXTP4crKYYbSUIDIGF/T18+RwCjBc6opoc69PX1ybi5e8c/RZZAGciW
6idZ+fAonooDl/UrYpvWmSCSnOQxtqgrhI3qD3gzgrb9Ed8txzvsTk2TjnBJIyc4eCeqzXosUph6
fn8zL4zAtGg7sttLeKp7oBX2NEwnNdp6kNUPfKCgTgWG33tcteYcM3z/+2xpgFr/xGuSl40Il/vW
rCxPuFj6mXNHYXETpnBlME9i8Wq9ThTIxr4j6S+aSIk3wkVCuaUwoXTenrXw1rCSZq74OwbN1ks3
G2HBRg5dDBplUr9vhuttgoU6mjoeO6n6Q33go4+InqbSZK6Ktdsh6f5FXJChCoIPin3hs62anOpm
hOgODYsWXCUgj/vJa0aXfW6ZPYl0kX8B3rH/tQiS0XX9bFNskm3gO0psZZP4Pdw1Plj/YoZEzwlq
Nz2TyErbjBOlBDhjA+8ortMKwxgU3DpTFHADDZ/FN++5IClcgEq5p9demOT/H33g0PwIsAJzWE07
/DuTIRJaw7eFZ7nl3tW0b/Fkq4Bi8TgYzStrsrl4n0/wxw7jxQ0aC5emge1UsoqT6hv5ZIi+Zu1K
nVVCGfpnl+jA/a9hmuwGMihIGcE2irFRUOaqMqmco5fdnZIqliz2wiNAGuvLYl4xAE/LwU35orij
0gCocB4mpQrZb4sOdU28s/4WYTqpnUeyGZq2IP/s/zviC34svAlyGdVzGsFwO7/9RkqF6AEXbzxi
K6aJ/qmFzdeg/8UJN1CMgLCsz4Xqxt/KfQC9yFMofKu9eaTW5Y1gpzSaKruUf8shzLVL37COx/2C
jv7+9Ca5Tl8LiZV2yhm77ZSwsDxtWuwlGELWFUal9fufmGyWi6w238hmkba40ttPtK+VUetnyCiJ
al4pObXDifSQLjkgCrHxZh3KFrC6jm7O98rE1pArE95uLrzs9X4QXrsMERrSm5+PSuE1kdDHMY5d
AU6G8Krd3ZGTt1oned6Av/1nGRwMR4QRI0VW8n8KZ6mBJ1RrdMH03f6HtiH9m1boTBpewWNv12Xy
42r4mwGsP6IeCqDvMmxRIS0ZDX2BuuCWk4Yd/d3XuujdXpFrETOBvM7tvKiADdfdolq3ErmwPxqN
utrAlnE+/OB80fTfnWx3wMjiOgwojhaCeBuMkRmh+4wejGP64YYMZRerXzqUYrMSqD2MQnPJYZD2
XskIM9npOgKrt+RQMb6gCqu63KQNauDUHDRy43MBcLh4oTwSbr0fm7NEtaKsjdUcw8ETRmTs44Rs
EkETV9j3XMyYrPJpQueORFddSkDzHcwj6NF0XC6q9aDc1QBH4WQTQ5V8eqR99AyWMUM7IDskqAkx
gER2DlGKUxmFcG4diuB92jKDUopRFDdkwwm68Lu9D9xrmor0xWyXJ0wb+IMwnG6YVwW6vOOR7N+v
TcX4oAx7TFd9jJaZU8qHwp2dINJ83S/Prdlt0/v3kCrJgodI6r1KQpkK5x32VJcF4AzO6I9q8S/b
Lg/I3bSolyi6YZKLmP6Fcyux5Tt7Ytyz3+Rfu9gEEkJ9u7595C61/WjvwedX66nb9jW4xzN0emnS
bReHEjagraiCg057hp5JKdmhhqKMd7YXxEUDWZVddZtEvfH87lMvv7lWX4/yQ0e8aaMmDR8gmrNE
UkImCdl6LiHPxqXPnld3YOaJbO8j8FdxjYY3QoLIbkC3VxjcArCCzOVUcDlmzhWM4VXQhWivv3YS
6n4vqfVv61p0gmyyI7dXTQLZnYdQfq9H6facZ//nx1jPVc+Uc57lO8bRpizevUu9f2keF307gbuY
zlhQOZ+dVe4C0M+Sj/Tt2wIXu0uyImNGU8mtJ+Iha8uAM2dseCWSBV4fz1GIHA4EjC+RuJ0/Fk1I
6Ne02HujUmuajSL50Jb6swz83JEW/na0twFjSQ40m0vhjF9SsDaQPoDfAG2XCvo8cFF3UnVZL9Vs
UBtJaANQDI2EZkSN0K1lCoKCe0CvdmCMAwoa2RT412CgykuxuN/2NcxlehtG9fmpyK0h+DBXX2Y2
LOgUry646EEfmvFFyfWQrBEqYm7Y0qdVlhjc20njAU77G/kuA6SPuRr9EyAJA7Z4xHyHjvrWiMrj
8cr2Oh7UiyOeHPOxZgaoOGlQo6jCUuEEnfqsi1j2SkMu/kSO7m2frtHMI22psQNNbFqWJ1DwkUX5
1LTLlRH2ntRZ33gF/X3H7DrtKLk0a9rHRUUQIf9yOZTfwUYZPRxsUGnr1KZ1ezY8BeuPOq/iXC7w
P4ZFQqVVHv5F9d+5IYHL5Z226nZhDFCKFAgTtSvanTft8lfPQFGADTG8TfRcqdM1i4c5o8oALgGh
+F1tQUFdTcZadTF1yN8Q15VPLijo/yAGxg6RZkwF/WfLR6jJ4rQBxmawpsc6L6gdzWHdwqczc8d0
shU8nGGZ7X3aDzF+kOdAoOFAoACBXoJELWltJU7foK1puIHAPtjJLjksLERE1XDjFVr4EG7QkiFw
R+3RsdBqTqw+2VYSMw7AqVg6zGx6FookEL7Id+A88iZqivP3SvibpBb0pgypnr+TGTa2yxIRVcQk
wrIjp8iDu35U3kGuX6IU0TFp/zR6+0KGJHtw+2O8u0AKsNwBsqse1sFthOi6KgNku5RtDxyQiiQe
epnQKZeVLBTNavyHbAxB7wIakn7iRRyhoHT6fNT+W69evQr3auvNK0vxqHBcpGqFXit5eYvydB26
hPPQeYKNxte/oWCFdxKYGHPVQmlKxUsj9AVFlc94ar936Xe+ML/5HnqhhJmWG1kiVZHgfv3Nelc6
NnF3nOmXqiqycV+Gf7qOmtg3xE5iRMPrr4oWyPgNmAUkvh/t1exAbpfSwWaSpcXbgGjObAC98lVc
Vffg7ehVe+uuErMIPrTjTKBq/Uyl7o5GvZK1DJuvi7iX2ET9Wb2nN+oTGarTm1i8JW7SW1mgkk2k
YMPVDTk5w7ZuzXJ8S2uTKhG5qP7ueHGnIMiztcSLVipDfZqvbQf9Oj+oA1BNP3UCc36w8wqwl7aO
3xEsKdr3k73DPRy6J0G2BMgv9gVPjH9lv4LR2KBH30vRyXKcVcS2Wut0hoVrZQRa26tuQKqety2S
i3LWCoUqP3Y7/H32eOcxXoG5TUxeeGKn+4h+OoIxV4q5hA9WBTjxBPKG+ZzsHTK/EdvcQpIJt2em
0Hk65y5NbydC//5+ZFk/LiIAzo9ZrB7LZpoXVMxO1vX9LxDIRHkgYQ6dqAUivhavNpjP1wD0ayo5
MElUluz2Gu1+dWNfehEnk3nSI73Tc1S1D0CV/qqxUUUn+XMafIL4sAB9UG1i9OJtDqENsMjaOJG+
kr2DYVkZuXh3449/q3pVV2TaZeDk7a6TyFCD1D3SpRM/EqLK0UehGibK8m3ebbf0cqE2ZfrqXhrt
hDgRGn3LuradLeEi6g2IIJ1QG2Ypq5xsxPxAihq6gFybDJHvivuZoVYjKxeo99ungbMvqwZQwgc6
rM0rxQ1/5MioaSKvctj4/EZHVQrIGpdqbotxDtKGVhUVV2hlmZSEJ5tcE9vGDgX1zx6AZ6zqNzqz
6PfK4STYAHFMLZh1SFUZllw6z4LPYLX4+x2NsQOOJb/GrKalsLwLmKyAMAJuvi/rEFikxbJXc0AD
WjqC387ipPXHiOMxwYZKHk1eAgsx2zdbdHJw1V/YFnoaJ9OW9JBXRwI3bsnwOKvR6kwIeSwDlC/r
6MJN+KjGIVTA4hI1itnXW0oQQ972zsnw4ZR56JoKqCMmNMmYyHeURu2HgVyjf/p75ARe6+oh3zG/
rg4t6JvTf7S2yQDLdFlJTADMC7h0cO9gbyIF+YGND/IoBbK+dnWSUNcUePgct9CuKhFV+wnkQCNa
rc2A7M+T/NNMX4FrUZONbsMXovq+3BKc73dG3+GI5T8UWS9TvyAzkRMrsjn2e960VuIlwC7wSYm9
ae/AyJx8ngRAVg9Z3kLz2Dkkn11gNK8G5mGdhZEGHi40dF8VBzw8YqITpyNJuaZ4jiVWxaeNUPJe
LLaGdIt28eobFS6xbTPhiR4ff7ThkBvaW291X/xEUIbhDtmzM9Tl2hKZH0ooS+QICZcaPGzDGl23
gxdD1iIATyiiC1dM5UjO01qoEImi6qg8lVx7biCEIgq7wYp54wFKwq9A72K5vb7tTTCAWU4dze+k
Hod7UwRl5zrPL2TYoWHjQ6vsLyJWvPJTdZdK4lkHEWXYiHzKXl6+P08eXzNBPpWSM5RU1T1qvSuw
LTw+RmzlW0PYb7HytVq4v5X6Np/+9GwcmT0IYtwdtpsNkcBMAKl2gzW9wnrWh3NonFMIiFA0lB8A
FmHwPi+VNbJwNCOyViXnIHWWjtvZFqTmNPmejbz7aRvTP1AIAzLHauzQkDXFgw0m6puryS9pNfFe
YYo03JUHy22p+O//U0Kw3Ndz6ifqPOgnnxBcaZVxUV6NXUcnqQ6luBnjh2GIZhTMisHS67hVB6Ar
py4wGroPVOJrYi2fYZQxPVX1W+tXFwixKeIjE7THwbk8vMXSLhjr4bzFaIslktiOaVrkEqa0V57V
6w70YhDWdVqyijrN+EHWznxORlcJotP9irLNmJUOFf+wNUFnT2sPqqPVWZymEXxbcnl/8poPA7FE
Nz1FvqKIyDz3AR15Mdlm3J1vQBd0UASx8+nHX2DHXEJMZGXhyGxva4CXXMS0mVAV/yn2RlssFw+u
KkPqrVzpYa6bKNgCJlFiX4vfoo2HmkuqslGeKNNQnva+swVhTfW/6/p965WBLNvDI35cUZKD6MIq
AYg2ySEQwShrCrZz2VqgFs5B4LFZzkLFl5RITBvdiH6Ts/cW/EiT/niw+K7KP9IKwOETHO/VD9GD
OlCR9F+2FMOBk1zhpepY6P5OfIO59SLr8KrZOF02dfQWfcHUxTqM1ySf8gPCOWlLsnQy8SGqBmJE
OepmwC9/oGZx3h8QU0KqdGpvu+Z2koyuN4WjZ+Zfjr2sfGk9kUov9mV/mjWNwBBmybnc6O0u5gg4
3bFFHEbCaiWTNi6IR9dtik/KwiSKsqfoN/fJLDcb9XIPokKM3ZpPwIh9+rpvhpY6aLUcvc8DDL2/
sRDJksjwcSFZJJ0oOpHIAIQ3XAXxHDQEeFZ4RU0zlfhLzesw/RMtBDqAB/kQjks3jJ89iovuoZee
JUFY8gya2s03SyZ6VzneIiy/0qMf0IgNFYJBaEDKzXII6N72PoKzyHr45blx9Ye3IW6KzKArrlD/
Ud+oDzkmE418R5DL+J2DQw0br/3PLfhIqXl9v0kB1TgWpDazIG29DKXPkeeAmdxZ5gskQxiSW7a9
BW55zgTv2U2RoG7FW+zVJq/3T8KOe0JNWX1XxzxOwP3FQKJ5WnEE/EmxpIcQFFs5GXuJGpEXJ85R
3/Tk8QxCJADz7DK15q1xAsEC9sZf10PVwpaQGEYr6hn69aBVZtDhdOYTSRcvrgGoHJawmUD/W1W8
gwpFVUp5x0hzrq/TWlA5zYGF9Sny2eRwKooOXOI4l9BTVqBXYAFQPlNZN6UKl/l0AyY8ba1hQ5O/
x8l1siNprm/AyRsfHody0NQQ9w8Qu1G67Lu/5++jYxyRfgHRJMv5CX3Q66Su/PRcCIaHxRYxVPjr
ZERb/9NGzrgz1Ib6rs4zu8i9kUsvZlyq1unVVSlqawvORm+iDsmWuzgaCWaFJZXsRAu2j6hO+LaC
srHGm/NI441hzSFqydOPqMV3ta/1baNp71CbUq0FgqZqtEfupltIHWW5DZ2+I1Y3UmiVW8PuH326
uhEwm+LNkyOjkUr2e5R1B7WAElueQy27gP/S6IbDnjJmpUkgDXIRHj5dkkM6mVa4zdlF0u/qxDzB
vjgOg2IZS6PCn1Btsu7mHTAv65YkgNbpsuMZLFYxeI++wCDJj+srNz1LM0wvquY8L1zXNKmWcn3+
nqp7ynBHijZE+ONVnEr0xMmfveX9FV3DYo2/EEKA9c9691TOzsAi12Qnr7s1LIWgCYazJAgyzRKh
E4Oz1VOC3q+w9E7dzUpXMVWof7PArh2m3m2q5CptfTB+W/tBnANdzv7QyrqlP0eYPU1V8j2BoDlC
Jxr54rLYlkFph6vIDbiXK0n7ZuBZVAHIvhAXnbzioIyyV5c+8w+gAuRmzP652cuNounh+jkSVhPf
qLEWbqHum7UtYhWhD7rzeFFBBfRXUkCWknlgOQRR6bjiwULe+lskdC5laRP3LWDfUAI2MUYsQqJn
v3FhnCrsQWIP86kwx1yoWIYD7okHMxPh0+zPbjlk1rAPYpVJDhCa3SLSDaOdWj/AufhqabF56u3k
hMncD2yP8nvjp3kx3epekd9RQ9Cr98IUjdf0xlVx2KCCrMJRoYKfiu2GhmARA/S1LVdm+1lFuMjf
LRcs1QwynlnJhWehEWf7PUJN2wS8t3VVX2rUmOrRi/s/o/8yrpleWPT/WE5cdLq8M+hhDFuObDkc
5jPj5yxr2hvHMqo+Yp9daF38UIy00XhHES8vIpVLHgbuUUqUZLnL48QAqScBAN5TBORc7mHXYz06
MHYvrKYrwbmqF1DRYafS81EULw8VirivhjTMpljAXx5PO5kLKcZ+qiqdwt3d0XcpfdjjJ/7phOBl
YOtCynbH6f21FcaDKZAs2mOs6FF8uIFJKWGT3L/xzfhL1ZRyxoKq0TUUDi8hFAgXkk/jMHfLVdKI
6UlG6A12WMUUWDxyqO2qxucuomy9it17LzPKMbp1VlzNic45RidSpWXX0QYi2ZKGSLMa2YzeYbkB
RfcgodxLjcXKbFHEILUbk+isurXNFuOjU83P8tFJ3MIMGIU540xgsdt8U9W6XYcdVfwgXalf1ibK
oBQkZnR7aa5d8OBiq3BY4UhIr7DmD/iR5E8SgBPQ3yuFZ2u/nsJSzB2tZmjIWzz+aXXkUC+6X0p5
SOEBfSLOCXaX2yKoL5GNzOpHlu78Ly8IMTbJJ+DY07CgMG2nAfvWCQyTpmmtW4Pss4lXXjG/cxIn
CA3U9ZKKofXb7BcF2FlnsMv4FZVVc5DX3s7+O/wdJobRlioXjA2qKLbDYmSPn7TcFeqR1d11ojBM
dqb5Ra6TWP/rpzBwKDj8rLkioR3NcQRUBciigCa/iIgMihQCAOV30+rnmaoYMdZtx5GC6/xevMyy
bQeyTEbg7xYE5Q8qm7O1D/WrutYUeKA9heDNeFw/0fV5rWf4tw/CCE9sgVTqMbkoxrUl4WI0iMPU
tWQcMt++qDNB1xid/YoKySPltR/2rzD3fQB4pd645MEXg3WbGY3PWni8bitMv0Y6EME5ODdlQUba
wptjE6PHphcn+8Btwuu6cEf9aJpKjC5WJLuWnCPclN0F6QJetmH+5XSQKhUwc6H0Q9PK3lCEVqMv
vqMNtjm4vt9HLmBFG5jOnJxku2Pg9czEXdNUWJr7kUTe2KjKsMqEfI4JTR1vhBskoTR0o3m6KSqm
lWR8IFPBr4ESb6mMQLDRcVEm8nU/wmLGDCrYdgsr++aLsGluifRa1aZ4gEd9p6BcmaWjdUpBch8r
1+R7c75zWCR30x8VQ2tPaUs8z1KC03Mv/tiHAeeQP5OUmWwkorTtbZHGT7X+9hLns/GiLSouRYX8
/Y4tsFQJRndVfaS9auoyXvPBQAtQm1Vwy/IZSovds/29WVxNnKOb0wngJQWg8D+QsgIkRZvrY+1t
I9atNhE/PPL1TzajaQs7tAOlK6xgM1Jmpk96zr73UK7PNvA7N3jB4FnlSlvmYUXiGoT0p2Q0Ulu/
VmeJFnF8k07YAVQ0mFhPt5gfowB9OPTyjPSIUBFILZoHzjnRc2AAxDR9GE1US4WDWt56m3uWPo0j
Xx4RrwyJWxzP0vFdOVEwj9BXU7AwdtitiUVB9y6awKg65NqIeTs0uH6UGV53Qtzrs4EYwccyxQCY
faWk04MbUo++dlVpR2E6/fZkbN5cGdw66logpsmmVVes5wtSyoWFsnuc65HzGL1wqTcSr3lQzBAM
Mc9acg0LLDukdtyseoLkHS01eCkekjY+7zs5r5CQuASJ5beqkshXeoQwWZMvS47i7RGX6YX+YQwf
r/jqKT72wsgR361ycbOeHmBu8Yls6M+dIkfRkuE1HdG+sRyqlVPjDe/j6SElnfGS7WvNO2lk32ot
mIRc6TYpzmXJqPVNPZuexvRUZN5AfwxyO1/piV3DWAdJusWq2Xs0hhjYiMZIQ1AItBbNVFEUh0W3
0K87wIYYAFaWKamou70nILClodffhhzR3zzmcQ/Wj3GD8MwCJw2SjGhAJNT9iD/SWzXHnqm6mUxc
bzm77YZBA1CURzGSvKMLSvh4yq5RuaUi/13Nf5tZZnQcHs6oiJHjfII2+cga8ZGv5RnkmMj3iwlG
2wlQE/E9AIhGmo1iyOB2CQGmvBLikp8hb9TFlUulDTXbqG36TCjqlXXxA51QE3nvZoirToQCmR7a
bWMQ+xtZXYQ7pDl2NZqiOpF2EPPqQegAFnb3W25WkdDpZpRGn8q0kFDEIjSKU2wLMhZPvCqgYJWX
Q2oQv9x2TSpUJ+wlTk4mT7szSnzi73AyBb7rkq2hSMXUST2Vlxb8ILisNQW7E6Gdouyo/LME43A4
wifzxJlw9LnnxPib7WiIpFEXTLWl5Foq6KdUBz5JI66CCiZ/ffYmbd5UwT2IybDmRngzLvQ1hIft
fIsN3p3arF3Ja90Eei/Bi7sInMzAPar+BqcdiM6aUknp014HSbbfugwtGjpNtT4g+SjN7yYjfwv1
Plt9YFFX+gdPHCqYYDGL3K4vjGqC0q5bNewynuq4YsvmYVQZCGpBxemsTwEqX9KQ01D3MDrB6GqH
q1AgQcjhPdZbF79VvQ/rUOZLCS2XOcgOT1iX31HYvqMYmdEL/vDrWYhKvzLVCYdnlhEt59KyiGGr
lwErAZdsw17USFT1TzHiG5GSppkTOx8Kfe43c35oS09OskVcumAjX0l8PqByIKdRPRXf6XTpN7nj
jvEvx7ov1K82wyjrxX3MGxtznwDLmbM5J0fWe7LLAIhJFxahHF68PDvKfLl63tLrhIY4Cj8h5gCc
WuKoN0BHS8TaYTFXZ5Csb5yZU43mZGnu829uQ9nvjgtzUu278sNa+Xfte4+1/B/9cgKIGl2H20Hz
Dkla+uJiF0I2UqflY9kfL8DKXy0/n9e5sLsgsR0I1tm0ZxIPs6FdY316clZujC4CJr2ZjY4cIJSx
osvO2pW6SsI2gYhP8cD3f5h1Si53ykF825V+3IDxAYuhanVoyG2Llb8OdXDWIqblTfQ50PJPPQ1r
L13Zi4SA9UYswWk1iNZw4r+5+8oL/V8bF8Ym+ZuZHb+yWkPuO2FUObcLydYNFi0Es730GDDkVux/
yNLpzM8Teaaab/AxdC7qvg6t2Y8pOg2kl66oTjejmqVMQKGGllszP8uiC1re2XUUB7WA7pxfq3ld
9UEcsqMrNfeMH8K0D/s2j4SWh5DK6YFj0OwQGUZggxfLntji/vYW1w7P5rcmc6O+DhGobgjDkkTy
Spxq6xz9GudD/+8hI3kIL/UCNcRWlMe+8whuGEbd+XgPjyYgpHVy7mlhCLpJEiNiiSpSamd83RyX
kDc0AMRPPIwNyUOcNI132lU9Uux3JLGwXeowZMMlV8myZab/1jDdesKB9Za7YlqG+uIhoI665S2E
M+/q1gjeXFcUlfd1Cj/BPfH3zlD7Umy7f2/mjXzsXEk+zvwseT+Aq3YMNxdZagK9lpO3PDG8uUn4
KGlWKRzSXsaM8D9RxYI4i6aXbk7UVJTkbb3DK9zdmqX/TSJebywxzKStirA7Hwdk+Qpl+60EnBV1
xPkC2T+fe008eR19StCLPZG99PXka1AQSh1rufmhEcvLqalhR3F3JONJxAhT7jsagivDR3ZVwr5x
e4n5G5uiR+J1srfCE36kPEPes8DNmqtoGZXM9CRM0bko5F8gQUmcBB1Nt6Ow3ZvYrnSWRl2MS5oa
+qQN34ZSW5qp05YMFUMaA25xrt6kFXReVuEHVuzF3BHo4+m7lS75zrGPoNBWiFUVUH/e67RufWuw
3kbC1PGJRa63HIL/rLvv5el/cG370MTE/LC5PZ9XJiNKDJloJZ1Xm7GgDp3dRGjz6e6DdNc4kBXx
0ZbyPyfUy5Awbbmf3iriwL+Vvy9cltCQdZ7bzg2XPhgbF8TTD4O27LaJgvQBRBivJCq6l1ykVGsh
DavOBi3SjvNY3ERyt2S5H7Mw+ykYk5057Dr5vY+o8MkXc5Uld/CvqtLTeij0zAh3zAnr6iES8FG+
oJtrTkGUgqv3K0uhziHUMUDLvdxJDPpvrQLl/QpxaoSGiSG30Lo/YckDajMjic62Yx+l1Z4U7PHa
kIVeJR5wW+RJbMfYpqogfGA8730Bh2u1AsqmOzhm+VnnENqWs9cH/upkqx3zB8CzBNMb9VjnJOr3
unVPcDiYmWzbCgkuf4DVCAmXKv1p0ZXJaRm6nUwumO1FZf1zVrTiVRS6RvJjjWtc1xTtcsjeVbMI
LekN0T/j15HshcWToJGwckuUliO//gdLRhuoxQJe4arQ6To3u4u2Ojg8022gL4TF4cO9pNEctPcS
53bdknFLjVSU5XG7RWAyDR6kaovn54m7wZmwk2TDvAvBU/nSf7S9DrKsap/1AmqZp/EJK079C5qr
WM33RrOmy2EQdl6qlBP3mTqUirFiDGKA/RxCPQls0gJUXaEqfN0yfg9SRIb9bjUMyAoaY7dFn13j
XXpPMKLcV8pSyUU7Z2vI0xbR67eqAeAybzWa1hOCJpLDjiYqYxvEx2pxB9WXOiF3camDjE501kL8
IavVniCR+ly+R4Z/1WDmAeAzkKprw+iXW2tcLAqFpe+NhWK+faKpz5LK+S2NiMa6q29+lJztacAL
h9ETh34gVzibnuJxS3amFs/GdRjhtz3umkiMO6MtpFK7gHDMBcGwZsK+enRGu+7+QO1NSdZ+b9sW
IzButp82nS7VBUewkRKTdcioXQgpE/FM+6CEmbHvur7/xGLNz01JY2KRSUV3DA1u42gGjYpC2WY+
iNN1VOemr6kIMqOKg4PRSg+y65F4ehpupSCn+MC+XA458LNgZ/vcre9JFAd+MYmw126x9LLfbE86
rEU0oJTh48jvMtQE4ZrdO0C2j0V4MWsVdsomKQllY0Rh3HzRnCJWvOn5gDdjYvHoVVmDWEupRNV/
LOKrF1XZCINnzF7yQshKZghOidEYBKgokt0aTsmRvLCaxDerZJ3E8JvtcovrugFNcgQXBnldprle
tajSo/fzJDt1DI/3NgBwAce9QcIW3u8CPCkqxEKUGhwe9SPgyhYjTkSgaiRJG/GQ8gkWL0O91TKv
8cb26au+EgDWNoO7L3F9mMfpTEd+EIKK6Eqkuw7fRJfsX5ztZ2tGLkIdVRYwj1v6TdZIgH8SDug3
AwnRgE4UwCg+V7iPuXuQuwtUShVUjiEYBR0UP9A+vARG6p9ohEBpI74zIvJ8Oz6u1f64eQG5gvEC
Fb6tu9gIFD1t6pnZbCyFgf1Nalpe8diY0UGVuXnJMDPw/Pzz32w2EuYWfWMFWaA8FkovjIOwrcNI
MS3RTuTzpymOekxeW94qhbts2vkWGJBjaFmRCCFocJvFcFApEqjUUHLgps704Bp+Zbx2F27GN280
NSuc6PS8jy5YZQ6lmNBUU84dSz9yLJtPyYFl9hP4tiE1E1r+2q9eu9G5q44Tc9j2O2YHgFF+hjSP
U36mhB5xubdJ8LLSkzSdPsJ29apJoW2y4p9dW3TOiH2b5TSUC9N7TOizLJFKixvQ3zXpAZgDCU77
dYn4oPSsWJtBK3YFZVw/IeitdENgnaVGtTJb4Jwr1g4L3ijzkN+T7ZFJwZAsnPikf9oyc9fcN4cR
37s9yVxhTxJE++8OBAXSyJVwp1E2rBHHTD04GMvwr9zYNZLkeJVLl9UaFbKCMydsHn0hwaRTkC5V
jjelBzKVvypE+LP+YCY9nC5wAIEcsRrQzDw5bA4wLQpwyBKVhTL/J1N7ajrr3wYhvp2TaHCRZq43
rONeG+Jg3i/2Y5ymF4Bjgo81yuVaEHJNjU9zauC06Zmu9SyjdhI/mhqAyilK2vsKMMummjo7W/hB
2y7BbvGhNA6qJBOfflRFutpU4+dyF7UNg/AGRvjfXy0tlZRdwN+mNzoMQ9cPd707EUXvu0/Rxiik
rF50BNfDNasmdNRG7g6iADg046ZmrQ9snrZS9AsYsQibVHU04rNcQ/PC43Hbbk4VMvED6/rnXJtQ
Vjx5wu7/+Fl/wYu9zXOEbcBwO5f020sKRTdkLD6VE0x1Xv8XgNWPtQr3tcASlPIgNwSoHabamZ4B
/hsEWRcomNohnujwmSs1XBJO2vSdaFnym5OBv4llKPSmejIDxDDjBbMXIuvu7zr957phIA6Qt8QA
oPhx4Ee6mQs1AP7KBVHIXUgCZhciXHUeE1gHh6/s/6UTGaNVXkuU8C0blDMJzg/AVuMCRHcd18zE
4MKca+5j9K6f2Cqn8cBnKAji0AKSuR/rRU/Nf8t3+JNlCIe027gJ5um9/IgNHKSPMOVayAbY1Fca
Hl4eCb6vlzmiMeLNplPGY92rhnCYh4CrQ7wvvw4lNO38B1HMW7YHU/Ik/SUAXpJJBQSxp9q8c8Qu
f5Wi0gOXuTxE48H4861pR3GEXYyYwHENr5p6C9A+P3/NP4FJNyMAA1FFlkkniitZOwNB/sNJgDHo
L62NpF7S0fhvtP9r/5sQEQ+Uv6GAeXv9Z8OF6etFLL8ekYByzK8WkQ9kVUCDGuS5stgaex5A4S1g
rFSFd/fb2oOl21BlPZR6Pvy4vpIy2jz9xTkfIspO8Kna4JvtfcV9iw1jWHbQBWGqaXkZjXnMikw+
EMEcr/HeXmQ1tXLx3RlGxxB/rP+GmdeyT6C6U9z+ortaOqW0/iwJYeX+lRJnl9er3w+T5duWNlKM
LHnkD6YwGDxjr3OgN6Sj3C1h+CImVBWnzNJlvwjpaoRoqqhKRInGspSw/wC2B+rrcA/KU25NetPX
l8GoNkd/O5kz0G2u2066IUmIyujw4s2CfXxtZtA8PKRYGal5mVb8g7U85d2aNUF5oR+qZyVi5L7m
FKeCmY1fuWPGasOUIBKUeJ5CPR+ewjTX4NSqhv9O37TTRKKT6/VeXdtszmKPDHFuO72LHE/XboVW
N/PwRN/eLbgalhjPiIwvnOKw30wQ0BZAe624yHA+gNfX23J0a2wUKcLgpCaoWvs5DHzsZ0OJ36Py
TFTZ58PW6auTKaXU2EBJs58ls4k+YTOYDaaAy98GNI73jwls42QxKUzu7pFDfM8QtmSAB89CVdex
yKBY+NrISnbV6XMMbge97Dnrb03HA0laSlNpjdPiwfcIO+wWVnv7AQ/f5D4t3pVt30MkDF/v0sEl
C1WheMds+g2CoRESKEqLCLxiHGUbNkEtXS1ce4aEKPXE6blHVQWDTwqLV/1V7QT+4BpNck7mSMPj
mHqyxfO0f4dgaTYVkbT1+khTyOO8X/UGRobryO2dksDrBRk0AecYOLVIm2Aa186KL+Hhfi/FGZEn
gDjZ3Y5GVoyljjzWl4DmxVtx9TnNBxes4s93eQPKOaaHn3S6vSm0qBjq49N07dl5XwOTu21CaBOZ
tgvwTi9/jRhXlspOLIqSdekPkn1tHIFCPQCwns7rdFnR24EHldvDT444I/1F+CTUzmdMjtbsVNMB
zRh6XD4/uIBl1lQmtTutQIVKH+RIXUBhPPboVR0F0QvAQKJLe3j5nxH6zw1VGPVC+aoMB9rpYrVh
rc6T1EQOfDpERocTPrJmol9S9tfTDdjCuhux6PnydKh10ryD4iVxXSldMYw9pJ0oFyFtuS9+YV4W
JeL0fAIsX5b/WnKTyK3LNXW/HZsyBVqzNvf9LHqPyuxG/qlgYPtKaremiZQ0E08r6YqRuQzQ0p5/
ajoEXKMOg8tkmdYZdZ9z5YOtRV9c5I069sO++Oi/+bJlHYblt70hkQXXTTUFu3+nYVKey/n79VjM
QDV0ggbxAfD+9xdEZSpB92tYGIQSA1Yt+4KutAcpnYEojWQZrvDZcxYnD/otEUOnnw0Eu1wuy9Oz
6juWAwyG25YRpZYLxAW01Rsg153xzcdYlr7FBHmKOBOlwXKFoitCQvjS0wRbiWj/JJwjpD3Lfjux
zTNYHVKGeKIkvlNEY9redR7i5xsvoXWTCQ0VWFrNSoj48Ia2+mbrhhpjXoxvQ7thus+1NTZWIq5A
xgmzHSiNsWMy8Pfu+60ICSUJZTMmTc5xk2KRpXyu4IgVelt7SEIx/Nh45YCcKfOw3cKK4jrAaeKH
0qvEoKnu+hpaBlcYMxSsahw+66QWBXDsb0aPX/mO9snmizQnAxwZcODn5S2Nee2MnuBnIJ7SVn6D
YCQT+CRuMUA8dJ4hSrJubj31T9gm5yanmaUyMZV0R6s3jEhrXKzzu0a5bbNyBcZ9vN9tC6eEM2Ai
5JexP2hCyyvb2j1j8VRhLzhur7ppvmdYvteQLBcSEM1JgZEEPeWYgeR80dPzWvbhg/ruL11TyOTK
WjKBiOEw8bqBERHagmSJZfd0YTypdoAbRtRyCnkkZqCDhXSb19XuB19I/rRaFnaRVtxt6MsCxwG9
IIKvRDRoaxkRs103Umpl6sYxAC3mBhmdNNrIJ/uTNxRXuf2i1yIlcsreNE7+7sIj9MQkgEZwv36Z
OFeW7FNE+H7ST2OQPnMQMotXfT4aKlIBMA8V3vLLLAWAUdOoF98BVHRPs65He5N5Qfj+vkdojz1o
8lw06L7383vqN+/mlVoNHRkuA5w4sjdbgkJtehgClxpNQq4XIN0MW6vl+gnkxje3NZ5heW6Nz29F
Uw3mqRvfSBN+mtg5cv+Og6B1TSF1xLUerHMEy1r3Bqpn3aEeoaxCRUNgq7S6W0T9pLTj01mekumV
U+StIykEY0KNdHKwPdm3BXDDbn5Tzp/Dee/riyne2vzgDIckxzx/LrioFRhddmqJ6C9NpRi9gmIJ
CMEGjZ1xjCpjAyUWPjoRMfzzl25rGjUnBOlBdqpwwr0bQM/JeiI7zbk6NOkkhEyxrNp83WyFEk6O
64toM/S7j3WAtHceKpVTEW75V3vXhgP2Oy1ahZjMDdt8lKYKs0kpyOm63PEVQ6DQBufbcOTAHhwD
cDIkmM8/ituqUZCDqdq9iu9kMBStKWvwP6QvUV8iUDYFM2wBTGR4m5Q71eAEiheaBLqnA+2Vzr3d
eYu0eNQiLLvERlgMB9QYdg40AtNrssNfuixafxYof/5uviW5nE90GQTdE4RoXmwH+P4t6q1IgXLD
ZV13UCD30oAeY4ltgzYsUPtcd82f9GBPCVoRKTPOkEMuo3ghkC+r8Fv+fcXNW6KNdB2nERToma6T
TWc5vWQDCHqxuqj50kMMv1bYk9qXBOvSF2gbLJfqu+aNh81cAot/QizmhJXtMku75ht4d4CXwDTE
VAftBOx3meuvqT5t4yXs5dC8NeMeRAbEnmTwUULVKJXEb+iN2lguIKd69+jznQP3iHZxe8aWPXUJ
pm5h58XgtMUY40Hwalu5TNujMh3aEWZrniS/5cEMILa88oxFWFqRiDUYCzGhv3QkEkiPsibKGwKV
1UY2EemDJ7cb7xq+jUFNY3oPQtCrp78zgpsBxG51RB1+AP1HWtpevQzPSK0EirNDImBv86hOp5Nt
KoUdjSRuzWqP6zKdDPMJWURawUJmHggfWuMpT5pd8YUAR/SyS+uoXATu3H/YLRdmUDwYishdQbkB
HC28T3BNmgjTvc8sk2vN0zaN4fBiT171VeI6xmWYnw1KlGvVd6jPtb2hSVirkc43hHDyoEL40sN/
rDZz9GCoxMV2v7RIaLPZucJMiW9R4BiPbQbzDfvRLuBWnttIb5LT04rYdpgkX4DcF8RKS+laGuRs
Uw6UXk8AwFSb3sOYkf+OAUUSxOVtgxRno6odUpOFAGodr7VOrV3myAgCCBEEkCeCjjckHh79v1Ff
DGUuXg9o1rn7qKmOYeLUn9IM3mi5BY/WKDXws2LgWU/xFxu2RqPQN0oyrlcrAB6aTC26593R+kn2
uh+KUWX1E2P+c4Re/o65wcM+Ugz0SecOUZjbRl0c6w64y4VOPaAdaQ6aaXTed1TahI2594avyePY
lYHNqRrDg71/m5HTPodOSaypPyPKWqaCW9ikbQQg+PEpJR2iLhrsnyxKHFMqOrdwycyhA2Uk9gBW
KY6K/3fr/cE/YXKnNbKCWygowO5zJX/8HPFF/2AJNuWipIJWu7CPMfdS4VZZont8nckUPh8vMCHX
rZ2+9epNJ/1ys9jePQMaukpl29SfqVfjwV7UbF0fcfGU4bY2eZlDz8X9FyOdn7blnRPMQNQ0a1M7
p8md5MuKuoMRWYtvfZpUANdEZhrm0bDbLBJMWMfv0hn55FL3yhJod0STXB123E0/wAIqR+qxHqnE
EYCmIbLB+0M60ZWN5IUPVPq6bRUpZchKG9zeQ7oMRJbHMZeJRqQhPtjl5SdoT9gSVLBt7BItEZYm
Agxh1z/zeXWYUh7Bke3AhWuM4nyN6ukjPVoQ5nmSX4gSDSKUoCW7XPvXkoHFWoMOU3ssWt5shk6w
WOPir3EpPiTiiWjCs1A73BQUiTTm3hJlIf37F6PUok789QKzq0GpQOUbto4nQDHhEq0wAlTpHxrU
fAKZr5hzs/DwDrpjfYUOJiW03h/wyrOHRyQR+i39x1kXASfo2H7nJ5kY8MRI6hgSE6CvAonqq4aB
qI1AsCff24ASwb07pjIdx1EktxmAaVTzbBJ6H9u0NJVQk5x0nfhu0UGzq/9iAGEz9EPsBuAOO59B
k7tSvXttwX0ABmPtMj/9jI+YT4q/THBeR1970bmHqD3ZomL3+I5XQsa36ws8D5hyRXMKkl+mRNZU
QN3Im30+xrq1h2CKnaaFV7C7GRkQx8W98Mt7zsnEk134KW4o3FZRfGnI6CBtySB+8LcQyA5JMjre
gCb/rOz4YZikWfHecdSPLgke5N5NqSGeIPtLW8AfCR8z5nPq0P9SDwDGx1ZJpuWy7GtInh0XSHeH
CAGmY/x+6OyapXD1u6D1xXvzheANxLPmvWWI6cOMlTxHTl6KZWXYgEixZPHTZSK6ZeQqofPMmUfs
aMomUwEnfA8zC1JmNdkHLkLh/3sD675z8lKe3WkwJT+idKGu2kiS0aJrQmTJyX1cWVeS2pGfeqri
5aY0015lxUkdfpUM1rh/a1o+rkWRtjyEGuq0xbGanzE4wiEGm9F2EbCuQTM943W6HQRMWj+O3OMX
Lu2nE4Y+E4TUPyMnmexZG3hdYfmOA26WDmRLipDRbDhOFrBWbYyWJF3CKPTGnm0aORinDyGT+XdH
7SuzwT9lL8qadwCzDcZ5SzEqDqLYHUrcjxPXdtjj4njMRPeIiAdviwZ9m9ZYvxtvTA7h5m/1NKn5
1+ex5D2yjn+FTDZyp5nkHjOebPInpsmNRku8C9eCyX/0qk3Qpr8RVooyrK2UiCZVe9ltYkapRvcS
wsUfdrjcXjIFMT3GAiCCjpp5cEcVjfaowvduSeApNa/xNDZQlD5zX5bvveTLvbtc+X8PYxg9qxbf
wp0DJCmjTcxJXJXzWwSlSIRB4ofViA2UtxQivzO4oUFJTR+Nzae97nBd5pT8WiTCNOqP9dFJBcym
Y6aC21siDN69p4B/YC41fa8DAeJeJRiuoh9WMOttt5wngUaFsFDhkb2QZGlyqZXxM84bGz5iA1WH
uUM2lSL6+VEMLd+Cm+PiXODWQArrxy9k7w0Ke1rvKA6yH3qEN4FBu9dQ1OY7N6skQdum9NT3p1cc
nS8w5jtUI297WUq8mxlHFEu7BcVu/Iw2jib41K2wHjUkKGGkong9X3E2vhBWPjg6BijAOfX72tZc
OzsGGxwm+TSwQOcbaZpnA7GHY5cWTYIITwgIiQbhXXGJY3AsFZ4sMnl9v9E9CqCbcGGSTVBbifC2
1r1Q8Mndcfq+3P759s46VynUyNIVBHFWef32w179IPjMhxro0cYSJLkJdZJk5f1BKsmBkx8YwnTU
svj0HMIAbKFip3aX393TjFLK+tRN9b6HpgtGZU1bTyxrUVvQkeeXoscNVuyhwfj0Kb91/egbWUeu
XmDCSTllNCgKX5ynt1IhP1qCzun+3nTe3gJsuD4vf5R7wWqWO+HN6LqhJhaDcKfpjrRqcUIUdw2a
yFK7uTjP3yyIoW0Uvyeab8aLXKBuPUTNg7QEgszi0dJ6MGr9VSZV0UxnTb78sg/Dvs3gfj4pnz1K
GIuIiveTpUsgIYzTHLZG6FD8KCq9+o2l4IlZFFfaRGGmLrFWJjk+RB+7EueeOAOfs8eYCXo9oV8O
dSV4oNyWjSzTmR7uxHYnrqHU8RJ2WfV0vBTMHIi9NM++VuLTqe5gZbfYiqU96zXlmxZljpaMbNks
EIU9FLqSDHs47xi/UVM12AI6aWIFpuN8lfpvJRRuZZGMrbyhBoSb7DdlVsqStCO5lh2peTRGyiDj
h8XuydxGgMi50dC8XFMlUuTIn2q9EvjNzY4KlgPcsTa2sW6Q4Z/JECutxLWsAJ8EPwznsEV25IQm
ydIQ9eYSa/iqxAjPLaee3/WTFBY3BAFXn5piTg+25OTXhNlCEFvggZa8QqaejTWBiH9SDgxhQWZ4
jQrv88SuXYbMJGL8F1fG26aCy/3BkbvmBBESn7AdWTYy0Az2vIbGJDFNvoJ6bbcF5knXaeGBOIG6
kDg6UsCNRhjxI8GmDhdltMNkrBcmska0S6XDCH7N8OHA2UEa+GzOZ2h5fkjVKD6tIQRVX6hCVxf9
/7FqYT+6CHONAEL41J93T05OA4OLHAUAYMg18oib/M31zTqlu9Zxc02cKBVWMsjFbHRx6rfE/+6K
G7+1VEKr2mrfXy6r5viGEaIQL5+uzOoELvqnJXzzTSav5zoDmMMxAfW+lPnQPQ3Ac6xBPYZakiPK
HSYlDMeQiOXycjTBbH0x/fkn9mF1rnAa43/Yaixuo3blH/7l32oN31xHcVGXn8mv+D1EgwmIS3JY
tOnhlFskt34ikznNknl7SEq7ANNtotU0RReqMOU2pYxfRJZsaiNZZLsgCIft9ghfgCYA2dub21vM
gfofMgqCY77YCmgxFX16Eq/3lXT9cEI5A/GkPYh2WH4qfhGUGnpbzH70vQ0HMDtegXqkmTT/1kgf
ceKxB0EfiUU5Gz3croce8J0TpESnHx9OuBGFnFxr0Zho/bMfhfo7QwP0bWvnVBuijeRcmFVBu1RH
4nVAs8Wo8jYwRkD93Xlwg7ZooYUOnMvGLxRNlTsz6r2z/TXuMhpufPIGdciPedFRnMgDAvQvV9hy
LH5iQK6VagpKWL635i5pjiXmvL++wlPhOLsm/IqcZJLZEP2aFnU92x+TnHF/iBZz3pfUku8v74kS
ZiFzBaHUOZc3ITincMHwjv7AuVJoKda+3jvvH34Do2zBlj4mA2NHmuJGsY3aarxsgyyUL3IwlsKi
kifwmTEKfdqv7NT03Ht1yzgCAfnKM+uRbA0LbEkZ4PlBI1CNHvdonxobaVSORkkTg9gMFwjE27Ud
jsIsF+pbtAgbIya3KPFHp7qE9764GGkVosuyT0eN+IEgfsJBu3JR2I9fAyGA/Qpf+zSPFdcC9zMM
juw6FX9kP9iliCs1g9ndLm8wM5Au2t+fBts1CBGvpRMO0X7H/uhiZBL4u3kSXkj6QxwdqEISkqep
vnQFNUZqkUronOpB2gVbCjFX+tlRhdqI6WEGp0IDOQPlxua1xTo/3wV5/osRC0accbPJhMhz8xyV
/C2w6h5VOmH+2UgWKcTyLlzf+LPYSBCto2SuBEYrdTcKcH4RFFzDHLfZEj90HsljG9pvxEz/YnH3
+zQsJAIN2pUdR0Tw7c6OvEMi/behVNpS7YAzAhm9uja/VZXc+bj3x1/oRuz0keY610+oANzQ/4JE
W35ws6/uTV+xEjQ0iBuObR0e5iEVNq1XKi+ZZ7yVaeL41j4lbOVK8pWurqQrAKcSqWQtIumtkWgZ
8HICYxr2vgW3hLUulfcnZif9sa6Tk4Gt0Lg6smbqa7onJO9OVwZSMIvgdpoRM84xHit1y/YRZNtZ
TbIFhQPx2zv7mixyRQzuro7iIWelvOywXhN+P36zIl2OoAaR7i6A/oX1J1wst8AJSFdee++NV6tO
PHiSRoxtcizaEzuzb9J13fyQtwg3xkGYkxGNotYiza2p/UtP8MAJEHuEsP22fCSokBI4PkILxJWW
vujhzrjdjaEpbWjIu7aljw5sGVVCt5MoYB0MB4IDOg/8jacAJvvvquDLvQXQKTtmaz824ca+VE1c
qYzOtD7uJNjFenZRbPCALFajK+SgmfPg/eJLYg+4+4UhRzMHjBUofQ+nbni3iO0Z16utN9cz/Mwk
+Ym5tpQIuLHflchuyB06arS/RwhsRbrjYt0MFrE4/eCb70E91i10ffbg4uzmaJSiHcdf1kNVcol7
kmbNvZFh6wzymcSHuBcNSRUeoWs+KAaImPz+ft5JQ1xx9QiMHG8WXadZirKzwDhoQiyzhU1VZj7u
GhMCc9w5e7WfA/fy4A+WkuVyFqrKXPNEuYtIMHArx5gDwYeBa0A3eD98qBeCJgALdwHaG5I3ZzVu
SSpCmjVsPGyqV2CRyBxpvqHiyzkO+tgnOPBtWqMISUYwWJF0KEXHTxzt1shNEcGlBTrhWh/kj7/f
wrGb4p/KRLZ3AFglPczlTV0Vh6LUVDMp5PwveGIT3bREtQxfntK01/IpqaR6rxVBsCvQ7UIJJ9eR
q/r4iBW5UxL2cfZrFT7TEzMN3VkO9jxlXW2x0e2JgdOfhXlUhbcABCdPHJausSBAulBSB5OhVa+1
cAV/6o9Q56qGsK3HPe6Ck1zJ20AIfrMBzZxDia99AQF/1zR3T5lpWla078K93IOgouOt5URXd9/f
+3sqohZCkFmKVS9IbGlJdzJq9F0mJ4mwxBevq8fO2Q7ydEEdms49Q6gOdERealW+XLGNaM5oP5fY
X0xcuZI9Ia60n+2irm8j2MxkAPfmXUaPTxWGKcgSC7OpEJF8OWLZC/F+KsruesN4+tj400xJfhZY
cWWtC1pNWaNsqE1BxZOojwzL+ub4eMbjuUUPC5oCfAMsc9AG1OfPSFrOHsxqPGIKV3ZEfv3PbCJ6
pFvlePk1Tf6YbXJ+mx3r0bMuQISSTVRrfjv/tkNOf9lofWXAsf9qAuH1CB6D8/+sP4qbaG2oBore
bBbwQyR1rXnzCHc88oJ6HQjIueCVSSQVYuk72JCADFYgavgla4yeFUbMg8uplibSfsZESJZH2MJb
P7uKJlsDhy0KU3VvnLI8c5FdT/NKvJhgCBDc5gMFDsV9O+7ev8I79jp5OD2YkbF7DQIJZWU3Adoa
ZVRPT4QffhAycXSzGpiF9JXt2oHhT8TQa4c3fjQfWdIpNHPiaAiuWVDuQn3S/zI0TUcC1bqbJ9Xp
YCVCezxpISbmVpk4giat+IIPPLJHicu9DdlKSI8txx6gY+6S7L+2Pdj0BvKH1hXfp9IPnbD3/Reg
1rugv0EeFpfmQsNt+F7a2qa0MicavujokeEbJB5YmUoT/i0xrXyARhwCsK/NbIX8HRCuGmjz8k9t
V/h4UKhoo+oLSW3IMdKLWS+lH2EFClzfeRWr/DszJwDunsUhPrOWFoOEb/IAUp9wPiIbA26CbI/I
3ZXwk0nBL8rpX2Gb8RzCn5dikv/bsc1N22nZTaZgEnfyv0pRUub68m/81c4t9DFaPE8es9uaIHf/
ySIR4M/rMKgf8CGoX5EAG0AjEwLWEJVq9y6AjKTK4bNE0zKP9GTqt39bcaiZ3JsVIjQKrWr1uLGo
2gLdHAmNbkku87TMVI34EhX9wnpJDuKydTaQcDRbSunLefDHUZCZdvd0lbMwGfquBStjm/c/DaCz
eyZ/HfeQYZfEce6y9UCQW+AfAkZ9Gdce2Uzz+dphYrqEGtCGqp3Xn5hGV60AYpDVvkBJjOFxNiAs
n0ZCesFwl+aa3OzTeR4Zk5tAk7sTUHDkMw635qfMooJS4TPywKctmKJbeMjcV3xzHkAwY75nIiNe
t+mTIlcOo0pVcKw66PBcZJJFwIFQV1yqOTEqEwQkaVXZ/3yUoLmPHWavq/oKheUNy2rRF5ehNEEV
N4siqVRXFFDmF76xTd/68kI2NV7q7P/iD6Tw0rZwQO7FZmSZvMAqFn4QUMzoqVPwNv/VlO19wQTs
T0tT8rnz+As/zpNPuxstHevaBSONUCdFfkR2IhutkAOPluigx53ccaSZch1k4TKX1aV0E8TEqX8V
O2xR8RzgwREcLOm0pL4VodD979wdF6kB4/bI3xd2FX0G1zRJ7D8jEkG6dSNZvhXvDtZ8gu6Kfc5x
waPj9S7N//lIDKzxdyETcQxX4TPxmd19Q0jVwHUxPrsozutdkiTP7qnApFyVNXRIa9ST5/52Vvqq
NlUTYjrcrHEubvHAFAjk1aCbn+iTPykXb7WdYxVypVQXYPurIN0iT6LuEWlfBrXDJaRoExuXuXOd
LHRCH7FS2nVxKu/3C7emZJPuoJiALFYqBQSkJ+X61RKOi/OPLbR4sC36sM10vJzw4RviceOWfGDV
GOBz+GZkxKTs3NdjTxGqHIMbxVJihOCI7jG6Lf7BzGY6QoypBrIYtzRSJge/yRK8wQQNpzfqWmNa
zsaQ6FwDk31mqR0puqXO2oMtRh1d1N60uPrOcyjjQJ4USU/Mzqk1ZguQ4hO0XjXhEP2n+GDDUPjh
oyh0hzm9ik/pjM5G3qrTts/G19UDj06OEklGhCVTO9gPOudPWp7V/jPUMsu4d0h3hx4HjpmhWMEC
mu5uuX0jqDwsZfUXdbwXsTwC1g0Rd9F1hzDMmMcvL8DOs1L5lk1+tzYwZ+Mbue19H7bHv3jU44uP
W/Xp5CRW9k0M9W4UDIGCYTflKnLerUZ8hRNm5U40EzpbIfdADH9A8fctlqWvei5GzQNZG5sYvZqD
oh87S8/LEDRpG1U4FqB3s9WTlt6RxIIE9ABSHw2yu0hASKWPYJq0OOQbB1hEqc2NgKY+RhVSongL
i3IfY+FiRAMKTgeAGFZ73C4VgXmeKYw3BkeTmiekJwfojW4IVMPIvh6i6Ss9bCcoWqG7sf+onQRj
162wGiaqyUtmkLKIY9YJkiXPspULyGWkAQwgFRzManGZ07yKOVLR053J+2epm9gDAXbX1T8wOjL9
IYbPbjAi5NEN/ov/nw0iw3eIcG0xiSm1k7bMmUborS0jayCCEGOoEcCAovOMsaaMcFjIZqU6pVjJ
V9a+JTZaH7HJjFsZv9BOhGecJ8cseaUzYqnO2FrIXtbpvLM+aXQ253lAJ2JTbzkx1CK6AqQJ/eTP
Z2NOVbsv8utA7za02TBboJiqTTqtLjNOeNzLuzOD7h4QD/ONqHw7MqpK2Uq/0KeHtRnOJ5QipLWV
03TUvCLkLPh9GSv6o90CDb22R7HI/slhAmgl43U4q9P8aeWsC9KatxOLAEXdQZHh4YBKzVXag3TA
EZqK7AFIyVgSvbv2AVasuhTdoOzSjLsdEjDzSU4yFrGn9ysHClbdPb1ascjWa8TK1VtTORXpBfEw
8LIYfULXcmK4ag/YpbeeY9sONTIk0flOgMu7UXPgNQr1Q52TYBlHiJOgpXdd2C3p9Pv4HNPSjXeC
T0vBO5w/OC3IlEMeplF0CtUSRzZu2yjEOfEsUesi8DiGWAhpVqyXRuFCcGc0chCxRoVjP8km592w
vPcPWKH/tt9BKBGC12f31jmYHyh+Cua4ZRe7np9u3nC8J/J/xCkgRC9ER2KfRAy78wXFlKfvZZEs
qUnSbRM0Vumto9D9jnGmTdwKM4P6L26LtOi2Tv6sqzyzWc+UBKYpBVBNiIzsbT2LKNPcwG9RYPpy
8gQlZajneLNGBCPWcuFSpSgFoZvpushjwYoTz66aHvNRMyFBCWnm1wakFeh99+e/eV9On6AIA4WX
k/np8IGNM3fPo6OVki08/mD0MLpo8fFG+8DqCvGhcm97rM+RMtzHiovR9jq2FZeEFqFzO1zelF6u
Tl759nymAqyrnczc0jH3eKERLco0cfIlIydf4ymLHN/uEl0W+TbjIhdnc7z4/IIwBJZVVsAAyxSD
a8hMUqjhGbIYenlC66/7FtG2Un0/J9Tp/0+FUYvdyx+n4sBFd/fmCiPzRRUo18zk/tE2kczUYcfB
uq69+0VtBPvo5IDuQEJJT++4I0KIZATzT9rfthAuS+43BZXrAVsPiTUR0pIQUZPhZnEr9A7iwhWu
cei6jQH1cY5PCS47KKKkLNlByiiCn06kbzGoEyBSCjZ4W1QqNEsC7b+eebmv8wfhZa+EyecpvxgV
WYc5ZGRagTW4GwSttkibw4gbTBBHQyHnoYAzV/h6Ic6Y4dzLp7NeIyOfcnTY1m4FhyvQvCYAtW/Y
TiG7UR1IpnvuNm8t+gT0qpDyUslwnO05LhenjhyNR7fApEHst20z06eegXpasdpHW8/hT/RgxxD1
4mVIqTxRhs5fZ4DGh9Gbq//JoaF60+pey7lZuLbbDq9CH9UuS6yRy3XyEbr7d9ZU3fDUDpF1+CWG
NIzUy57zB/FY8juZfCWYeCOCoosr+Ks2oc8EcaDHS+3bglP7mSLHXlEZ69KjpaBW5sDSMEydGaRJ
LuSkqAbgcttwWnK8N0YIvL2Id/gYjA6hvWF4W5Ra9KJ8YR1hY5Ie0cJzy8zwN09RggsW7ys6Kmo8
MkPIL37W5uf14uCf3UvdKTpxXzZQpm//SoKQsTf/LtCQ6Q3JDx/ScfYF9yahX96V+JC03XIxahgC
KBwp1NS6BArZoQYujmANHNWJ8YeCksTaNTYRjsN4kjO8vsvVfJlYVHL+ESnKLK0wjttmwaa7SRjX
Gp0WCp9NwX4OS2QrQ5WNNkStLJeXg1YE81PbiqqCXcr6PRP3KRWr7ixpMEZwimFAnVDctWMbCZOY
PK6HL6u/rlj/gTGtYQlfj+prL/PmwZGDUYeJEtVQi6bON6Imeb4ZyXXN3tLRKEQCnJNB8eCQcBDa
yfN0DRAeMMJqqVmJzlQHi5RrCM7z7Lc35LU2VUYicCBI+4O3PWl0wN5LJaOAcYXVZ7jUrPzqvZqe
l2+DWuisl/UcAAiJOONurHQCK8exZKyELI8IQooTSw0fm0jF9mJ+J93l/1CUE7igKrQA9SWUHMif
TP6Y6OvTs0hEJzV66cviK4gJ7ZZMnXM9q75SIvez506eRLi0eMya2S6EvWQ6bi5qkTXhipm82s8A
kH61HDlBKqV4uw2gSs3D91GJVQ5PTlbYoNACk0IeixGLZ1yoam6LpXVSS6ny/t5w5uJb9W8MlQ9/
qDII1od9p02bbBD878STy7cJLLc85D/xXwvqYpOPybPZSn3p880GypRxGJNznZ20EPEmMIiuZqP2
V3tEQCnK2AFCBdFL+7llfwhxTDRZRG/2oLec1CrmnLk7QnB9eKT00QsofP8fVSnjgQEqvSPQQFFl
IBgL1xG8u82dUZhpezJZDVSGnO/ExlGCnGmZFOBaiU9TDXrRv25G5O4IigPQ+FhwOLzbKcajHKHr
oymLtXyMx7czvnvNxhOWIXWYRC80vDB6fDuIAW2GUM88VnovL0dQcgBEmsYXJC4YEyEP83AoeTeu
bsD4TKkaM5qReu+/E5E0xtzMjuzi+aJ5cmGpjHiYvZIwqEfXEkEoPITtiZzEfWgLSXDZZ20oEa7X
/nf5W8aQTlEdiVBUly0mxFwENtIGAcYIcvasbdqiSCk3RR1nUeAZwlVYCGUiqJwDEw3x5x+JDo6m
4yNYcHsyBpjl+NXk4Sc+fkgy83iB2xvPFpFyqDA9u6PBSnHoKFU5PsIWBhfA6mS6jSiJpjK/bjdI
qneYRHhWqwM4ZLYa0sY4ijWf4FUJ9fhn8xL8AsMAqC9Htrnf01kElMvKpMvCOvO11MDhvNijO63I
G/BVUHVoRhcVcMUli/M91aZ5cHswBALsWfZYymo9CLdogF2omXjRKfcz2F9hSkEoANO7p1vqZ0Qo
6mh3OnJ736PtG9Iz7zxDe8GSi08G8Pw4SaRaRYb6XwpD6qxNe5zhA4tbQb7n1p2+G+4Rr9uGKYHF
23qUGgBv7gzAlVod//jVBDsDGxCHkiIlLwTCwCKfDLKEFawlEFmxbfPzIxCUJ3BJkBbj/MjDZ9fz
ytIQHOyTKXHIWVoNw/89D0q1e1fwvk8JouHpbx/WDOV9+kJiiJwb66Q6m7WddelUCp33oJ5qLtON
JlbAsuqjTSnqCxxYCOM0aB2VBxyk2OnRVnU7Y+7Ru17w9Jn4dsYs3ZHmQxdxPMJLEaiHVzrD/M9Z
ag1QidFNM/9DbdNcWbE/kvJoIWiQyLvLk7U8Ju69eV/6hydykXgI+gZXyeYYru7SUhbuWbi3hRRp
HJy5SQWaoC7Ljz5i/LsbSPGEQoHqHOXCl+GGIhS/aojFOQB4yWA6SLyH9N2pfc+d0I0DAlY6kqxA
jY2mqd+OimvaNLgmlPyaLCGgPr1Okg9InmDVbkep4QxL06gGfZ1/zSibgfBdTGjwyaQ6A9mczW0K
XcUezLPhl603YhDSNBuapnmgKOS9QQfpaxfYFfhwfGNB+adgmNo2Fx4FlWisch5oMSmQ8EK8b+ce
QvkHDGuTcobwzdmGnnJvrt0h6qxoO7WN3NPJD1n3xE0evyjDb7q9cqdhkUyIxb92yHuUe8Y+j3b5
WuVjwQhmSaQiTMTF0UZBln/FEqz2/WaRZaPahocSeAwldFCsTToojTpVna7JfLkg6EJVPn8P93Kx
RxK7QnICNDwbbB3aSr7yLnuh4u7UqDtdaNSToxlgkoy7cxO3l2vUoT0qxbohE9TC39OldUedupBZ
DzjhK9jsLasNr15VMYL2RU/cnFgYVPeIrVyPoXW2aU/F3EXruCVt6pJlN2hGu0OM4oTVlb2IZL/c
CW8jTQtnhmJHGKf3dMcm485KyvlHPvBYLAQ9CpJhOq5Tckk5scJsMAvTx1EUxrmgNmAI8APZooVl
g7Bc9nE6vTqFmZCeGKFptfYmMJUcNyGZ3x+hYFysoRcknreIBRA60J8sfyd0FoIengv6urrouDwQ
YTMy6s1H4gKj7JZ3orb9XDxrKQUudyeeXmKswe0Q/vumT6rYKRwJOJ/Zr89RTExnMCUJZGplYadG
UJ5jTC8ho4D/wTmpgsVE7DF13a7itxCzR9njzDYNMeZYGBr3v9qKzlfyCd2ZbLQrN8pc4blh2eir
gVcSniVY1m+HRGoehF0pvT/ICSKDsnx9xMJHD1ygMD1BaaEJVFpAg8EKTpacTqqlTZ9hnjr6rw+w
zOaQqkduedmZqMod9zw/EzdBYa8kX4a3aiOzLAubcoWAypAs+4lzhPZVfmkJ2mWLJu551DBWFmf0
oK3CAgXzUz/SAY+khGzV2v0xsWg+FgZBDl6a9flosYPm62fdCHARr+APoDZR73MvPvJT23uS7K2b
WykK6Gps0V+bqPSo2mGLyCmJQPxYulzxAsvLhPWF8qEYdGBj2HWD2Jp3xqm11Uid6crsf0bJ9ol8
v2RyFIPtMLiB8dM2CZoOJvq2nSVd6ZSn8oxO3C4SnHLNSyr4MEIGCvfktqtzH7w6/xcN4+ywJtrV
We91Mf8IBXigBR9sv9B3rDy4tJs5+dfH9I+XJX5yRhAjhWwN+OvSFD/f9vqQZ+TvvkqGUj9yq2wj
TkDrvuFtSuMETMZQjBupu04hL/A/Sn3nKCPVopqpnLsPB2CQAuFSv6fDTSVYv/AzdLxEXPxrT9x3
xHu0YOYWEYJl0ATV196GBRBbLQQoZ/OU3zUi/YzBVycd6c6zR/olW+t2ULu5T+z8fkAz8bflx9iF
Kihajtr132VkLH+9hBnd/ZHooiZBv8bUlQyBC4NyeoBS8CScVIm5a6NCB1hFSGASNp/Q7KxNbKkb
5GlXLU8sTVfl+pInIDoRAPCcO60x1AtIIipTx2CWr18a3KRvw8WXXw+lohMgGtpn8V6G3BkNh0qX
25fHlrV4LO0zxIA6YGT1e7D/fCY4P1KgPo3OkN0nQxBe26xH42djDO8Q36ilcXbcZ9JScGRlRSrq
6OPg1Hf4/2KZNgP4+JIiKtmtNfNn2YPrK7aASvhnDgi7kd6c9t7dE88A/dF7gBSwoUWHq186UyAr
IphlpX+a0rUlQPZYa49AYemnMn4CAtjnW2mZrGTudNQx64Mz37V+9OoEP5kF7DjYFlW3oIJ4oazW
8Avj7vPxEuldNj2V+97wKlsw7g//YNGwSupv2mVBz9vmo7m4emwwKb1wJzDP4eiCoXpaqHuYNNmj
CVQnHaOWVwdriI1ewObhncSYnANGYxFqy17Rh1Q2NLYhKsaNdtFoitmFEQlITg0/6+odtKCyD0lL
dC+U9wLLPaEltiTHx0bll/fgvJBlrwS5Uf/E+NgmcW3EpgdN2HKyaKpv2gs/06AqoiDPt2g9CHRy
h0oxe2VZY50NHTZMZjrauOBidKNilKRpOwq2PwaExXTquU+3+EBn3UFq3DI/b4nwygslx6Fwkgt5
1Vx+O7lAj4IcKieZcJzCxQJKc/23ccNFeICjcPSvGBzcmrTM/H2ss85NaxxRJZFvfvspLSCYTs/O
m7O80/WchWtmWbJfG/pYLjJQ56SU7L7Sk0O8nVUsyT3Cz5krAhAnhZ7kJRML+GjkSFKlNi6Dfvdu
gkSwgorfwHUMCWwRZKxdZEew+UvaiEhCS0wawwfudJj5eawAqz+H/VYVcZZ8QJ+Q4ud3kfRu7qGQ
BwJdnGd6k22mm4vVO/8ZapQDHlLfQAxIrnZDZZJvsCum+WOChGn9tkbX8Dmh0lc+2BmovhWOoJbB
JynIsiBjb1iS8DYl0S5MJ82zoD2isl4QUMVl3PswYa8QevyDJi5kT3IEy+Ts3KFOPnQU2P7JwPcV
vXBeRGfa6xJr+cvgToJS3lxSSAQoeq8yJyfIjR37cLxLcv+ZJqw/v/KaBWYIEfbTxisYfO3OAiyF
BYUFjPbAVhKF8QfJeDcjtsCx7EtDrU+rav+UCCsGWLkum1ra4OP2RUeJnBFA5TerEDltyTV+3nYF
eKklNLUfpaCi2wvhp5cAI6/efsRQD3xmQztWNN9k3uJA5UiqYXuMhhhdJt+QvTtsVIMRS50rlimt
6Q+wk+xqO9D//FhG2I2KgX7VAEW+e9UF5cjTQQG8E7xxkhfrKTyQapNuLewUKRtk7A6aZZKNubUs
aEXIzkgwWPeZsU0neYhnu2NmRFwiJS7zBvRD7GeoXA+J2x+w9JQpSc3LB0Vpew8DPf/QTbE8XCQ0
I/2uAoZj+Mg6rYuJxpNPTihntcNFEIhke5kuOwHLNeSbh3w+lbRd206Lk/gykUEpsANFIs7RIz8S
SYr0OhnJotwFICdUjeLwVnQqwxfYF3XvaZwl2E6C4xaYEFjk2cO8kfTWUiZVApmTzHmzn/ifAh3e
jQMwg0kWd7RTr6MZh4SR8hN6WF4lM0OJHNR2bo+xVlws9C9pYYlBMjzYAIHtkMoKF4P7wDxR1rPo
JRuDmSsBJwT6w+gy7esG5DrwaiskyZRqIT1pZ6BPVfKA9hkAWsjuQobfUbtETydux/UnkO1nWajs
/yv1zgrilfozMIiHmK8b2+8vEUQFlSY+DBakbSwCyQPRRv++Dd2Ldz8d+FzNncn8HxOYKOz2cnA+
HpH+rCBv5BDsw8PKwPyjflI9cx3BvswJLrQ7NnZCe5ycbuC+TEzMtxz6EEbXv1kyvAYBvRPdRmN7
MkfsaZWePjFi/7rDZsoAIlidMk7g1st0QSvPm53qZM7FxSsYpv51L28tDzIdC3DU25gLIag1cccl
/lRKIBYJtp+E0CcLIQcGS+qzUg6P2WydyF2WeL4ZjECKQ5qy2b95J0v32UOhZFZvGGxcGEh5jK5A
M68luGWiE4lKOjSbPGD+TogNP+N/wxPxDObwJPcyhtjzD3qdK9lAF9+EdxAhysF2tBKimiiaUBQm
jCz0EjRrOZ0Z7zB1v+SXXJmumKkg4cpIHIy8OXMLkQr5O60MAL0Ta/otNrsCxpuCwugiOxK32TBt
IstNZMpCsBNpsGC2MWiF2X1qaiqM7map7o5pA6tl6/10FzsYvNK0dSFLwXJmcrClQWzWO08aV5jK
S6zzXx7aTdIW2dIaJQoknKQp/dlTuK2Eq6IKnO4LFGDm/U48PWDsIIZIKs7FALgdbfECTGpofga+
NEE5hYf8WTNND8WcJ6QKs29JfV7Ph2U7C4InkD1d4VsvoMFjxd2BAIqA/llXNsFSJCgLiEhLwZt5
dqsZxqF0m941tvbdWY950NXD/I6RTH6ceOUEHgZCV4LNW93RxJ1GSgDAIjS+jNUYvm/ZYW/UxN2/
pzUzjcFSRHqOocv/+Ryz4xlkQer3x8/7i0R8txUrIU9e0HupE1JqvtkGWYH9RqM0SPOdro0Elxe3
hApSY6zbNvxf19duV7aMsinjHDukLjjCEQ6X56qy5r+Xxej6gvqcuV3MtGRO1JcUlX2FmaEnhJ/e
m/jezCZWDSupKErTiGrw/iDHz5bYpatALFNhwnJMtqRX1CEmufJjBKedGdwbDzIxWMJugwMwL5mF
XGVHOblMF6jUsqXu0cpg9eqWPpvSovSmOVSQZ0gEXxoLsnWaA+pVQhiOpnrynjFpP5uJXky2OEQ7
pvjUn9grF/hNqgwLulRdCYp/N5Ibs1vGOjAFMdlngEdO9jQc0CLUrtRhCVX1JD37JXAODyZBNI3Y
1yXw+f8bxMUtrEU2sM74hRkq4p7BKWlLpgPF2Bo/Olm03ty/MBkVtfreJUhFLOA6H6n1z6nNDGaw
pz0bsS9o9bJWRwdEja8Visp5vV6PONxHVUGjNG5+5lo1D1rjDyDYzUO3BDSTVmkga3nA9QzLkNi2
4WLzocqJSAii4V13Wb+pN/isBRe20S4FbBJo/ZmT5RYQkLWhRmAgbOAUE7eNJCoeBOpC1Nyp+uf2
mipilxsjGE+pKJmjlKk0GSTK4QGHck6ZzcbPGD3LP9s3kUA+ivk7+xBPIeo8iFK7B00P2kZInBaZ
lRSYtj6SnFbGOUFzU92B+RbyWu9n9Z2sNvlVfhYqfRy8ErFEndZsXbuFO1s42iwdV/ckvtsyVYm8
51kSLWZEipp+x+qd8Mi+fLYO1ZNnbRQRu+QNnP7lxhY4M+qJ1DZMCtPurqdpLWZj/OtxGQ6om8E8
fDSFn38+xNr5NUZhTT5pmz5RyDTsoRxIjZPU/5SAhsvQhandOheEclVuCBmuEeb9oJ8H50DpqucX
wqLDk/1YiDnYHiow5jJ9mEwtWy1UKOV3/dwiiSiJCx0713pkJepcVT/O5KP6aIAKDvd0WnEp0Nj7
iyfM2VQaE6jWXu/83JAH8evC0jS7AvFapPgnKP/Sm+3O4ptFqv/iECb9e08KWbQOtT/br9rdBtLg
ngndMYZ3jQiiIdAeu4VjC7NSvA0Djm08JScT4RER0ea6Fxb96fFLmjo2AlATj7ee6xwo1KL4pWun
X+srSxSIGuf7JCcFwqIn2bLCLuOSRzUCXCHWdJA+i+Qz1BM8K2z/xcSmq/1+39R8lE3uJBwMIT/5
QrcwuYmn5LwwEYEZ/y81Iv8qk/cWdyNrQpbPp5/5eOkLmDNZm9ryCKaDKDcoAHLxhYiRzo4bLodg
RJfp0RPF8aGfMi/us5dTPMwJJ6tCFkXg97Pesrb6xESqQ3hC4T+c4AfK5avAb8Fb1oHrHXt6GPqF
oy7xF6i7W3KBwXFbKdq/+EOZkV0kXoUqIECaEZZ9TR6K4Od2hS56uKzmPLopRYdHiC+t/l3hqklX
0SSFe2ANqlA+qmRqVMlgZFBCkPosZQIaSt1otkd9c3LqFTBFtzSWUBiVoBbUZRDx6OiwCZf3L/em
IeM2TjKpC4KEZ/jSJWR4gtJKTj4qwPww3K2znNjIN69Q6idT8OIzLDI/IdKhGq1j9IgV3xfKXHBq
Lhdb+PRz/1S4E0a1LFS8nIuuUAslhGzmsjogSja9yhVjyTwme8WAgPYztw8KjJsyoVoGUr6Rneo5
+7a3KipHnqZ12sdUqgV9ttD4T8IEP0eCGcebESvLLyVwkgtOzPlpkMgtiSH74keOrpiwxn673fZ/
cQs9Weo6aMC3sSdz66/BSWO2jnJ7fYMr+WO1r1v3tHUyQ44Wp/0VMTv/AFfZrgKCnmERd9ZHiEBh
ElUkTMC12t2blm4TzK+FZd0U0TlKJphpfw2nP8fF9SBciPou6PLBGKr6iis6pvIy2t5yOTxHCcP7
qEF1/1Gi1L7Sl1JUiR7Ay/Jnknx8qKePEZ4suep+DIfVVFPsHpbJtgEzEXlltnNTAW85MQJ326Zh
k0o0l+y6IdyajR93yhro99czwkCaZvZBBSHerV7c6d0+9rk7fOmGvS+0G9u1bWV5fEsNQJyhmd7u
bbNb9K2C//fylVmvXdc883M/vwqKxSNPwBcDSVWjdUsV+34mgzxceF/hHxx7w01J6wqKivNq3jwI
tjYeWro7lL4DO7JD9DecjxPJArao1WWTD7ErTAWKAeYGvLcQGlvgf5K+0b8yO7pJWMs4+Q1J59Vq
PdrF1vKbHLtjDmgexdCH4e97LgWJPuZbXGPunJDP8+5fkXgjvTjNBTfw5r1/8HuftYysHhYPaekf
rPKWRhu2XOi6Uqg4OyJaCgPkkEdme9GAEets8peLDWmPD/mWiTFrs41HsGoT3vEk4hteLRswW5Ei
YwgXrwAiV3L6+z5K0oCazcTuQ6EBNFovUHHHAeeymd1KQnUzlXDb9mUPWeI+7nA0mC12RzZmZaLw
xv2FkIVLRzDbgapP4VHUwd44NfZCs4OKe+h9dpseT0l4RnyIz4CELWyexHGinqSnSGyaRVa1N32x
4n7W2e2RW/5YzmTHD6NO8FW8SDcvluEIyCHFLgy5zP0tTAGn9gHw+QaEJD2gPIQL055kymFziive
Yu8cJ99Cu3HB9z/Bny2i5ewuxrN+3ks6F/vQ2bnK8edkN/FPUttnzGsCDTh9iBtaCDjOAnwrlD2r
kILwFWgXNtHzjBI/GCdQffhRIS2rxr8+S4osUacYrQEq9hslU52veO6h/DU87sOeOG6q9L6EO3PB
oE8w40Z+fGjf/QRPFNmEB2ep3C6TZCu0kdHLInsgzK6mDIXOOTqtwVX0kL6xCvZnlCBLORieRhq0
l/0rkRKGEf+84pULVHML4sfvjBUoYiVIkRxnjBsF+kLT6ojqZbHXWa1JuLNnrrvtmGlflNGtU4o8
G6Nfdd3sQMt86HtCD4XNagp8g3+a/SxMZ32lBbbS/gAkzmuggazZRjVcmCsAUJkwMQH4SwTdFU6X
zQAblRnSZ+Q5zgut0ypPle45PAKBTxaySDtu3s/oQ0Mqhq7PFtp0hD3NSZP8zvVsVdpfF4NMoE/k
hb0WNvnT/d8rpo7T1sLCIPtM3p4qzjhEibrEsuHCnWd9NYbJ0YtvQQdm2x54LbryWXDqjhLu1Hoa
n5wDyNy9Qs3zDSGwJWG7bg4XdTyokwHBcuBCz8/ZJ5ue2Rs4eLHiJqqsmwn4Xz01qUlTEZmqQWVg
CqS4r9d1IMkxZ9BAuhNsFlPldbtxLOVw2PxPguwl3LVUSC3YuUz7xaH++RYjJnMkt/lIHp6ra4Bn
y73moT0SW/RSIHC/isXKWz+xubkDRwFaEbS2BzJQ0bAblirqQ8qhuM8EPIPxcv5S4Sp20cVs/8IQ
e7/VUFJ6LIcU5ucFomqz6fhKg8aOdQ5OAGKS0sEYu2grSmb8ZO+dc4I6Y43I8i1YTJoOmwmnvDEV
va12ntKJDgGQ4cnUafWx2Jy4S+6wVIYFl2s4gvUL6JxMy5i76fzjU0w0MgWEk6gX2Cb7GUhuSpYa
IQdCU4ImxbBdhk3UhMdPP/x784C7LWNzFHVQUDeOe6QDWlccOTjZa2NoVvaSlPP13JKtALRgzomC
LU2ssss8BfBLEhWiEvMzgvtnWVzfF/IaDsmDcumt5qUn6ByZpO3fY5OVe5dy8En72xEVKE1QaXGo
spe0JBFIzjXDkjB+MrbaSg1R+3/AKn2O+q9NWriQhDxWrYaikJyl15w7D50he7XvbiLXTR2mj+6R
lHnb+ncS7y5atNGuLOkNMxzChQ0DRmOlBwyur97aBv/cwl+1kNPl6Ax9M3r4fYF781NVlQmE9AUg
OsIKXNUfv0iNj8stIA4odNSTDtna06HTV7pYBhfcQQmEqgs/p8iFVwgJnEw70haCOD3T/Fq4MN/t
ZWhCDS5ngmWVuXUZcF4wDBFoDeOHzyRuZlGkcU1XjkU8pXW57MNfJgmRohPpIO92r0TWWmSACZN8
stFzp2lxJpG1GXfommtBVqI/dQp+zuDRDhbzlRCJ7GuCSin9HKrHjttoZ5DNqQNpz4Asuom7sw2g
wsyxrSWYvX/zvJivRONLGJUwOKy9bWD8/cykxhtYLXjBWNYyJX2w+iEv6BSqnlcX2NJ2ALzrIosq
v2n4CemKHvN/uGpQ2apBx0eGdmrNbJ/z0stYNiFHZhoI3BwnRZZay+JnBMdFfeyR+mu7QCyWqpll
SEeV7Iy7NX82qB2/ULnTCkpTPBuBYgUZt8c/R002j662zFdjAiOCsJbJWmbGU8SIkoSYecppgxb7
lzCHVzxXh7L07r/u+VrAE0AKLZrv/hxZMQRRx/PB8Ump+sPj3pOWu8H6gI4QzehqukIRJC8oi01v
CHOHXkd0eVUtbPbCFewrUZEIzAtg4eP8toI+y4Hi0Eceoy5yp02GcZ1dli6i/E+kAo2JyiLD2LoZ
UxHfTqRv39tDAV4IJFt8O77AmYZ/TWq06qCEDpzeJLPGEhCiUCYZM8pyefWryqnVhQxy1Sre8gwy
raA49h5p83iA3Ot7lYPKa6vOAJJAlWDSRtJACmwfSshr52NIrypNs3DY/ZCixjPiIFe3jWi8KyAJ
BwxeEH4/ImDWJNI0Y1fsQs5IvJ/LT49Iu6I/j2PbymSrh331xYz5MF8I+uPiH+q2EqvFBlVUwp34
BsqNONtql1el38ynIgElziTCSiW0z8qOqBPvIFZJcTvMxfgISjtYK5LhREziV9jH+lwbZaZQxsl9
u+xezYpWqCSqWnheNCLzwJzJmT4/OafpNJnHaRlCPgNw28aLKmfwy7wjDnQACHOzcFxTQoEeCq3+
JYp5duAo9uuja02ZEvCT2q0hA/3nfQtcCA+KLEvkEMFNTZ+N/heDpLyaRm/SRR6qxSIrmSX3qQGi
wvYTikbc4fhmDd3CA4yVitS5iFerEKidE0mQoWF6l1+feYCaWeLYK3cd22EYMQ3RDRnh2t+kj+PW
BAw57ysUL6Op5VzKq+rlh6mSRGHmJsZt/20tC/jRW0muWZ+8kN8DWtNKHqGG+rfLRMY+EIoyRBq6
LOAbaeOB53bg7u5/xgNKz5FwqqogzjESt3j4MVatnd+WsrcXJTmlRo51WvIqTvQ4b3qb5joH38yO
Vw9MqRLX8ji/cWVz2UQ7wXG5qVuwtJRp4D3uQ5snBXXMlv1Bv/hT7FWx/ZIUAp/e9GwBZJOup/lF
6FqARnXpGRan+fRTaIQnyklEWLX53NRe0yjIXZ3lBTUMvMul5i3eeuYAf5GV4jXrj2doCyAfrIde
xvaVagoG/VLRXMaA7WPdSWmoOF0+w1dLDVLcgW6xxUSrBUTouOc9ASCpAk3P8qFnR3l39SMxDEd0
AW/xu6asIvvniGn3vsqWFSVHlMZjWobAuNvEnIeMBBf/DOOpPf+CNE0cG0j79TkOVZeElK9lNTNR
B+pwOaVGEuckDISCKGk9Z/HR7/RTetMmIoT7sGf4o7uMgrUA0aOm3uD6v8vEWRlOOBUr6PZ9syQR
6mq4xzAkpK3+Gm56LNSFNO46uRMTlWAZ48ihq9NJjLtd17wsYjJ4xhmaoDcf7WWJb7c0iMXDAy6z
d+K99D2EEY56lvliQ9/YuFNQ5Zd6LUCpodRg/9iIcxfunEkIBojAmA1uN+vs9shpUjWX3vWalacq
AywR5yy3eZFPH8jpBJrledC8ec8q6HilY3+LFggjcSrEjc+jSNVVUySvfsBj00jEHXQbAUSlbyA6
OPhFoQUDn6/UAlvxgTsOhhkYjMes1WujrBmjoUle8H5755YhKSOzAd7AOysYeTDYo5Ki+lR2TsCT
0xYujiVR9tfseeZnyvJEAsQieYR9x3WzB8+0ObhKtqgXQSESeWCYZN3nry3yQrREkuAZgP62KEEr
YlCQ8nJeBatswqBDnTxv0U0086P10BswdWTGkMzsv3DT8gthxSwH7XlFbR3ykSdIjvTZ7vpgsV+z
blaFyfeoVgdxT9IA4tqcytm9ha0qRNjwwk65+I+E+rmbJl4deT/WvZD1ug6hu/lpekqxl9afCgjJ
lV/9owSKjlcfqzaV837G+PMw9T7bHuthpbxmHX9G7lypVRLdo9rA79zwEEUa6pnPMtpnwLIF/OGp
kMoo4a5w6NY6XiNlS47YMTevhFVuRuulgA8AQUm7Q63k6JvuncZFl9iX2tGp68iX1zD4kKydzB6R
YoQHFbE0iCCA3ioa45Jgfon0ZDrAxItelImF2hewZF9CkEB6SiWMTsxIVdxhUwPQvHAl80r2H5Ot
AtXqvdlgK/7PFw6SuuUmWUCdKSQog4p5xR/FcGEETyE7cG9WycAXj0dnpZ0KlInCrindrO4u8as8
czrFklKg1Lr0vMube2GbjFw1vvYWsMINULZL7yK2TywtbxCM4z1dQHV6hiBhmKmFiuZfhW6rYZXm
f//iS24OIalU1Q9q5MCtaDmtvZHBASEK2gWiawmqY4SjN9Xwbo/vFNb57iQVxcsKvgJ/jne/PwGu
PybB0Xsoy5vaJORTlUUiI4odizHa6YEx4AoHAoNod9OP1Y+PA9gGI96bR6ioUdhels8RnnIEA27h
PRBA7vZ3UTCmGvQTC9uWj2XziVYv7O1MkcPaLAxQh0/6ew3HGblp7FSrXpjRyxAMnhTj/DD2sPnL
tRrZo94N9NuxWekfETDwXh8f7m4hoCso3/rc+wyvAqRqqMqo8hIjruPnFancSPwRPuzxUUya6FxY
U429/lKYq+a7u+XmMarBZdog0P10NdpskkAPsIIduf1VL6yuYKz6os9QAmZ8+fGSirc5QLNIDnsH
kd/1BV0XwJlcQbgR3P26bNlAgWf+KkfDWYl5AQLMhUHKMmvdfIs6kCpJ9u1ihGgFvTRu3v9N3fRt
otqe87IyHj9PFGoy/p0VwAZnyN3xxtnKec6SNZZrHKn48Mfjs49VOf3Jjy/HUK4FOYB5rHULmhKr
DngSN0ofqaswemo6jLK5BVZFf6pfDSm4UmP5lpwbfXq2OkRIKgXrWNR9zrNaEQfiOLU5oREtW7uI
rTgrxzcmj+z1LqcMUygG20kuEivt5IB8YzgASS3Pjbvb5MpChJIqYRBaFGf7lv3NxVzPp4eH86wk
ReJLAmQg36kDfLhLzZC1ZtZf7yOxzgjJM9mZEHAm3cNbx4pZ1ap0mF2UPXIqX7+MVdULibjP2AYC
ZxEIhL8xUdthaWbKi0wnDTZdzFLMiHG+vsUvzeCYWgUv1dr1Z/DYJMgIdvTRpCgBL1kAaTRi/Vor
DqLOOwo7sWjVRnp4YtYKq7ngg/4bpERYGwPIXi9E2UMQTwG8aIKixeODQza85P7yrQR00Tnws8d1
V6bscSAH0tP6eEZhg6URqO62scGFOrR1tZJ6smG9t8cmPWbLXQ8lKF7KO3sCFJdNQBY3qPbyeb1r
vtO+3iiUhOVqtYo0dcQKNn90iktWFR9c6S4mdY8bTI8bgYihlQz6ssZGRkTTe1b4RT2rlyeHkAjN
I2NS8NcBCD1s7qwQzaV51SKgOCyf82nkvwNo/qUpiY8sbT/VqpxOfbMoPuvd3CdZbsUHZt+B3juE
zvQ38HeTYTT0qOX7TiBO3tPCtygjPH0aMAIDza/7CLsgob5v9CGsjNPbrHSS7OQtbQhREkRUKgNy
XQvXmJsLf1B5DH2zhmZDKoKupG/zu+Vj2/FRO4ihbQMPHffQuAzEPdfFCDJBF73YlOFD8UV7FLhv
A5n/odNX2IpQj+Se8dgWLnqMibNo6QQqTYGsyPPRggqh++exEsLgiAfbH7nzw3hl0GmFedWbO+YG
WWXWsyPMNJ/D9k43w80RDlScCs/xIXzlCA95Sz3m7rHZGVKimdfCvoH/2m/J22f9D9Iy6sxDowlB
b724ThSiQvrXH8OrMFVxG31n/xDWo3DQYcNqbF7FqibZIGkmIjy0TzjDSrhWPmCekNIBp08HhbSg
/2xaRnMTSP1w3SNkpSfN8/HHNhg9W1/9R29Hkk5IwJ2L6MWVfCAi96cq90FfSw9PH8PoaOziWitF
PseXBrWDhB/H08DKNioh0TtgTQQG5hmI9ETqr+AS50wHVEgXfSVeCPwKnnxSHAqDKKJXk6JunsU0
NrVSxZkKBDhQsOz+gwsEFfah2FFGeT5O1grbsGWGPA1fCMNKLMz9KwUaCfgUMs0TwOWEBeVHuozp
0HXTEvyGEsSMpLFjVkt5E9OSY2/YPkWCnC79ex4+qjUIxOenY7qgLOz8FWJ6sjEBirh7DZ9qAGFZ
66bMdsfwD69QwW0eRngeImz4Fvtm/ezrcFW1rRhQUbEDmV8BYnXGnjNLErN615xNMfoaVW/BI2X2
NCMB4o/0XDoLk31JSHmOasGD9FYgQRigBUuW0LsiHMPgHoHSH/rssAC02BYMektsCBL7T/0KfDyB
3Pya1xee2TRkxp1LkEcszqFCrdhz0bV6J8g6Z2RbbhTzcUIKCkpk3HtS4oVlZZW+14JpuQ0e0QPB
I08nGL5C7I4nM/wFRx5tJWF6DlKF4L1DHOqK/8bKOX44c3kEuN7t9g7Qnqo/HcKEBtOSuK4qR9Az
BoW5hJcb2YE6eixWmGeQNMOsYUvNbqY4y4pEfwXp6740lUPq33JIipUmp2M1AkoeN4LSOjzGAJjo
+R3ikrRFD9h/8jZdCIORTnNppJfA4B6lCo8SpQVO/K1cRWWEIPnZOGo5+58rCPSQ63KbnBM20wOs
k1CZPCqplmjtBZ6laYIjBInD9Sq/h1Pw5z0bJIAevPW5Px4815lz/NfvbRe9ZGO/xYnPX8AZjoz+
hM+9UBsRLCpd6C/PC6ddjnsk+upvq0MP2yq+sCKOSALrTiM81OhHO+oAdaZ/bigXOaEkV1wW65dj
R0IVhieaWnyatL8/5fdVLnCVDRyihHuGS9nMF5at6LY/CxkKZvnYEokHLe/FuNa1/dftWGAn0UF+
23e5wdbv+RSoQsBr5fuOAmjtSjXKezHj2yulq0uQLOuImeABj5Dd1MtIbjfc5aPOVosRciMwnVF9
GTL/tCeu52A2uTPydl1b6Jw2ar2nFYaWzvZUW9WlSN1x1g6pa9bRF4W4UccpYMaWmtcKfaPzbWWD
aP/sIYcJsme0vF1XX0gK5QNBo+GOFRg5NRXuZYQPA6qfbvu+L6G+7+1b4KfLQXI4v3Qk3bGel5C8
rse2EU5sT2CsOpoXylAUaoKW/VquuWunmYUVnSuFy7WGv7NFKCfix526A9W0aAPrCAZzhzWd8jeh
E2rKdP1DLSF2/5BAkHzxrDTHdKJT6g8izYB0DFJOlQF5OFF9RRwqr6HgYw1VipzMvd7e2eHPNsYy
jgUM6FrSrk5/50fAiJJtdohIT5ftXAPvNmnIA6WFWkm/TZhCwrJuL3pNuceLxmCphIFCeXfzCBGt
FFEYddSCC3F0+GicHjejEtoWKrEMEge61a7eAyy1udmlPaeaXsL1IgIC3E0oyU/ni4xwc5d5e6yz
1Jz0Wo8ceuF9vUh96fnCeSbfSpmGutMSIIt3SkgS6Jn7E8blkVgG4Vq9NROIpMver5u6uLOftJO6
IFoBGkMWoRTjZMkBUJf8i+xANPtYau7oaQ88m1NJ2XGsq7yP7fUlhG0TmqD+/P1gK4lTyLQeJH/x
4izYEUcTULC1gXODH4cvqh+rsEKLoCLV4yOGqYFzAPpzPyJ6wiOAMy5JVe/xchODG3N1cZVXVAcx
co0ZlSsGHdV8ptMpMhqGU8IIq049uZUGoM09YI+cqdvvTugK4mpSCWg4T7YxngmVr/z81Kd6gaMB
dI02O+mx9tG3nQpvv01q2thzVB5KtOukZ3Lzlm3aBzurmNDIk/7/MP/nZ/bc9lHLqCHtlumXoyPS
Lttu9aad+P16EFahsPs9hHOLZqjk6OlEIuXMtljZ+WeOxVTLSkISGsymjzrkRm5kx13huhPJn2Em
+pHhfli6DDHzzc9sX/6n9l/SzII61N06rkV81Z7wiWoCWsNGrV4S7clV+T6iP4snJB3G6vCumgRL
UQLq32/MGC+quuJ+gvLeSwXwRNk9Q6M1vvVj+OYUB0Z22KIhPigRH2Ijy3a53jcmXw03YUwppXIK
843zIR9nRXaJM0GbTola7mZ0yj17QvttSDEX2eb1UzHy6la63Y4M0r8xIE69WSU1692gfP7IfCfO
kfyBGSzJ16EetRvFdFzXJUPrR0MYZZ23plTDkHzzJZfKpRHrK1uX6h8yIcJyTvUkMytgH1yYlHB9
7IhNrYd4LI/9lv6riolj4TY3lkWSsH6TrdsS9CNoaJbSAXmIAVW9N4T070nHrz2YsE4gE+HBhnQ7
99knMJjqutUDLGG+8gi1g4BAkyAKpxW+0vX/sTuLbGINcPZp8zyVxLKyWD/3RZiAavMUIDp2gt/p
4fRV+b857TqNa9H7vxoeA4OT4G4pOHwDYUvepeR+EUgiUn8ASoVn1zU4fC3Qpwfs99NU9ta5C8fx
uWAijbidGOSW8Ws/RvMG881e8rffAtjr8Cul8dgAFkvOjUmNgJDc2YrDvGdp6F0Kko5ECHlbDEMN
WDXmqnCruVsdZKeI6+ADdXMvdNUoWQhJ8Zt3OIItEslWXTf5tf8JSdTOVIpSkT2iMhrPRgwjNfY5
/ZqDg3OyxVJs90Lyaih/2YVGs/LW4XqpTKIx1blXuWUa/KNENUZv/V0meEVXXhkntcOnmg4MSuPF
BdORIsQcyazotV+MtRi936NVNrMwwP796udWeo1JdCLzb776FnHK+EtjHyE9ElyGsBL39KJQfh7w
m4opF3S9+GOA+fY22XHNFxfE0x+lVIY68XM0naiIxlqQjfxFAtjyINZNCDFmAVUxRHpaxrEdSLtx
WUYLCTxUK72/pUpebe+nbXCYora6/Sye+GN4NLpZ7fqsfD1poseGOB4UUZBWMTnNjy6i1yZ5+sY/
uavf9KLdYCUAYVGspvZF4UbIXliGSsIMhlExfRTQ5FoaeIhdiGcgcxo5MrlmQzx+ENzltTzudqdw
byoYlwecTR6Evp7OHpjNac7OU9do4iJrQwy15ww7T5Rii+3yHu4cHsbhWPr2Dauh2FHb2JEonDCF
yK/dAjO2ELsFasbS5XXEhMtdmN5GUa+wYVD2hgam1CpqdJQ0l2duV4CAbytCf0ZyMUeLjN1BfTzf
mpFyHWB2pyWdgLX/t/wSV2ZnXw6I5iJQj1ky+Lg26vCS5fmrdL4yckF8ot14EW5zb1q+8kCmiBMK
SEiDhn0rzXdKEtwPbARez1ADj2K1CzYB+N58u1d+AdY2onMBAgue3f09tj3+ZMqjll0vloKkWJ8F
W9b2yNPInVwxPVgFzP6jyJuD6JndelSx1JhIUI16C9DmbdJ1mwt0OxNolKYlSgX0XSVAcs1WXpY4
14ujy6OQ7D5/3Ob8cZ6kCuLH+R3qCTNu6riKAkCMuobxrPxnLbzeFOAWwtQ+Cguw4UGCiUq4KhyX
bY43M00e9SNQ0Rb90XoZupQKKhmi94zObjCb9f3JX6PQA520Q9xTyySkIEdFmUDXYoUabQuTvkMy
z7ZUoe8RatHiyAfX1tYawfbThynPDDVicFz5kCMrDQuHPhZ10PnCogZiz9a2Yj0v1NSN24Xaf2In
pJeu+sUaNvditZZMvlM7uLlWfTF1eRrtoVM197uFt7wO6nfm6y2/uTsWewdPpTJIF1gKFWGPm33k
z1Nl14XjAaiuiC60eWQLX3DO3fMuIh8lOc73b45T72M/jeH/GUok+q18B2iY0m8k6BYmxUjvViCK
Vw7vAk/ONXYz9Lz+GrPJKJmrSzaf+1DH5d5HAJCQHLs6udTmmJAx0+gvbybOtu7tgPA9zMJ2lXbk
BIgkH/McjdXvsUi9DmkBFZGC+RpG8E3jKU9k65Dy4BTEcM5dzDp4MKcnwhOr0rKII7L/PswwHEyW
DdKJJbpfiCoBGoadFHV6Sz3v77mdeLRT2SsHUbsT+ohomAXHDYzE+Qqj2l75Uh+XD1cvCHbYdgSh
1PYCi5IA1bENTUXfrD+QckrdsO3euCgqzy3fBabIPj/pfDBwhtsn1nIY7uT9CgTX3oQehmJC4zDc
OGUs1myNuaUBdx4hKFh87sqSv++S/UbTj0lF5k1vi9lFnRzgXWiDvvjuHcOHbKxCGGItjeqvg6K7
5JU3d3RRBHUmPXyeTaayg3aSK6LZPQJlFqBnii1E1AiDyXXyG4FRubpuQd96WBAj8QIIgXUQTKrR
mSqfZJ57AQJb2VsIP+04gSlNWMLic+sWws6Lt4S30DpNQjcc1jQUxl/7e7kX8ECAD2Axh/JD105K
kc6Q4GmpIKItE/bs6SyN8ZQMt55Kiz7hOnQ5TnPTVwwzp7EeNAfyg4ecA0jQ/WJR1GetVh02nsyo
/obhJ+AgcUlI8zopKvmEOXYY9YhB58KzNfdGlSkKwom923+tUa7Tr7bmN6EOS1kif8XK5c7VQM/j
lJmltcr/zTNXdZdGIJPMqGgctznb/yqeomzLc9y2MpcjvU7XB0jw5jMZG/HirKKhl4TZ9WfDXtaa
8YetAKQ+612I+NHSUCMIK43jYj9L0JVvRLl6wMcHRFszQsnYXyLCdJHGFXezuSpJgFZ4BvsNRAaO
k2OW89xzWTYKsM4LKYiaZltBtLigVux+9me4L1oIhHQvVqm5Rp/ZeJNyVDS9l7O89ktZjVQA2ev9
U/+ce0ZTS/L8C+JupEhl1J1ccbKe3IVvvFm/XftXfGNCHXUwqHAdTXXaqiSgbtQHZc/ww6dXvuEt
CM2vgKF5Zfjt3TfDqOcGWyUA6KLagdUPv2I5y38cGpY4ZJ1Cg6rAy3W0gBX1Dt4uNrBSZ9S7saMn
UJbQ5miBhhFxCJyCwcp3/cOn0FdXjY37Eri60q5XWjePp8plDxxHrJ0ZN/1BVENGbysOZupFlfHr
dHllpOECM5ywBeaf63nAxU/Pa4RT9HZSdZdIJADTJAQcwMqerewi7j6bildzZQamB8gLGhIl7vvz
AAKT104lvrtv9H3c4ttgJ27m0h3AVDPBoyImpLAZ9yZ0n+m46yUw3HRPShcf92h5MaGDY7VCk3no
kTrJmP7FzYz9Anbebd2spoZHrPY6RxjJn/AesyrxOg9C4mEfZlvLfAe2OdU4s1hIRyNPUcXuAYvR
374V97bf4oT339tc1tiOqtgsC2eF0SFeQYG/+69PM4dsW3/QgHSKcNUx8In7uoSLV6y4KBmxNr6b
6/2RvMTWwTkyWPRO0+KwpF/p5HyfW7z0fKJKnrsRv+3/tewI7X0SsXAik7phaQ/nSWUVa2+yuEFd
XRSbU+wRrkxbAVMXJ1OfhEiQqR62sXApaHouYpjQBnSr0Sj9tWwtZwrYbQqh47nu0W5ccYXEGITF
X89kEVAWEmmFT3yHfhe4SOnO4S376W/G5UR9Xo2/rMzTjDva36zjRZx01E00MuMRHPy0s5u4k/YZ
eNlpGu2LCN8OeNvtfaCcKmNvvchgtTCaRFPfERfISk47KnDNxIoHqEKa7cxOx4SW3IpVzVFPK75Q
4O+XPBOYNSyI1LkI7J4NqB1KUCeflvf3NsakLWJxKA/LHjwmG1fqIDIAkZ9bHU6BwfNIklHJCbZU
q0n8krWU2L35MrKhgcXeew5X+K4ETovCuqhOAj2wiGyZ/EGtUu3OLGyUTa2uToiRmriIv7l9qsw2
5rjBkjgqx/B3NRiugLE6xVZ4vzNyemYWusWIuQsLLy0aEH9ApXAgsAjuLKQepuddnVunT0kG51W5
SkQNqiyHrNqHgiZvPNuH1BhF8AIJoKRu6hT+B1y9icMBA/sOUwDJjBR7qJYw1EqZUXpLuDaizLCr
0FabSjv9r6jppkUEXp3YE8EQ+byy6aH2p5TCPqJyn6D2tuhAmuXWVwRaJk+Mi0Qtk3SDQBGSfQg/
Hurl5P56VyaAZ8/YmkRbb2HL2UKcrNTk86SaEdBhbo6rhoaHvPMK5jRO1IK6nojrHGIjbbpaP+zA
2gWlwnKrR3wVP1gddbBP/xYF+UVxl5UgkZZ0uk09zf8JyWu5ySR7cjU9hSaJdYpfrqHDjG3VJbsp
v17ArEZSggzpLA5kajS/+CqrYXSOgeU19KF0DSERbcTxylrl7rroXkdJYSQPoa8GPUdYzDgWvIM7
s2nZDMciytcBKjslSUpVRgAHcpIBeACEAVfIUn5xCOSqLg1x6lYMiK/s4XGVCyPeBcFG0+3oIIB6
cYMDcLVrfU180G01DUiHv4EoFXFE1tgt8WwinBoIjL1+1UkGCZTpmd2TMQBZCtBtsLuIO2yokL00
2Th9xE1qKvRhHcLegTnyH9aTrlfqNfy6m0T/+z3yQwRz1/ysWp7CAwI4VujWBqqgaLsBpbsvOhSm
WTk7QbrYh5L6oT3L6QeVShCwK7qAWXPI44XauiG2vcx2RarsLs7vRFb0klVXS/t6182QHdvN4OH6
v4HpS0lKZDpCcBAKvwKOZ8H3s5RK5AEJIruK5LOxFPfsLjt6QSsRrhUr82bCzhTbpgn3Wj44NRUC
BuKZ5ej0vxvNPpzug8pBlxr1t7W1MTxvFPMF/yPZuEQl/8fnZf4WebT83xTboreiVekh1dF2V0Uk
kwIOif39JZCOBryNNu4mJesB2Ki/mbkgQgegn/LzcN7VIrTvKIf+1Pjz8E7NKFWU9XUxvAwxQmp6
V0U4xCz6BFGgIFqatfjJJIYTi/cIyXTvwJTRSGdzP2QAXgrhjqZwTakMNqZjql1p8mn46CfaTo8p
kzpG/C38Bk0ufgstseklT3zhlFVeWj97qNQrhaWEaGAJnhHzQC9izMBDwzgkfaVgx2vAmLPRCwSD
RN+3NY3RikEaKEFWrGBan0nsL1pYCpgo6Mxa/lu5wwCkzlUfEch45g2nfYQyvC4OPCTNxxobNbs9
ljuptHzSHOAabUVL9I16G2JDvAK8Y7AzTwU7taqjqtWyBcPqNZHWiIr190dRI42jb9Qpxu4dHpMV
oBJWPfg7w6utP9z0oe+IOO63qwsMFdYX+0ikt7X68Ta+xUom+KmcGrOyL0o+6R9xOvUA7X95QkCd
k4XOQN9ckOOoLqyli5g/6nr0rapL6f8gDNoXJKwK3GqBFKelU9FkWPKod9ulIllUPP/IL7hK1USo
EWVTeIsP13suDbSlu2ktbtAJ7hE22hyPr854VskoUr1Mkq7HgzHa7EO2zOYRlB1x0IcizHSX8Oj1
qK4WMgxY68sTgxkoti1qymymMaA/RUSrJP/GOJwPglT9WGVhcTtNU05eUngQqO7PGcqVh1junM4R
1pkIGsGwT6EY7/kc96zfCLmZOwzjXlkSKF7jIS3nHp3iIdzDvam2tJRyKqRKsGOW/8MgLSGrS76K
5OhPDM6YrQDe8rZiJbh+DQqtKlomZ0YcAjWcFXQDZFbctJwqTU6V7TcfZy/rqGjwuWKbolUVwJp0
AZSKziPUDXeGTLwah6042zafo3MScZj77J9azqXDpYSSz2mn0U7r4ASadeP+YTZOZFHa/rg4J6l7
YW5m6F+zG9dwHsbb0sFMj8a3Ryq6THQgEZk6wh6PhL35z38lXQqLZVjWypAdxgoOevQGYtUp46ri
pvXdfCG4qCB1+LEZOga1bfT3YFtisMHbYJAfofKV/oH9QBx/9WnLZzuZqrCkOFgb+eS+C5cUwe8k
wVDu/Jg6JjkqidP45pzFS7G5p4R8r3vM7Wk0xqbprhiQvKO5w9+sxfoirvTNsImrbZ6r7Le6k1AZ
ftdrSxfJpfq+QCGm/iIioUMXO2ZQBH1P6FVRhdCzFX+KaI473UyRqN1LiegbWipstyTE3ulOlEX1
gRO4mT5I7FV4rAER0F+aUrKA4ywQmanSt0vZwIIifppbDXYTcYpx/JB5wJvE89DBQ9X4oNnckGbm
VYPzlwnSy7Nabx6yrBvG3MJl6uQjVePHbtTD+oYYmzILVs+Z1hLDecwQo/p0v4B34tNlH9wD6O8I
D9oaIi65adF+V7NPISvOsuAz55xn4sLeWldZq9kbVb8GUeBrzZ4C5A74m1695ww6YJaYzkNwRYdi
Dys3Whne8atmLMesBISgX9LA/DnW4AZXGMP0P+TaaIkev+6Cq20oE4hbW3GWM1XaZhxz72jHB3b+
goKpXlThI5AIQsz5TETHf41AalDm2IrzIQiNGdIznCR0tNMn1weCO5xWBB9e/Ttea6MWzxpIOpAy
OHdlcfjTS35wei/tekxqdd0lnP8ZnsRGHeUkcGaggNyBlN3gDt11Wf4rO/OE74bBVd4hBcjDzCis
OETGVlLp8zVXkXjXehr14LTVfDX3H6iYq/X8kS5qv3ZBoiy6ZWhRnQK8X+5862QQoFl47NKyllP7
/uvUCpuHuHYKXI5zqeIQtwvWOnpNAnjWcmp5kMmIlET4nnVjUS0SY7hzkqpUvm8fiYODsDVZGOwV
G0WGuYKR9ChKxaRFSQ2+s65TS0zB5uS06XG+3RaQpBeOdTRrDVpG/CtOhysUXbyXonFOlTJ7gI+b
aItDCKdsxe71KDIpCa8liCGMgBa7tgpvIh1xwdui7hQMYafpsAF00Sky+0BdXv4uUiRNSpJdIGNc
5xtcMPH8DpiqFrYlDy0D96Af2Zno6LZK0I9NzAEDYDtV6XlZ9RmBB0XEuJtVgQOIRCAByVWBigzr
+yCH2H8zHyyi5rYQZx3HxgAOOENcz1gPIlWvweUIe5HvvUq55Q31dmKb2HCJkOe+5m1SLMzkJUAI
J6+DeI9E+cOywu0IhieHruAf1+j3DLbC4tL+QWn7D9qtGxaCnB9SgjMIda3B5Yl8nYgWMr277nIo
2yNzER+u7X6IfLgs3jvDp6fNtoJLVBrrH9+dcqnPC2joDkYiLq1oEBxpH+XLVEhKXx/jZSzha782
YdVUS/3lLE5zR5hJ2J0Iz2QwSJ/X5lhk9C/aCbumQ0JPxZZooIwmMGTF26uTh0PJzXr7IwlC18Ae
7SCinpGy3Xinmjkw2z68mzYi4v/+Mq/UC0j4cNLcwidTYW6o4FI89GV3rUWhzB4TklJOknRCIISX
Kv6AKveC/wLql+G8dRLTLwZXL3jtc3qtO03tne+JV/h2wG//fEtEIFgr25YtBOqxWkryeHMZvYF8
QarLB5aFJoEZHfWr/LUJCxc732R/0Bx28FcRFMlGpiTUYJAnAjB8Y9BILpplewe0u0AgzEP2qIsK
Wj0Z5pfZOupmnAV7P526CUkEoApX2NguCRMoIZh4i9gT6viJuDu+tkNlMHCDsKzqWTbyhTg4pMlF
dGS60bIQhbiCmcNUE+/5q+PrmuKmplh54X3j3rngAXX+XlJ+ZQCOW9vBA8aDQFfRi4CuZ+kYAaZd
j8kVrwN1ydllQCds35a3+zVSh5DRsx9tyIP6jSRZI62u1JYgzW1dKg+jBiht23O2VfB44yLp5HCo
KVrEJRN3kM4DD0eqHtVesWGVhdvPsMKiwVcJVsbjgNKP3O5NcY0BMfrryrtGWFiI43lVLPfc4fZd
j1tQV38s1oMXQaOIy/FV6AbCCOG5ixnLN0Uz50ODP9fNeEMalDKcggbeSbUdBE+Q/NTWapWve1iI
2IknhPTGqx+hPp8KFDvW9kaY+SSP9JagncLc5WLh89/wivLyvlTOvtUGs1bXazv1cnnAf/5dBLJf
CTnzZhkhmrPLPWrkdVVKgKzVZX9LYy3OjNd6BbLN9t0brsXlTkUvLafpJ3BBo27DVjSJLh9qS4R5
qHBjC8NN7kXGAIUnIKxlUNwg43OWYHi1JL9qg3+NbPS6pxvljX+INYAOBdiiZbA6go18rBw/aBWi
u7AMYBhkD+5F37CnQkARPjrvhqV/fSX3l2YCYPGnsEz+5U4BFLOdAw73uhvLZGsnLMV01rc7AEGC
ZYBY5YLkJ+ZEYWIJUJDoCggessI+NnWB9dbd5KrAgnxdeXKsuFNjQ8KuRGXWxJ8vCpLa28buC9np
tUid2GpG6xAbIUe4U77P2thmO2mmeu5rugnQ4Zp2wb4pK9Pf4r+2jiUteePf+VXTe+6TM6fBoZDB
sFtwfALMQqv1Ri7Ovuk94ZeeHjqJ/UUlo9C6XPdKxkHX8Vd1tGOLDZ/dTRZaFJm6Mk87brhc+rMF
jrZzfA7ZIwb5utoVy6vzsiqcUp73Q9yTb3A2Fwz7rAbPfVZy+0hcwhWu3t6ltw0R1SBZWP8mEWXy
jcNKbaQ8ID2uz7O6MQ+f5PJoBB93TktWU6S0OBz4yAHDn/cuu4m3mORauaSB9TtfKRQ7KrGwdxjs
IngvOZZr7v4VO416Gg65Q1zH/Iq0zpdg4m9MPc16FLBDeCaRjho1c9s23luakxtC4BQ0tsNzu0Bv
5EKI1BjNhLL6Cb3uennIzxXzJJYQnTWaGU3mNG7vwPzNpQPFOEq1J0cW8mG2U/10TdT0Ldaakhck
C/rfvp8+zcTRpaNWG1njj6fpLFloWZ4z31xmYfnyZwyZC5wQ4/ZCN6HD94arMMazKbyx5cYnj4Nq
ac2hxqjYFykYMi70MByz3bBYgypVSyOuInwM3AYzA6+jpVgUJtBl+755ShtuhhMbnA4/FfDqtePN
tRFEJrY6bREXVPUi0tZP3XCHKAHy28gaQ5lLRgCawEFk3dmqYAHIXq9VBfNPaozLYbbH4ihZ8T9S
WCVrVceDniJ41NlfW9l+bwYcJx7A6LGe87EVL7HB/aKXN4nsCi9QfapwC9HSlxL3oNXy2m7CI5VV
dCKQ+TqgfkLpY+3TnJTnxgZwwZH9SRTAKA3Opq903ArkIK0gzyAdtg9Ys/VRH+Yxu4c3n/iQ+qr3
vd6cr1rDU56wxN949SrITOfCdW3ZC+mH/f2HqjpMqG+31TiKPfxI2tUS35/cFk3ZLmv82KZtUNBO
DwNo9nfGqb1ZEnxKo5Nuh8JIW+ug46XwziZcGzC3sXRfbSkzZr8qbi+tEQrwgoi3Bd5aoXhP8UUy
rQWp1PyVNHsOERIN3CJ0qXDln3KeDvg62jWboTr67cRdbpg9gkTCgG+EFzalnLd6V6eqlPae7LOP
AxBpmkZvUZnnN+ORtVsLP7CIPk8O8Q8HfvcpaaEazPIgFHVDz+LtkyEHZC5SEtpvlvEEkYA4vifC
Yghxuw2q1I0PrUwx06PkDVVcdw+hdcGaHF7t7Y7M+RA0IK9kN5TRElXjbf4++D7bddnA9YGMyBQA
e4b6xhbe4bXKenK/zGtgdCv5ZJS+bU5mhJ9FKcyVz62IV7OUSBUbgqc6IpVWMrccLqxSZIXTFwwD
o+OyEwEYL6F7rMvGzdGiTEL353aIuuufZbJXnuVv72eCDwWtWMALlwxUaD5XiZX6IbkVkMuM8Yye
JmaX0c0MT0wkPFmrYT1xv76td0hB8w88H2X/zF2ssTfHY+KHri2OruhLdephUiE4tjbv5wSzYHEy
N9QcmStJG0TjxzHF1Cur2K5u8IQm9jljg8bTzIo9m1ysQ+0pYmCLZYCOp3sLkAz3xXqHbtB68iW0
se815c9IL3Ns7KiiuIUrVRGal02j2LwOvtfUrlNBRLU6ykA2X8I26mOZth422WbYhJIfVVHBXOBw
Gxa62TGuldjTIsgm+aE3QCjbhVNt3Do/RAhSVsx20M0iGr++uV5pZvQzNQwzxbLlLz6u59c/OYMZ
9TI3KG7hxCt4VUBfqd6b/oKDWjJkWAMlDXYzRjuMms12/DUJLWAbf6Tg+BTh0QlrH8QsBzva33d0
Nd3Q1NKDimaMyOeJ/zMvpqvVpzfBStcZwJuga2pTS5RO3WFy8pEII76Wh7NBUQvKHnYWAKR8aIFQ
U4G8CtfJVpR/6ZvyUdUvdLsZJEnQiz5tskAJUni9pW0DjJL5GA2CBZkz5X3S3Bshk0Fyl2gOIXzs
eOM21L+dvZ46GMzFt1JlQvRTkSY0YBqiuS5+ejj5TJvE+iPiuze32ifXdgd9EwafTen6IOA9yOdQ
ZvxKDJKZqkN7QXULAJwo5QzkXqiyOPeBS3IGORA+YXgoawIXncwQF7CxVCH3vZrO1AucD63kReSj
sefcyn9eJ8fdqk5cnMscka71KqYE3VOEUI5yXB10hAJ/NMVyYocFYEw4yHFIV5Pi40RJ6zGMumJT
eXD8lkBqx2A2ffjWeFqBwJgiATfsX1m3G/VPepa/48UZ+0orgP9lHgEGZEW2LhPt1mNiXkZfcM0v
vUtI7Es1tj9wM+8wyx6S0YGQ7QHzwtLBL4lo+cgWRsheyyDZvh5sZWDOocsVhd8c+U30YLaAe7M5
u57q//Olgy93Y13B1c5uagNJoBFrrE4v4ohFabjrZODxHnsSuLY+PsDI6GcX7+ap47PWNSanOeLF
9Scn01b/p4uL4UNs1P+6xHMqTzu4JkkxBpybxkgpz5T2IprLtkBCXHYo4UK/nYn8DupsHnq7sWw/
dim9aJ48s+vVX4z8DhnGaz9Yv+3VVfcCFjWWYjUQxOBC9cHrrIfl38tbZXL4+1CnRrYLi+nmcsfX
GFCuMKxu1vaIxHQwLu4YdT2bK3Tep2Ic8VxWSJP5rj8wlqXC+koVIfQY7qI2KXVi3ph0arocJZjR
cUWl1jH34Ot0mfOupfqpHQWOQSmwGflsVXzptxYMcMJW+CyMtbGqyzZIN+9OQVjY+tgGiNI/hG4Q
Jn68N/3qtFB1RsG7aKpDsee86bdsJyl2CHATCxkh5GBfcZ6YOy/qzucGMXleeCvNg/4GAjJdBU4z
nue0V6vpdiA1NSoLU8WPUnx8EAJFVRY6HgE2c5dY6CtLjI92XiJ/RsDH7OYXo4afZCDENLGxdFwm
mkdFSh5TuAHj21+kJlWJSp8j4ndjnQ7xvUdLCB7wBddaZ3QsZiM04ezNsX6nQeAmdjxZNJMpCdkc
iQrgu9PzcsPGi2+Hbgt0QNRiJd/+Bxl4UpQYmjpmPU9oM2yeJ1nO0BakKr+tAgSVz86+QNfkCKn6
Gjj0MTYAAM88aFG5H3yM518oAbhru9gDHa3XQTPYHYS+IYhUrXbZnTjcwbRhnWCTJlWvVzT9eQi0
NvESXiXKAUntxT4/eIfnU6mkeuninz/RODWe+DlhI67obJye1qwiLRGxuImTs/NR9cCFtrq8V+DH
aZDXKd2Z7bWG3cOBpvNyWPg1w/nWmETNsZCGq8g2B4MPN1yrFa9Yd5tXIKSvxefxolLnXDgJza9N
z2CnLYY2crpYeNWd5kh4vCx01xu0fO34Rg+xo7P6oAVduZwNjUKMHhc2Qw0baDGOD843a/04YJZ5
rh9ftRzzEo7m9oYmrZDiXXNzwtiON7Kf/0OUCS7JmKibu9B2MpNZRE32+DhkHiWudaof2QVuPUOv
k8QIARpxJBK5tjC6iDC1bTgcZE7+uDWX9q+/gf39quuAhA3Y8gc/pSUNQHacuGktoHKyVFmD8GRi
SPwR72aZTT5gK7rBmYkCglnd+nwY+l/54GSbOi355UbL2aymk69ZS9oD0+Sy/ISdDLl9qsmM2lF+
gZGLIQHFa6Otiu0JXsTRkxx9al0v4p/SCouI4dHmloA8ICmQ1BpOJhplFbMyzP+tU0NZSl9sHyE7
8JBWkb3o8z0JSqyL9UUlTOwVGG+Gi46DYlMsDXJmAGXFm2/KWlNjM9JetfffWSem2ih3HP8ojSvI
gH5atyh9XK1kj4JVEVDBV85jRB3Y24YEz9JkXrxgVR0dX71MIIZ9A3fvxFOzKUwWmngTVJ5zqdiI
nKYfDOyGGqTWkfhnbD67tn4mNz7yM4kia71oRL7YdcGWe1fxG8tHGXNA2CEd9Dxnb+ZszHpsD3If
+YEz8AC3nXIC5nOu3JheGOCGFt/no6QvRZ84UVxqWQD4XX8CYnCtGOgB4V3S5r804WX5CzmnvxCR
+uJZRf43q8EqEqe07rLnT07B/GGoXJft+f0etju/NNxECccnONL+SdUWAcX2u6ULQLSpF0DGsFfV
CcEKMY51E0lfs8xY4pxoNJQCw8FTFTLeESIZB3LmqulnUtrGofU1uiHIfnngxUhkepLrOAiR5QYs
PkCNkvP4+Ln7rzPKKYk2QYQdj+u198nK3kHxqZNFlTxjCz/2Hn3IDiVphn5ZeTV3vCWykoKXR1Su
RJ76dvXJl5hC9pklgLcnN52VRDabZ776xU+qBShkBBtX4WbVFJ+B8y/iPSyAI0d9omajFSjn58nX
rYXKNdfv0DLKt4mfb+3pgPylhToVmfsHPprZtW6qAe6bp+i9cOziry1pvgkJaq9VSA5nOzZq2rid
d3Fc7pjazZCs3S4GV5e3YuloabXtrlnByBn/PV2P6HiUUbqfWHtpz1YtEslEo/2E9UvTlrfEGJ2X
XYKCpywW7JNUlHO84yPWaCV/c/7tKlEPUA8QDyuClzaeXuBFl76+2Y/bmcLzIKBgDS+7BrqryKVO
OUy2OEh2qvPd2Gq9Ya5+wkUzl6QnmRvGhhlfWKOTUun+Qowzf+AiZnaK2WI4YduImSX3CLLNdt+K
u1X8I8yXQgM7yHuZoKA7WEI3d62xhLSWWDK9gaodqod/c2numBpcoPS5HQOSHLVaFLt3q/ngOJds
+nA7WSzfBnQZa25TIX+7GZaQnEedFjlfVI5p9TNzCPKXvdlUrbe6Ft9PPXBr601M2AbMYDXmAn+g
CxlmJFarE+l2qqhJQdoyw+ZsyTUiDKODcpcU0DwodRnQGYX5hCBgePIZ3Ls6ZN7+8v16E0MK4jQh
R1fpd2/Z39QFetrmtgVn8yBbRQV6Dq+eU32uczn1vxzOF7krgvYn/XQaG+dc2qxkFKOgoOFV2VyZ
R2eGKBR4Op+/4MnmsQRzaxMVebC9JB/cZEpKt97ffhw42QEqOQVLr2Y4MszGUaLNLoNFov6IuNXk
vz91ghr6aFTvZq4DfvBJ6ZbFFQDATGfId0o2Y+Lhs+jQK1JzNIOpUkBqsrtHllfG/pvhfv9hq6Nh
CiUpCezTofY2TO3PDSb8qqIAbuUyQ4wXw2/JkXjsc0ohbjood+LUO1fi6ORNRzWU85T0XrIK1MWN
hnflwXQN7vIEF+5Qri7qsFPbrqryd3rRd8zC3vYIC8ZZeeXCN+Vl6MP8VNh2li6HtKKvrSGakgq9
nMni3l2tCwdogwVf1QbQpZiqWpIDNd4RD0rq9oZYjEBnKLJ586MxyrpRVc3F+xhpTxrsbbIADWYO
PbxuPnWgCOssSoUgz0AKsTlAdn0sUihXxY6z9xgMh8VdcpMFFyb8ebHCfsNyZU2UHUztQOiuiyXL
kw4yKui8TicGbcd1QFU85g0sw3kob7BdRn/wsrUvhBppcmcZ1pFYiTaEdBEOPm7pWOoxd2x/UnDY
CYDPvNO9zkO7Scp0JIANV8mV9zBnZwCzT/NKLMKB6OgeP3+0miHbRSRZcLmgorY0khcD3Iem0eFG
P+9HcOISTM3kLYuoawGg5ZCYDzEyRKeE9GwblUuZV47bpA7VNxkGt/p1E89ec9IU+ozdDdT+Syja
1A3QD0sRASN6neFJ7v20zzMFyesvfBEVRWmsKUeGzhkOTwNIHjkcy2KbGD80aGEZZwFxMRPwIz2E
eoMitXHFc29v5OMKPYfQvNfO9QMtH0CLcrSNuRXY8GqBpPfvlTO/TTz5I1AA/DHW7rR7t5DzQHaX
kwZL1awRGznMomtMBYdGxACA8DKKZSgQmsk12MWxbur3kTGJ0qninOOPiXHvcbbkaNqfO/G/JRq6
ZRkous7+Bhju4LS9r8hxFCRpV3MCbfeUFq2XIelhkCPuLkkw3s3fhO5+X/5QOCiXMsqQt1wAR1Bd
Yzndl1G/0iaLzQouKDu07jNTYbh4ZJ69dazjQbIpZYgWY3tqPxv7stdOhVsKOqMRrWsfhqaBLnEh
MSWtwipYinWE3gBpFaPK2OGaqe9Ta6ZDHDFxDXBPe1C7EHJuIHxgI5SYPVpYxHcJOEWEAg4oSxTr
AbVEbHL2kk0fRiQHbOy19LSqNep44m0+KTAxIAP1hsoygqdFnx7oeTqRXZne8QhPPWYetSKNMfQI
Km0jt6ZQzBeBMDvjG3t5iDSPlaCCaHVZuTMXNKRJwMxow18lo3/P/I6w/SE7Psa0ufoAUdhICGQt
eXXHJu4GpAc7BNS9xsIwywWPb6QZF/eqrktuQ3l2vqqB+mmjmpWOvSGpCUsQlzjWMGVrdcjlbHlY
1KnKmEtA0Tybwlz2WYxEKhNoulCHf7y3tcj8r1L1AvHA2rLXxCgVMTZBOCRp07fylxCnAc46+DKH
wnZUvJF2obGMcpJeokbBEMp/M65wk9BVfAI5ocVEaVfmKuWC6R3MZCHQRip8z7+GXR1yklvstxdb
mPc1+fslRD8J1EPH9DhYHnNUu9qF/K728dQj8TqaYDQlKFxMrwSwoPbhuJQV+erIweS5PeI1Kfjj
mmsYpvw3YstZiGQGurBSImj/vE9GcB+1nERQ6tbtK1WOGBGDS3mlzOnv8HmWWSxxOVVu/9DA05GH
CVpYmUQo8otwNPWc/aJJ4lWJEOoQoqTPu1wubBa68lr0V6eVsLc0VPjZqBYAaziAkrsGsZHjrT/p
LvZupmX+QQDEe1l/BUY1ZrZ5exA/u+wNRglruGvHGQBwE+t/soG72y7PidrQ6RpQ8qDQ1/vN2XLT
9tt0q+diLt0NqpHpqGjjiS/XGf8hq5/XA87YD9ysK/AdLMEcoH6al3GaLrk9LmdaoOZnPwIzUbMw
MGyGsmWu2Ealihnaon/LHz6KwtGq8qjex590Ht8O635U3GWRjgVD47zttXhgNGpMUFNF6rV+0pqF
qgdB2Gvw4kVLGEwuNOnvaXonP+Df22OdrD1enLoAp3SKugDoPTzvdAkvFMkgkNE+ijUBJtc0Rr0z
XS+pU9WN1PCw9Gwch/3k/eZVNDNZPwoWQk+P0jKXK4pW3Ya0Z9fBouVzSSeAP3RR9dZftXVridos
wvr7IEZ6K9pu/75FBPBhDLeUD2C2AGTs9PiZts2O4j4EUMkd8PmCZwOQxfaDhr9JAIokK8aOTwfK
CM7oEBBmjis7pi3kKezP9I8Iy/FX4waoVnUAN5r1g03B0y8pb9GxjNXW+bxGN/sxCRhe39ntwKzz
GUDNuzA9kdI2Vtzdf6w75YvUog0PW8KmPP4zyud7H6ox/91eIB+0a3N9/iXBHkLaMZ5NReH2DWYw
fGmnLTXQIMwfSja1hyKSVJgNxM2pY8g7ulrDihMNGjjVvcPBzeS5wJ37iXf8GOeQPCQvJuUGkEvY
UeElvet+9Mhh1KChNvb0xyTgMtJjjeuO9KkYVycLq6F2kPIzHZEY6iVLvE7Emt8ua6vFr9flgGl9
LQMgJugIZ5TrTykHUchiTO/N/oIytyHa6RKSBlL4rJ7Etlqf96nIeyl3onKbj0lWM3JrIan0Oub9
6lhTqKLNkvAdoI8HEwAuKBWaYp2rwc0+lwHfIMp35c/mxbqJ+Krv8hZgivGzWLomDYhQ+UvuCM/E
rrqaZedOhpn/In87YqMlbY0pXcoxYfOiJfMXXpjhMPo1XGZCXB8a/UqhK7khEYfvVggeSD4Zbdsf
vdN+2+UMOtIcPI9Fs/NKjAvFHBIpSV3O1l+oRoMHn6JxudBan0R4rfsHLJkQWYB4qLyNUP94R0lv
6soC8d0z0y3JnGZ821Y1plmw+KZJDm0CO8KcVJxslbwKHKXGjibg2p6iXzSbbmgclGkQqa5YOsg3
ti3robgYRGWqM4XeRMdiiHvWmEkA3QxOt27VN61YTVVG4pjvYXa3kbjf9NSbvKofuT5rkejDEAeS
nrX2dfdwPtuPCodyF3mvM4APz5sotMXNsCnyHGmPGwL7RF+ImVL5MpijZ3/ptDRMzx75KiIvt1hK
XTYuY0GRFcgB39Lk3P/YrpS+mG480TFI1LmFNgX3ZCt4mrg35pHJwN/bT1e85/GEeOXkBwJIoAkF
9BjIs6QW1aEo9cZZzV92Y+eMmmZ2O3inO065aTgtfk4EcSZVxH5QG319tFupRQCNc7fh01tgEUUR
MGLUHSajl1EADR+2lf3mHmkPTwpTgiArZvXX8I93lqHbuhcWwWV00OUz9KcBsfwGbJxRmj55HR6k
2MVifLVu/YKGo/LNGHTaAX2ASn8OLz5X+3fVLcIL3FB18BYa56X9yhZxwBC7YLG50EEgUhVmDQj/
IugMEmJThTDaIVBIhJbXc1fsTfprcOIQeJa6wmfcMxmCvDBuI8LUrxdaTDECaZqIVZAUY1exs6FK
IWBOVRS5J9i8PyN1S3IKFPvlkfET/QW4UDDdkeLgUaME3jX2D5nk77DKFq+dbU33losn1TbhiP8a
VinZXNhqnutiNG9R9eX2jaqeh+3xXha7GdY6fcf+ZZ7NGzVJdTtI25Z219KwofFq9Bj0I82J9akF
EeDcImGBhEHvhpUnYsw3+MtB6R2TD127LEYA9xqKvAwot9Azt2ISqV2tv2Kex96pkSlZn75iQwFX
WZ2pigHWmmOZLyAPg13HaSamEGpwpH6eLbLjRsFx3e3m2ZQcVC19sPNo78/RHog/jGk36XnCpuS3
NtT5Z9kXou8kJx3F94EmS3891DGo99fXZPrP/jNtDl/H9sHcxaba1VXlcoIhHZWrOAJV5epqhk1j
fd071s+VepHPlQR3bZML8nZZo+06lvf+FmipjGd/Tiwh0quJRFe+nVpbQi6mViVhnFTyVl/cy0NO
cU1Z45mH4vT/pWOCpUuli+xji49m+Okm9MEJeLxINO0jsEWsWeMT6PKUFALgU0h3gzmnhsE2anBD
6xWn4WwPdBny+NEF8od6L3te1eG0rrMvIui9Qez5MQwqOwXhGCo6kXT5hddb4+PrPkip03Pzvwqh
C2uzXKmLrNUmBhPqeER24oXmewHQpJBLJIkVrXX1jV1FRzIxhhOmYpX+faf8XzsGpPyYE6MhfHqq
Ggw2GVnidZlAXs55AgzPEOFiKv6JAap5ZpVwDevyR0hqtnerIBbW2RM69DFgpviAHL3vDLN1c3Wx
MWubpCUldZgwhJgkxHWC/1RP2+B9WH6BLTeZ8CA0gWlZqkIZbkvjuH4FU7OXQXDiPp26gg/6EaqH
gJdEhC13+Irbn12I8wNfUtJGEv55duqtiwRFRhupKdkVvohuF4VLJ1uy9jyvUjoGQZgK89Ga48q9
8uUnN1kRIPv9O8YpIlyxxRs5iFEwsnC/8DRJYLGQzInHcirINUdjPRixbAl/VnKdp6XxAStc0+9W
hSxPe3pcpSSxt8G8XDZEASt8M1t+c0/AdEOtMMLuBmUtWapjnkq/KXMxhOco87iujlawYMqdswyO
Hsy6L2NPEz0npG5GNwU+th3d+k73svtexrIoGahO+KhsyIv9FyTGV+DivbKU83VXTN7wRB1LYInI
PYgUedTJ13PsKEzS4Xo4a+oxGuQ4A943Z/sLCAqJr2iBe3XVXbzeobUT+hZO3J0cg8jN7csQK3en
pDpcu9A9onBU0tiAc4+SsW3WqrS5JF1g3FkZwL8lLuYWKLdBchYlts6Jb30KPRuIfHhRbqQTn/n4
ereEyIkjC4WEwA1TnWrSscK0vK934oMrU9kf4AKxqo/r1d/oX0Q1oE3jfKfhCNILMqVCjP+o64IM
J1QLR/8fcWHLvCCJIg1ITEhC740shJtBsc/m5U4jnnVJXacbo4MJN+nkb3kO1A3GR5SCdVvjDNrY
L2Ns0v/Q/5Sdge2qnH8RroDCRFN10Iad8XNdb/0Ws4zpICDAzcOxTx4tW1N1eEI7MXE6m93YUB0Z
PBck1KCPGDVUBU6lN3L2ev6voarjh1QPUhkgj86+ROuqzkR4JjbQe2uPQ+IkoQXIkS2jHp3DSJeB
UpC86muUraZryDxX0UfdHJkxu2cJMTA1Oa30377dxSwJBuZAIQgLDDdAnpVf6vTn37MYboJjD8fy
RlpzTE1wdJBjMd4I3Wlg4vQqszBVuEI5mZeRnRZxX354i/GNedxwPVBkWFMjEurCgGlOeOS13XWz
DIgO6VEGQUYAC30I1SFN6faVYyzZ7aQzIQMykDU2NqkamZ/Cs7j4Bf2SPZ1vH29z27fEljgv9Quh
v6lSft9pVlJqFvVSQGQM1vTJu1jBmK9t1Q2g83CuSm5ilJIH3y2zmDko0NpD+D/Dm4fWgxPEpBC2
LR4i0CwIgBfO1RqatL+CO5q0wbD07BXWYDN742VHD3UE0UtU+O6+5cn9gPVd//PIHKd86ZPomqlo
EdekxIZcpB1ZsxIpnf5eXFb1FhQqQIVnksv9bxdSFwNFNb17FCklT9CccbgcHf3pAubTITLFqlk2
/jtqo18tWJg3drPEal+w3/TcNlkWRp0e3kRffrGUAQ8nPzUOKoaT4BNOCcID+TUDsngPmr3nSo9N
Fzgq5u513QyBYDrTwqUTGfQyRi7UqhNutOJxhz86dSZ44/8ZHlEwZP1le5xwQ1WtOHDZPzgaWJRp
7l6J522blIXEJQv89OMfuoBGyH4OQrWmM7CXVON3nEn7Qp/bFj/G25PH1WlpXBgbSUIQnoRiVdYq
V1wZCHtMGCKeKrTqDsnvona2ny9+1mfwT+D3cqtNG43wk5hwFBxFE/OX9cS35xhEHiGG6aPIIQag
e2XorA6zyvW4DqetR3N4Wy6omy1yZEWDXYn4OpWg+Kl0HpcAFxfT4fJP5tRD2IHe5o0jmOph2o63
EYPWbm3mINNs2ArumK2+jy3AhvOgYKQaOm3xOBY2pp7ObqzLVMxDvgT9LV3NavKUVB3JRG5Yf5zK
nb+XmMY+9b4H8cP7PpncaYvNdJwqKeEP0ysdoI+Rf0YA2hDuif0ZTlzx8d3/ElqzYzFIDH6dJ7Nv
rXavWE7/C+Qh1T24T379qM+WwqIkMsGq0NiACu8dgnvh18Wal8S/X0m5+q50hAGkAaoOC5l6qaSs
FrNJ/4OwSoYMkghgvL5/H+S4oWKXS6y66fRzuWICfQdyj3/f+XNW12r68gldVo+D2LS3Q5yF86ow
Z4IPP6VjG/EO001vbnTLIcbVsy0gIg3T4gxYIKTlwBKpKYJWN4MtND/Ic22S9R9WkXajm2Dno7Dw
BxGQJMy9aJMkubLTA+O9I8OH7e4VPA0Z4hSiGN9aW34P/kiW5KyBQlK652l+8aDV6mlQu5+y8pUC
C6W8e07nzp5Zd0LMYW7dzQF1+epw6StrhfV5VFgX3hC5ruZQ4qFAiyObfSMos1C0AvXneKum3VVq
tEt3dcKMYa5a+JP6fa6ZdSsnZeF3eM7347JowV6wKsZKghCB1LwKeTdOy8iLQounNKu1DJ6syhez
tiP/T0vpH41g0B45lMYubXxtbTxm9ZdfpxqwTbDEYDTP/BkgN59t3+GKsQXrfY6PWTrMIe9QJ683
z8opSLOd8pxeQmJCrwU/W+dKrrlcThrBKYhHmzZOJ9LCyn8iJ/8UQGVzSy5p2F1iMZNdYNEfp0+6
vaNUcBig78vH5bC4kVbb0tHHhhoCsKfU23HJnjgT0V1WLHncv3iItVpsWVhqyQlBeWsVeOs28i8p
9bC1fC0MbE86SHMSCG06vNMzIoKOAXIpioAS+LS+WupEiGhdElO2q1tHXNGnHPOfE4x3suWCWulR
TAKMQPXPtKjISc62jT7P/XBhQ9wNY7aNm3vUBXPqLtlWmE5hOm6XFpR7lmJDQo+JbyFUocyOf+D9
7SyY3Uiu9+lBORjYcPxjgHKIwbpHySYl3tp/MmmqLyM9fqBNpjLvw8KjtHgmicXawDUw4ezq5bn8
F2Dkhr1W60JqvxPXudyAxbxxEyJc2s1bC2nyTC7QwviAvy50YkMIIV3qEUYr2L19PNMpFYPwJ2g8
fR7AEqEUHd4ySGLNshsxAN+iqmAeiFqG8uzmJjHh7AjvTvD72yzAPkwKWgfiVxBYQK9XUiVpSNhQ
7Y9jqjCd0nZU3iGz7J2qUA6YF2WkQ/rAdlwxiKCAYGWt3dMEd9Do1hlYSKLlDIEhgERD2regcKDQ
FdZBHkekC9n6kBkMWkrpbaKEwgOgE+lbwctAJHoIEejRFxWXfleOb6ZlEdjZ+XuA/6zcENTDOR2y
m9mCbe7F2GMElLdistjrsTZkNtdmt6mq+07U+snoUnMZ3cXZ8h/fdzI6N0CpYSZqLOl8CEAsMxDD
NamoXmXWxPzthEFE1zl2swd+1KyRT9lylEGH2t4ucyUdO7GXDihheyW0puXVHdl2IaMPlTt++9NU
OamoOzamlruHkXeT2JGq5V1SJHfexElmw/z7oZDjbjOyu0OIoYEVuxLlhlk6ljHZ36GKJFfMnysh
syBk9MjHtEB/8/1Ll0seTxKmOrAoqxOSRSmgK96iyGmNpPTv3XApgq3Ahvt6/JfBPXtg2nmjx40t
MQh8SuE+qyU7KTt7pC7RqEy0G/AYC4YJg0FLSiJb7H20hk3ukBxYczX+SCLi3wPKyd3hKiR72uh0
wba5dRL+vkepjCuZTy0iDKObPMEsSuPN0JHM1yg+RYtYGQDDsrjLkRQBPqmVj0KmSAVFNTw02kED
+0POxhr83H/xT0jIIXzbeSEG/IFj1Luz0X3ELuSOhNef1fIcoh1cHxTz33rr7ZS976Q31tMk+lhF
bA10aV11fb8d0kdR0M4oAKqw496XSeKTeAaYCpQjYoLvzO7kjWNWNzhsK3WCnwIdLTew80Td3Mnh
NVMDm8OObqTtlqkmruyFpD5eVM0BsqDjPHUROtElRnpPBgzzJZzzPFpYqHvF0vn6yNvnPWcs3uXj
ZNj6nwQRgNZmD6B3RVZZxsw96BzZ0Aa5ghQPP/HFDPv8vrtFAy1AUGxce2gKFe+U9sTxs7JrISKt
dL9ANQmAI9xK5+dC39UaeIt/X30TIiwZdS0BcZUiJ9kx1Kt6mTGmoMiDurXUJjwJu1Ce4y/0Wojs
LIuYQ432BH7FBJKOAZYK1lVPjMp2DS3WaDJEDBLayb/tqNwyCjKBpvy13QD3eefSpd3ZT+5jQqBy
KMx8C+iPtDyapMXSkIxtsGO4bdG/mKTEX8Tivmf3cY+uGYeZUb0qrVAO6L9ub6M/pRy/0hFTvURv
YzEnchWk4MdImCB4Xlts+P4niK5d4uvRUBw+pDXCTQVSxtJrICugfDdDSvd2kTj148HS6txR+d6r
5LJ4hfE2+PlIqGitEHfwhpwn2BMU6D4JoMxMpOSZ4qO5t0J4/QUblBbpApjKATTYogG/Gx8j5kgg
CgXWFPwBoHVzzJa9xyhcxGOTO7MuYSs3DlbEFXLwaFycPF4IjDbdUHYeVoJFE0y4CI1y1fhZzaKM
KbB2O6jpYfBdLqWI16Z25MPlAb+IEtbqlEOWZUHHaAuZlvq8dDwXYy+gg+3wAvGE/uNyUdPnwvaV
dE2SUZUFpNDKyaMCRQ3uuaaewcd2UWgKCzPmABAyhBS+fP+CAex4HAXrrNqrboE3R2wA6WyylBA8
M/d68AulpJ6jijVpYxbV6stax/f0v0wlegb+NqNfUMTbqfuKHvsv7d6bTPVQIdOclFzxELJFrALL
/lRV79nbU1erRbdAtoOPmcTjEkHDHoEMotck8OFgR7qdVA4dQF/Tw1cURgcVa8SznL7w27vVZQmz
9nnGcBsasqdBkEDUPALHN+6Ok1Hzy0FVtvbTeSHT3v86J0PNBwI2bxmN0WPDBEUAlzN6OMQaxKWn
2SSPmRD2izEKMf22gTSI+6KMVQqqZAKHXAIsvbDnUx21r2uRhgo3C42ejT/9xirK9J9eakqAXUaW
OlXolDR12Gdey+a0HaSkiMgpY25Dz92naxKJA0fl416h8Xs5QrqPpxBE0lyzG29SanAvDH6+h3FE
ykOL9VIf4Xurg984N2Dbkmz6cHfXCvmQbciGz7TiAZTormntpbl9wOGHj6Io1WJC9yryNtS7OwtK
U3MYLLkP2HiangKitN3h0OA22UoRw9GYyo+QacjfqSXPowXAB1NEnyQVTYLpKmPVNNEAQ4nJaLZ8
8dk73v8K8JmCdWywUQ6ZJVtPPlSIi/o8boiAtOszWEeMgX0yTDDOC6Wmfaq9uYri4n4oyFVO5XlO
Duos5kCGfI6KQ68I3WMBJwyeIaElLLY/ppgsu6wjfA+XTdllRBSV8n8YPETlSfOqzAftNG5g+RSE
EZVS4XjgdjbEe4sdeGo7o2st8lnUd2hitpnQkkwATWkuYKKqdzS80QN4+8feW+tbG0FzKu++WFJC
CQ8fnyirpKQHUVewD2g8kAXIbJw9uavElXD9V9Px5DaN7C/NSoH5Dx7Xqd12C+RSn18blVcooFUk
zLzTrOnHmmZj4tlksD4nyJIAV642XvOB3SdBkSTT24Bh1yDWKShy+um8+PZnaYodaQZQAkWF9BtZ
NAEIqBZygRXIdAVQuH8VhgQ64rm0ImXrc17SxC5r1/UDQa87OnxARQiZExz8FXvNAyFlxp5QkgMn
6pNWeauXQAvDinwTWhkyuMcwBXjVDOXLTmGcaIS2OMiWozYOLCfnpPSoywncksPtmUyap7Vfaqc+
7cmzxp2plriTkOHU0/lIPGWwBVE3mI1S/Jc4umjPQU3obyWUBq1A5JlsdgHDypTYY2vl3w8wOvir
n6pVOLVVXgjDk4Gt7RaY4xi5SinY+F36gPwOaKaEZPtaZUGUM+oPmAqFgVcgtP7VbPBjI1dMk2gV
FYc25EcyO60kpX446iQXc+jSZqFRndtyXxop70zE4b9RuTkgY1fKROgrx7tfRGhz03vfJsfzYu/Q
HG4OqZugl8VrhHcipHMONpKaug4VEfgjE7vys1/Ip9dEXZuKi8lYeNbYHl3cOTbzVB2BTDPkbedP
ooTUs0LJxRsZT2kugsJ2xdhsnR4GPEAOTQhtZ6pwbmxQURiGUC41JhEB6es+6QX5zjQcyfh2093t
cQjrLdZtX0Zbb0OmYSipy3gEt2ILVufFyg866en8kVARypILnhV4wLXLtLLIATIbqAqRvazYKhQg
lfcBG0xs1rJO6UtFJGPMz1+0VQssgjrIU027f5A8BhiBJlcns/oN8PGAaPP8JfzyVVsa1txEE0Vx
fqM1+A5if0pNViw9AJbSznAfmz7qK8+S8+jahEwrvWbQb9QrYEaHI8s7CiZobok+D6LtUyMXvJ85
n+6DxxJXQjFf0Ag0Ok4l3Dfnr+MzKLnwE2Cw4OTcWqXVuHcAdJINdI12E0s1K4/dC3aZ62w0wqIX
44WgFnWIzVI9pLibA0Xt0XwgkytiHMLq4RGDUwNexZL+7uJFLTuhfqKt8G0al14A+VoIFgYI+TND
8F/78MLdxg4XCJWD6zpTMtx419WxcKvh8bBSlVGLNbht27PpOh7Zx+c5z8kMBM2i7/5SF1yK/xNS
Yk9fJuV0+FZgrBRYj7mQrsDeSMUiIo0KN24uXagBlFB8VgmekOQBQ/Xtuc29rDByQPISjMdu/Xze
hmsSu5FIcx0BwYs62/5apQMHFHUy89UUvp38kfb1iDUjbKu9e6XhUzRioXbde5mL+PZ7cnFtsHC3
JVUW9OcPBjwQC3uJLGfh15+UK/ZHhhpQqx2Arb/M/h5eGxjuNIsxbbyZdKKw0rVeRmHATPF+6XGj
mb04OrCSuhYQlvJh7oMpHAXio7W7i1iKnXHsli8dJp9yTwYAqGQenu96+llqbjDOJVxFVNfV83WL
BWKF704EEkhVOFJ12kFSQCQEfZ4YwJyILAz451KrUCok+yTHxxZFMlPXVwA6hmsREfmJ7owvwim8
SUdZEY45G9CA2KCiALH6fWGlcPOg0RjbKEbC1XBZdhPDO60tx+iCGsB/ctCMSOGapTiQ3/F3N9fW
uvLVgJVXKicJNN7cCfnseBx0ueM1L4Wi/GmrJ1FnH+pnbIag1gArTNd+I3DjpjLuN+hwSkLsfBHO
sJvAF4IejHZKV484OHbAlU1Q/qav/ZA+uxrEdOZbVjlevlym1FCxPCrnIvvauXpd1Qs087DkapvU
tQlZ1Wn574ZBq/oEXHqViGVm+BmIL7yNZ9+mZvIOkZR0g/t9c4pUYNLO2BBeRQbeHryGIohguS0J
OZUtvnaohRVaX/TSzHnUY07boBHFknSJA2D15Afst2Jznp/g9/N7N2wDbmxREtpG4nRgbD6p89IZ
mc5vBfGRnOWsC7SjTLV67SeqaXTnfk8ZFpH9Kd37CiKFPoAIRjcL5s5Xzrp0bWPf5VaHfHy6MiMF
EdEO0gRb6X94Yuqx2ntbhutkfxwQ+DlnU5KIGIWZHxu1cD6g+zrsGp9rOwmumbxmwcqSeC9L1yHr
lqpr8uBW7ozTF4HU46oW31DRwZAJJjWqROaLUSVmCb/Cjy/50kP/V41yHf+Qb1IEvbgVP1AXDlSd
lAlcGo3cpRAutvw+39WmBxvOCJz/Vas0yN5MkS6O9NntZgAaEhXaWxUsWHytBGhUeJ0Kzdc2UABM
6YZx8nXucwz7nzK4xlklsggrw8BB2z1nIiR1sQmYgjZftRfQYkJAZoQaEkUyHxQaqwIWRtS6DBjZ
TzVzcUwZzceWuyID6tDwPC9B0cW5O09pE1EpHapSlRu6UVonhdbHJpd9l5vqoLViRWk4DDKpzqS6
++G5IrvxMawIEAmRCTWc99gtVLEgXg/RRthfewWgkup9vphP/M4iYvSLyZms/JL50a+GjBUrP05v
vI9K6ruE5nDMQ0Jvm5H3unKY1VZPqrLo2rdqxId4iMFjSBKHMYx5P9N8iOT4D3caM0v21RfCUJBC
sUYMSpaAWs0hqHIscg4mcVWXCuQdbE13f9kJGLa4I9VAiXW9EGQcouNW1Trma2C/6HphLkoAoWqX
vGU9thI+029uBMOQ0hQpnwzAGdOGp7CHWIEzADHY9nZm8P5b1mlWfMeTtiyw8+HHfgRX68Q5XGMq
amU6L+i9yQSvlXr2qPZBMKTR0f9xuZi/DRfY4AT43RtvinWqDo4EHwvn//cwgwq1FKGej6+c5yxW
YuaJv8uhafanTqv+umlfiW+GHDa1X9+7G/xT0DSwqwpjOEa20n9lVErM+vme3Bsn78UYi/Yfb7y1
j3sNECvuwueN12qp6uLoB3QEZ7dMfMR/Mo3URLwhFnt5ST2i3/URJBZxQ9+LLr6LpIZjTR+rZnEX
UJzTOcG8Y/6aClObtkAENWOR5sKbvbYjsS2t67i1FPsaer1X3RFHXp5PDI2UN3HymrsZOmmYdkQ/
OTe8wtdge3xzuytQbl0EqQ0ycvcfta4uROHACv4PLz9gio5m7qaelQTbgB0+ZiFCQEowIJPAYw3j
TD0kREmcWQoLNv3uP7lMrJxYZC1lkvAEb9K8A9075f+D0eON3+hZN3+keDefemRChDEIQ+gMpgb+
eVAWuG7+TIVlmukQAvtTHEQ87zb4csR1JucAnsMW4xDRMvxus1VelcAaIxpudwX3LgESYeaLqxyI
lkoS9cEJE79WsSdyng/sMJbDLFWoA+Nk5If6BHckEfA9l9rA0wxVSQC8Pm8qog4OQfuIyIrTaOW+
tPw6ECXiRpIvEAcYmTUopxzqU8h7NwtJ5zM4xuiVESLYCSOD+4NR/YNoFGaFzXnOxnfEJl4BjoNZ
Sxacs/yhVNzCbRm+iPVVVdt7SPkWzIV4ovf3TCVed8XofAd3w1F+LuEaNhZU3t6Qg6KYJV7FxlVP
wCQQYLTexvKSOHF6QizhLnlU5hvQ1mmf82kvaqAgP94nwIQCR+qLelSI9mr9DOpZ95bAsbVQ3zca
94T+xKIMTYdA2qzqeB7VPvZ6tFgbAzxpGlG6YEWxOzfJ92JO9B/xY3GR9jCHd1oC6M12ot7v0UPR
t/z13YOTH2rQH5KB4tzVYDhuZ5beHyaGMFLzHWP/pkWsYkNrBv372vWSId3zqMENKWSlhORijgzi
mIvZj1fx6pIjQqjI4sChNGv2XLE73qx0KdeT0+27el58XLzJydZiAxwp3+6f/0RPu7gSssvtPdKk
iq/1EoQEsyVQtt+R3NpOfdzd4rAkA7rla9Qr1eiaO3PBixzbPY8YBLgO4eJ9WlakAX5iGqXdB9FD
TIfQbq1fMIBH7buOK/nNKQVzM7y1XWmPG/JVPqxPUH9dGpgZdPPfSfKaEk/lnaH9PfE3dddtHWp7
maAgzLjN/Q6kLSqOsRJxh0ve5xFyJUKioQMVmGoqOcK26HOakeBGr0/wazkqywJho1tsse9U2xCS
qpGrNnYXFS75YBv8V2yHgPST+YpLGsmO3kCDNEI8HJtbVeDZ9nY4aMyWl7NAWO/FlPOo6iWCTKgb
PmdDPZsvxp5Z1iC8wyzeX4TTLAtZTWAzNHlIej8SD7CH05C/w5jyATBn2Kkdywl07kIew3svYSHZ
T3dAvxJZXWPcaBvKTZJz7+ng0yprou1Dg7Zq1Yqja0f9RgMrGdDBsdJF9d4EhUEjD/yqs97FlOYb
9APFs7nmYWClxFxAY5gsD7dvzwTJErTuVDAClwcc4iLhwfRl3yS3HMlz3Kuw9G3AkQ0dVRD+w9SI
CIy/+fjTptrDwwRIPx3gAu1qrgvDk68yjWiVNHIix2G7zIn/TqcfQsu+1C8+R4yDYHWwnSyP/aSA
zgl7C7maG3KoeUiG4iJ4T+HFHRreiy7hdKAiJ6liDEgCupFBhzIJajDUsG5U3FO/RLUp/Cwst/BL
orbvAmNazJn71esgz4/Oh90lnpcJX2sZe8vNtjl1+yZA04YopuI2DHJYzyUoDw6PDwh1D2CHfK14
Ghdlbqg0H7EkcQ+W/IsI0TASHgHGJT6Tkr/tHf5LKEnAJ1VrMJt9n7KmiqB1Wx5a3SVdab8yJGb4
lHkqUe8O+8b2gpJ92c9+17i+cYlmgTwNoEKH5ukFcxAsPl5ovzwSfJM5KjILT6Yw4yJVPm9Mk/ED
4bwKdwG2fyozxq1RfVBf9qyiqUcFNz1kcr/ln4B1VWfAiq+JphWipGEvzUvD4rZaVLY8dkKE3UoC
IH45OtSPt8XjQvP59l9FiLiZMrJdtBrzEOOno86w1VK39O3PANJnr3vCVnMQ6JQGVLBkd7MgEx9K
3qmramX8Gnms6ENaokv+ltzZ1R+oWIlY0cOQPXky8PDQawbXqnQ4oD8fg8BvD8zhdLJwvYuuREHp
LL6V+FKam29N+9BmEs/77IhOcqKwUc3f8JujzzEMf22Bv9ZSIDigw//8rooY2gFVFVANf0bPmfH/
gaisw9jqapu12dInKy7dvwRhR3HZq+0tQqvpO2D9K9Qcr5O6Kf0e5m4sxwNWQkspq6tlEd9zfgN4
nHwBiZybA4AtKpkXZR1V1LosmDgki6YY9K7vG27tsLA1koSdOknUJx8HiRoOMvS1fX7CJgKIOAEJ
e4gpyBc3z4n3dRwQYJz7cJrS3afI/J5In+yYZLxhtMIa0xEsY0vN2hZFOGDVQjazJ76YtYLqFRTy
pjtnAKnAK9bz3qj209OvWMtrkH1ggCXPbBseHHqiibzCI7A+nCWqiDLfW7iQDKsmqv/48IeAc4+D
+dprpn7D5f5k+P/K1ueKzowQKhWAwtwwS1WS8xcXtFMDyYF0Gm9wjf/Yk9p+BcQD7JYPID1L5o+0
LdJQjHM/z4sTp2oRQFywJp+IWTFTNmJuMAqdo/ih17zyYS10flr6QiCANt+NiOKG6mmiyCBEurdD
U704IKkGI6sZ8g+90fBfRySi4YO5Bdarf2QDvJtL9R9hzjpLYqCdRSpNTg3sLrTF/SqNDxbmDyEI
aVLc/5LQ3J/mpbEpcLNdtFeUvkz/6SEJua3Kco6r4dhXYe1jYIjcm8dHN0N1LD8k87ZvEB88gDwr
9dHSgMLmwg7LN3CVMX6lYE6g592cO390KomqK4etzn+P/FSMFBSX4IIgiHnlrB+GJw43BCPMfx1l
KL9vvNJY9JvPf6b0Q1PK3Z5wvufITLCZYiZ1F4bU6Nn7uepw2Dbt4/I1atWxzZasISvc1BJteq8E
ZvQjN6GCPaIhfWbt1eRPv/oETebSJRAfVQdn4VvwZgi9WEJFNo+EWqVwIsRt8BkSDss83HsQeCmr
yiyfIMoByJSXtS8PzCLwuUdxIMSX8KhKqI3/t6IicaP75oUzCrtYIBpWNYXNaiyUAunmOcfl4yYU
IpReVmmx0mxHjItAJnfDEFYpz+tz4tMMAfQcS1XEqWq4LCGf+wST/3kGnA0Mugkghfi4GYjzPHXn
sNCLZh3OxDCWQSZcueXrgrhc/zuveqMAByw2zQ6PpvKcbrnUQZeaa0InEghrMteE+VNnXVV3WpyV
wFAMYxUBXLYsBj4YGlsPk0y4OSp9wfSPI8xjjSQTBCteH2837W4kIzUaj1f+zhq8X2UqwAhN2aEG
6xmzWcVJneNOd1Ow2PNgGzmnnRxGmpbdGMDoaTlsYRnKi0ZNjrSC49ICK3Xz6X++oQeXqcVvQ7Q8
QLokHIrijyMmJx11SM646laPM425Z49CSfceNf7GwT9/M+nfRQwRKtMsqBUsMa96JK+6EbHObgKq
An17geZnJRwVR3Hp2F/7evxgTQFIUW8l3GRGOXUBqxKU4mnKHKFOXH5JK+eOq6ybCsql43/nTn0b
7nX4KemRQYOTZB9xO1k84S2lljwqFAEhYP/T78QD70boA2lnbAUf0Y/lMHw8cIV5XbwBkK5R/hKE
3ckA7ZizuouGYYG1We3crJcaDWi9C5KFiK6mq5KLfnPy1lsKGIMc6bGtYJcuKNzej1j4inFNQ8ra
EdqghG/BqKZza4wO5higmr8PP4qNmDxY1VQibrtOSXj+Tf2FtX2OwMToXZBRA6c5zKZCpBHT8Mk6
kzhykpn+1XOFSo6Fzmo9qtlt2Bt8nMyq8Orb6dJHptXavq44AxBEs6B5LgHPSbILU1wNzbw/+Vt9
Ll7Fxf6q2A1iuaAkK9q578c6FjkmWFLSjQV9J7Nx4/D7UKJyhYReNyVpeA/yxLVc2j1qZxzizPf8
TctotHykkyZNHhUDw7hvgUXA/hlA7AEa3fkgnpbtKlJ4ZgDCTqSmCzOA9yHIMawjlhZDA44vqU1Q
DpzHznXVk7mIqX219VvFF5E4ZEncu3itFREhu5fJWpoMaWp+mA/vVV/h2sWNjgnTSS/4aLMfYKQM
HSuS8b5698bH8iRBcTggooaUSTG/d9Vp0SfEGYaZutNhV7O0YWWPGn088PuqHL1egqcAbYtmcrB/
7724srE4j2zW+9zWCYlpXIN7ZhzIwFLwki4JAKBcSFwwlGIV/hIsrkqQQmFKD51TAl3R3rCnVpVR
tnGsAkidpaQvAyVizIJIPHJYMb1nznS3uK8m9xxYvfGb83YdJbK2ISJEjZ9LFUQGT7IDmtA07LJ7
4PEqyioZCYN2dKuf6V+Bpyfds/25GVCEDyyFp6I+sIND6YkPMD+Lp9I8GipDQcu9AkgYX9k8TtEi
9jRV6zLzu7Ui2NfWbfsgJrgLbSXzN0DopVrLZ3j3MMMyfDeyvoRyddNPSI+jYx/kuV1MMz10mrpu
jLHeBQDPMz1WhSKooGiNiSbOtdup3YjqZP3Q60SEMIzgqMTnXFyOUKs7jBKXQoJfWharsgtzDzxE
DHbeihn52NwGhsvIN2gMuM9+pw35lkWZQO3CJKrbbdUnzriZODdEKYkIYOZN9P9u9w4I+5dw0KIN
uQmOk20hUEK1Y3zc4A6eqjOiqm6Y+qQyc/1H1OIqIk1ghHIR+mBP52lmiXeWtiIFB+MsIaGA0tkH
2K3vKkFBp6Lj7LGbTJCVRK7mB/YDZts4uB3/Uvn4x/KV/A9ljBobKklYVs3Vs1z+WTB4LePIOWeF
82r14coN3d/y3gTiDAJWWnx0C3GK8kgXhSmlPkYj5iZAEJuPTUXVnX8CHNaAewIUgBuU/NPRygrp
mbq1cEU84EOpM2lnSxKbeSrTmkmzPLLONvW/VusJzAxGXp4tM3ntgnzQ54OplonEwkaomF+tN1HA
t94YBccySm816l8qoCMD3uSiq+CweJeWMwPIr70etT4cEB5gkvE9WoEjzbrl2g71oFYsz3VLPhtA
OaKqPvcIpNgZpAv7unErCrOnKwmPA62M9klFRALk7jZwndXW3+NA4boN8LTtoaHlVrGiiDyOcdID
Qe0qgw3TYzRs4ycB46cB8UJrKFw6VMp+jO1ZxDJKWoUHgPMvr7KgIINFqsw3Nt4GltNRmVtJ8vLZ
oaqgTbtMyJidUJqeMVG8aNOP+3Klc+RResF8eWbT2RBqomQ2y5L90uIG98Oq5SfD9am2EIMAJcQY
lwn7ZUVL/QxD4h1QZIZVu4Am/3xPvIeZGq+4CB4J8bMKQoZG92WfCvQt5ZwNKXfg6mazwlgf46GC
aq4mu2NCBu5E6iJrDwl2OyhJGVU41UxySoPJFeaXhK6exJluO+YJezBQarTmh5TW7tycVpekfCCq
XHqrVPDboEsVAMUdeZx3a7LSAo1SjkwLLqovPESUZoiri1gcr8rno+RuPSt/WIUNYDSgPVfn5sJ6
Qd60SacSRCgGfz+MpVCcVc8g+uBjVArj2He5vch6lCcbIGsEY+sMPxljSk0yGeqxa909w6uPUguA
u3Gc6qjnnX3Cu7tEa5mHgSmRxhYCfQFhOUzyShcapEbpz07LQGDeb+LD6QpDCSO5ETcQY2uDgqq5
3+zc/V870rKPHEAMEZe2VxKIqEkUfvpVpK17QurMrpSahtT1dxtpzOlbTStMSCdQFAXsMZE9zg3c
YcWte2Wu90Y7tFx64OOo6vp+Cm7stZ2n06Fgn6GsDWJYZ7WF7ni+LhbuxoWee+YaU5u3Wvbz6NZN
B+AcI1C0pGDerxmRXMCkeN0exn1DSs0qq4pItgPMIVcskguP0oqBwbvTLHOik4UOKdvWXa5zg9Dk
U2WKgfAS8Dupgz83dwThgaZ9oyvSEyvM6sn+2F79eTW1EYbRdWwqiXcQ2HZDif+ps0WVrYtiw64p
lmuzV0ZEQcEuLlZO30WHToZoWWzgn1hja8ms4pRWLjzg0KaRrFH1ezcVUPA91q+i7VIUe/VpWgk/
UIdA8AzwC3i0KLzT9IL6+E8VhAbkYsuXlcaHzYZmKISiGisQkRuBFUR4vMWSzREV0vwUG5Db+5hu
E87Xhng1BY1fcpf7OYd+a0XerP4RRYEMekvPa0lt7TBAAzHKd4kA7Y/JenzRS4GipSC92OCZtXi9
7Pq3ZN/m0MjX4zfoSMSIwge5Jh0FwIntewojxn/oQxvOaGrhHHg0BrqlhDQ/IZ0ApLAYmoC4Uz8E
7TcTwe+46Zfc5oj2wBUZKXV+xlRiQK/L1aKnyJzBZrlsLQCGMj+n9o5Kte8Xre1TxA7uxNPEXKxF
Sd2ppGw78hccWokLwOgC90UkZDb8KzXL8wKTBfXPkAF/usgSImVJu+1DuljZC/hT1nKioBGnFWVl
z14z57uTRrvH4H3hV8HsOgmOOEKQUK/q87+T57oXW6jNb2kVWlQ0qESd/BszKuISg8wM+bYCz0+o
s9qICVLp6KeX72kQPsU9nCgz12XqMZ1jO1I7VYG5GmEInNmp06BH+0P6hChPurTIHyZiWU1PiJ7p
s8MuDxlFNJRklqOq+NigPtJoH3ZLfJTp9ycQ3QcJkN5mh0Fz6FVQe3XnfwaTeBx3ktTAy3U+j/XQ
kP/mkZFsiViU79p5URm4ynYC7MpV5RlgMdN7Id7HcoRx7HSo5tRO+xHIwzyKRKpTnnwPcjlNesy7
G3TvRkEvnK0ZIqd3LLNdT+jgTOBorhGYJPP2Y4oWPUbAW2DvU+NP6skbXey4DN15qnOgPpL69HLX
kMr56WVZQoLYyxYFFd8zRc5Pc8+m8DQRwBJxOWQzS8/X6hCZngdigOdwVSFhTNIaxP6dHICaBQ+w
3zhUF1ehKI4UVLqqatz2uM6TtmtzTmGWKnkW1LtAcGAmBIRyNDJtVG8e47zMtjP/yI+80Kfnw49S
rAyILgGtb69CUzmgl6hCen5nOnfIFAaNcplRw7pJsvO9Dm5lzZclZcsf77b0EGfzwwfk+MMK16nR
tKfHWtAzVz7nWDPhH/f/GqGEHR6O/BW8FlBpPkAEvkb04BucKcaRMczFYm4rfpOCstskMVXW5WWW
ewETNTH/3hpgT1G5glHCA7kdNltuU/r+iNuE9o9UXaGkz1bWhch/4/G0y1//UlD13bP89LJe7ai+
YLR6O61yhe08Pu3WimBfX6Ox3x0AMV0lWCg6wz/2CclzTBMr6mTW2v9a9RQyCtSDUxSByBLQe/yE
10cCykpGOfs5Kvom0cxP8/EyWcvk1JS8haWcICRAdcTCRRR73F/JCEXtpQcCS5PxPzInjdhTXIC1
LvEFc4RYocNPbaZImUZ0GCdC1Qp2V/DqurqZoV7P8bj8OAJGrp2CXZ+NZFNqwUwmXsLTkUKICQ3S
94AJYRtBDspUHPXWPa0R6TQ+5aQVZWYnMHB2kWCAbYglsOU8c+NUb8zcUpSXEAGx+aUa3sqobGYB
h8/8F0Hx8sFRT3mDXjk/6OJ72dFdGGoYY0lDwAqpfN1Sfb3s+XY7oRb1ckAmIdrW4g4hEIsBG1+l
YScE1M5c3xyxWTFPgNK510npsgifF6Mg0UVM6xSA1MJ6CZL2+rSiJYI2qd1ECvQVPjk5YggExRTK
ZYRIK/QyARdNRiaP6oLIiCiVvMNc8OBHo3+M0Df3y7e2JrnhlNIHoYdF6XdaSutB2x/IDzBmjgiw
zPminfKfpA7/3YSTZ44QXcwAN15g3ZXQuZffb5OV8jwc04fDd6oysvdwOvJBcdICWPvjPh3/sUfA
jqNP8E6jrqjtI0JjMnOhzUBGwTchKjC6cjRCZkOIbkYyDwRvk+xcU25XTsumt7mMnh0719T40lyA
mB5drlmsl/4NRzKIQXF/5TjB6UYiHmGeVIZsKiD3W/g1XwwdXr8FNjpmTsV0LC8OVSxdRkvW/J+k
/x16aMZTmnp0qbwyOZ8YBnq33HUlfA+Dp/IZP7H4s0PPIeHEIL4+HxQsXmN9RlVpvgKLBhJUuGWC
YisV6NGPZQX3f4/dl+uyY1VB+N07gkdgYCeqlGsUizhkTGRf/vY/6IZHaqY9msIlKe/H3Wej6/KZ
RGXvuA9FRw0C6cnH09m/WlyplmeGscwpjAJg8GzJtMpKJIBzwHgSxqPs8YQp7LxYGjOWoQ6BsOod
Z0SWjpBmWymVk8Vcdf/jP8FCyIAj6YqQ5bP9imjgZIUspR/Iz4fublvLuC4AmHPzGTCDsEhuG7Io
aKaEByS+oKDCH2ifdFUIXHQp/nykkwVxerQOIfV3dwog3oarXPWYcPkm7Zq5aov+01HC/l/mSGJk
O8eaA0OlowhZBZlnvOzZXlICuyrGZrIA/VCEODKsAV/0LKT2HiDmmceGdXCWcCEoVc+RtKEQGevX
4KBdCh3II9sSpx1DLXrXTMXSPV5jujajGW2Cio/0apJAxh3ZQXKA+gfruIGgHLYEM51u4mmkRQ8z
3SzCi3zW2sZyU3PelXqNHDDpNus2hlPCUqmhtN3rLoK3hB1/Ko5gpMeqW+rRveS1zQ2YYOz7E3NN
s/D06C2dmRjjL82fC36cpo1unvSqBlH3I2IPXCzZnK5btvNBGFjYWvgbcXYHFFi2mrF7XfH9lIFH
5qG1MDhPkupyoxQSYnAncUa+6QA7A5sQfDpcNdJ0jVIhm1TdX+nJroxE/esDz2BB2NRPuOgSHpnt
K8XhEqsNSavdIVgw6Cjdx0l5p45QR3uUtjlYt2Bg6PsDab2dckb8uKovYJY50uSQ/rcji7rMHaXq
lkWppQxC1obHPHHisxaYOwhIi2n97Rf73KAJ4nXv5s8HzWbUnSWcJTnQskWlbYQEbxGmE7c9gYwz
+oGynNuhGy10MiJk6SxCVcSFXogZc71Bf4aZrqTYV9Tb3jybSpOgbxxmdHekNwJ1NECXwkBVdSRv
DH64Wcs8MgSaCAvbxJPmmvtGCSr3VxnPWBkPy4Ya4VFdcKnKKWBoid5tlk2BsgimWorW7K1c+YB1
DpYgolIZRH6e7YHWxeYxvMqNMD5X33+suG3dLeAmW8gBlaNNDiCQjLmN9t/fKefGIaZMqUwpownV
tKwRMT11ZNJuXL/dKUgqYrZvaG4TW1VYIwzX4ZwwwlEm5EQPK9T2Q56y5NJZdnYTiSq+nNj0WPj+
WTb2SppDISQ7jqITs0ddvKFfX/MZ552W0jGU4NqlliJ/gXZLMFahNvIhDIKCOtN8LBAgoNxNacV9
KaJbWFYFoct37BnOR2QrNw4fkIqqj4R6r83rb8x1aYXKkrOVSBAMFCTD/3+ULNbwmYXe7zd0jJot
ZQqV/i0tu5dFvj3f8tNnKJzgDWBnFavxWkcKjDhyjb6Am4sK6f0vd+/EE3ItR6xoHvf7tvFytbat
cYRRlf+EL2qQC3GaIUFPgxcR1RkGRQBdtTlYbQa848MD7AMx4Vqgw2haLSUTwi4PCeBSqYOdNF84
o+Tz7dpgk0Xyrhtsp7cantd7bZ5MvwnNq5O1ITF33J3hbMNdocDFqxLF8jGG6DUjzh1fPBQdvpGS
7vK1uk+/tC4KByvDL85spPWY/iJw/ik//V44zjV6Re3lrwjJvtuZre19u1UDwnL95AvOzsAWLCWC
YkomkilGYbuuyZ7uCDSBUfTTWPx9mR0HQnAAunVAyg9XBEIPkg/HA6A0hSJIaHTU1Lnx3yL+Jqqp
8CtNtX46s4q4QRlkMPlQ7GH5Hqx4Zfh7HUuts4NRTCLDKB36ogFB/rv6KJ6j4CApfEyQ6fZxQEcU
5H3NM3CHKCbSAKHggVGvM6Ckuzq5LfrSIuNnZcE4a04Lv0Ol+H9rPXRNeA2aUAqywAUZyITRcX6P
wgJ6OKT/8dc8e+WyMl4HXibOy+YRetJ/l1Idu7afsFtyBc1Lv/FVmsfbvx+RLwWqsXCYlDGUrsZd
RufA/Yrjgbuygn46jbyJAsz6Ng8pXrwPfcRl/d12BBnM0tO0VMrEsQjWHxowWlavIx4MI+dglQ8+
ip62sjJcn+hiLQhhotoINOz+AaNZR+iduw4Amz6GhLWde3+RRtIql6J6NOhp8P1tkXuSznr+NmZy
Mg2/xr3PMsumxE3oVgfWJBaJJe8qDFTRBUQabDGmAchUW78f15fgzxjZ5V4vK29zL3fViZeBVvdK
JDlwKNMK4D2+/T7RPHfRg4y2jHuUpAc8O4KYSXYVvQJo/gzfTkUGA3ugTY3FdmxjNmlQyPM0e8ed
FGzISgG6rN4158IUKLKqcbFDbK7W3GBG5Ui+3Zqyn+HFuCjfn7VMlzOduXeIPazee7tqlygReNWZ
Rcj6MvnPl93gGqDHDkOLqjOGR0jX+mgi/FxE/gug4cr9zaPZbnB/kjSlsSCCufEaktd+rQCbhgX5
8FN/n8FG9qLMcXcQBE/m38/PN21RnwXxT6NyHM3QYnJdx2uIrd9Lg6g1t/fraR57zEas6xMRNlan
Eren2VAFxXzM+GS+y2Hd3R2egsSV010qPJinRt8+BS+rjideWnBhfWYAe8Va419sHxndd4rF+31f
YGW+yDSaG2wZA2deSLnQ5qvxtPA5UPOKwpPiBYEflV4I+F16vZTd7rh92RrXNXrlsyW0IMgHEyWz
9vXWHcJaD+BjX+kAY0SGpbBTWwMZRKNCigGaveiGqix6OeEmBby8GO3ToNQC6H7iShZq2Du13QbQ
fGvGekodXJf+HPqBP9PE33iVoTyEFRwbr3aggevcPCKTSVCcNq59hzCShRrbKIre0I7wKv8iDhFH
DgKocSwFlutylQ+4BO+PkQv6y1bzq1AeTCbqWUpNcSC+z/Nppfo8o0Ile/AW2BbCyAXKpWYbIJp+
aIll0/SclJlCu2DMzLBiAoY+nhHJZVLPNkHLuuwPxHWxP9BZd6IJQ9da1WvM27/JjUipdzzw8MDN
+bf+CUyioE4ILdJPaz0oakGgx55z7ruefua1rxBpvazbs7C+6Gp3VHOkYBtq5g9eEf7YCrrng+SH
FnWXkix3Fx6BHgMoXxnoNDXmgmzFHkTHywtM4G+nwM45BiWRy3v32T6ogPBKd0VRlUFnp3rMQH+N
j1h9IKuJzXq7zcHsXKIy4aPDs70mzAjGV4KRbkwZjzweQLl6QxZFzM+18A+Og/RohAlUX4qVyHvs
74VIZpzstQwoaMZRzjtqFDb8SLA1wYLi/0jRjh5FzEnHv00kpXM5m6qnVAwarQMuzMbq7Nkig3VA
01Qp1UBuBTOIsDy2VccmdXbdtW2Uq3PJxWTF1f03UwvAvrBAA8x3e5zySKf+zHOwXFduVM7tc3gE
UXQJANx6d80iWV+Jz1qsxxZ9KUXL3zj6yy+VebMwKKJ4uWBSs5DbcB1r2Qkrvx+5Ykoyg99W+74r
il7ARYIjXKPurAaHDK+VrxB/RHgaED3+HW/J2TlzY6aRxmDfIFiC+ibz9d32QGWbhcGIOEKvMSxP
PtjW6KxuMSRq/AJRWEww14c61q8zIbAWQrAIygyX5YHBpf2nuJ1xfrnYYspdceaydlk5QdpA1tVa
F58woXxo8WNzSsLiBGIynEPyo2T0/SO1sW9UsLeOV7JBY0ZZ/985e40HVHJtwL443844GM5jn3Fs
jV95n/tAntodsOHDhziQzDp7tdhzRlueUzRmEwCvZlp2rSVkIAxjUE651zBiIlSSEsKiCOEIYIl0
kZDaNr8yFNLF+5XyVSVmgZZ2IuY62kun2DzFbV+jutmzJkmZSVhcFi70zV1vHpm0Kd04ev7cOwOd
/NOzne5Hzob83cO5qAoO4mi5nC3mJ9C+4ASDNBlBJna9qIpdUHSpMtWDaoedvZD0NWLWUebWf9zh
EsIxVzRj9ew0YKZiaFBH7U9vcyG6KR3bn6ALgDve5u8sNO2iWEAYLxkQJV3jt8CMNegAsm7XVwta
osIEO13rDUtrBexc2sooAE2wcqOlKiuUZnX3aYEXKDKSS/VF5RWZYkocT5ezZ9lg7TnuOvgSqyYm
A2j8I3Ns3en3N77qD7oUXw8F4/5GBjm6DEQXtnOZV4FZ6aGbxeRP4pA5Tz4rcWwIiq8dgMKchWXe
6j6Eq/SYCVcQtBU7iXSM54eTVdZNcXXYApbUcdugy9gLT1zWwZpplxJwFOs2hzHjIt5TPQZ9HBmC
C46quIHNztMfHBSBIBBEqoOnmR6o+RZcMp1P4FxFdSMG2hk1MUaLIyXxb7UgPU9h3h742qiCWeR/
et10zCwnEeZPIOCkdORJPnSQj86DJ+JDkw7I31eajWG6VcJEpY8elKSwbqhatQmftmdJGZ6T/Y2t
kmMYY3tVG8i42gJgv+yZy2uxjxCpo48bVrCGxMKTQHcQoGFgCJzl//08aw2oMvFtDyLgRWuRki6I
yPDfItonXzJo+qV+VXaFZRAoo37ffQ+EHEaUC4a4VR5gpK0ev9ClNLVLHHGp4TdZRmUuW7LdU2to
y5Jf7hTvL4A0JBv/64de5FY3PH/iUlBCbb7fCLG6Yi0Xj3w1SiBU0bKR0FmZDDDTQhIGoEnLNNm8
P8102XwzCMjPfHoojKhzwuBCf2iVKpGrlxSOJQOM1zhrMdXoDAyhgjLWZq07KQQQwpQ2tzR4Lz/D
1oBhr17e8GAKzWaDYo+YCbjIdKNZgLuVSiNJaBICDsWZwwT1L4Pyp8KRbOfilgX/a/2nxwTuIo+y
OXshYdnC645r5hXzke+HtC6s+Tbwr3xJQug7KfDW1LfBIfhvPmXDKeoTpaI0gQ11FbS6TgYvnAHZ
0N8DWD7mSyu/F391h17hP9tJp+fh2C4QdXeyGi5+30Eqt4GmhzCaorEMR87fva4RVZ6PCfhs6+st
Evw7pxrkTcxspajbHl22s57B5JeK8xZWj6whl4rQ++D4gE1UrhXipjKyuANEOXY5k7nlm6H6QnBQ
0sDhox5Gm+3WhxO03NVLGUJGOZ9b4Vfnzspty4cr+Dl27N5yKjqmanbr/hT8A0ea+ps90peLXFCB
yj9pFl56TJ/Ice/jYPyLLALC+KR9pHeo8voRz3A+NoT3JTcs2eEC+E+tDXhl4N9eRXxj9DdHsQvS
LBpGujAoQikrgII1om8SFGaBh3o4Y50uSkb5w41QRpGg23qKtjiA0GbRtRlXvMbks3DZGy/aBEYt
2VuihZlXO6uipUivciaxpoN73sTPZWCQSEFUQkffXc6ZOFAcaB+Ra49Paic+0pJIvpyZAEg5Dhkq
Lrfof71pQFLeUm2h/R8R16SqibUw9NFc50yw3Zni4ym0q4lc2kLbZJPRjuLU/58tAY6uL1YG4G7j
WQR2+8xkXSUMKGH6UTSDd5KsFd0T8rSi0qbgY+jEKfzHAep0p9tPHh4RzYKAkPszIBuyIHxuPd9S
9Gcfh2kHg7oqkm3OrnFf6BnyLwEYDQr8XtMUimym7PB81aldy1Gd7zVMbq4xaTB0smy0EZC4HBeE
LRp4yKL5pWirNMBsHHOBjQpnuqntkGzF37jK/8qsR6O/gcJP12Om/Sv4+UPzhtdyb4zvxDOqLNtw
SCm9HPRQmNgw98BHryhmbaqp8fQmCeFqdu0Nx86MpfRsPRwdHBOX8LIbINJjfnZcHGGUCI3HG+Z9
gsWwtee6Ite5xJ4BuU+coKxHEql4I9WdaeWL9AN4jwJVEpP+UP4hHh0pffq4oPA4eDvQ5qozNv3g
iN116D/CZv47e5d0ipKa337qM9/crzUW6lLGyO2gilXZMgSmthx/TlLOc/6Kyc4M4igAmA1WB9kQ
ZJJRcyT+ybKWM6/C7DDSZN3ytCjyb1bp3qjthmXM3JW0r6cqIKBgOGNxzMu5/lcd55asls6VDO7L
FQKIG5ePFztN4XnxY0AkW5YlXKwr582VdHHptU5c7pQAyhhKQvqXJGVVf59sI9MgGZ9os5T7P2Rh
dxx9sxRqbj0OAKduBbY9K+hOP+sWAsT2zjELgQuLzesXgY0OniZrKO9YWfMRCLTpI1aXOWqsbV3V
BZkFvYm3LIoh8debyldm7nx/0+FhSI90qZ8nyUNzwBbNpIHc7DSr9dfwBjjvPsEgDXqy+xrBKsem
NuZVYxW5IMfwAmG72oZdP/w/MyxgS4CcomhnpH9utjnauCUYshTV8agiAK1sbODtqFZhPQ0hG7jG
hl1bo9JgiC5+OX8B/40HMNRreQy7CeNHLFmnNTsUnlLO1F6OzA16lWVOhExRW/pmdnnnn2EEbjv1
2xO5GaAK6+9Fs2zkMx7fN0Pc3t1P5Bj/AWfleJ05JU8qmb4b6tIuHudkyk6aQQ68Mmovw7YeS74B
5nzLWVdSwrhw1CeaRHdvpDTc6CTzTVHmWlBh8kVEBpOZYatVXgBUm6OfL9Z/xYzVGlaSZKQnMChu
/GmvnWOeGiKYPqFrI1z4U+5bSWU9w8lsuLMor15DtrkX5hKmacpiIOu8NfDA3FWsRH3zCYlUFBTS
AmidxtqhqVvWnPM4FtdQrl9yWKd8riF9K3rlxtT1LViazZdJmGzuHa9Ueekn0QfNK6tjVUEUWqk+
g2ZpLkPJYP/eAU9RaeNTbP7u7msNoBleysiSUMLXxyorqhDobH8+8GbaONh40+lArD7TrMmXi7LQ
0gI7W2sx963SbLKZAwHKyDlNLzCRu5adwXltoOno3DueJncTKMvGm1eB3aTn1BNlrE1qzFsq4gj6
JQFANgw0m7tiUoRqXLbQfxIstv+UQuV69gMCr3/Xc59vf7z7/3+6/ET46zeYQ2VYeNR/++vvV0/+
ZkT6UbXoRXqEx32jhKU5Qy/I2RK+b0yyGrC1Nb/wYnFHYD1z558whbUGHl/VXU4YAHI/ZlcN8WvX
qpzQ5ibxiyvHV7N/zH/4ifRRxDcRT2cF9I1QpYrwUlikvf5HBGR67rXvv3M0ybCQ3PmXiFoah+Xs
XKjqXJG4JaFZ0gW+QsN/QQgjU2NS4k5JCd8bN6Qub5TJKL1WTmP+Z582QOGsskGfxpQdEbcJ0Fjp
9hlCoMDFNWgwaZG0fkpxVNdMt7eS+OIPijh+8D9cuQEUIyONtcHzihbN7bmYvauOhRMG5fzOq9mr
kROc43J/HFStjq3MegNv4hJmgJ1dC6tP21bXG5Jk8vOZL6M61fiQSLYHQrfLdLe4p6hBrCD8Oehj
B+rH6tc8O+hGe3yBGTEG7lTmy0SjktOH1c7GayYvOkcCqi7T71LDwGfM0XwUxebKAx0ZXlKdOSqU
HfrGrBfOXAq+y+wIgaNKvFXLAhxuLV522jwH9RSY4QmLLn5eTLPHWCZ9UdAqK0Z9jcXOOa1ZMvJV
RTAFzrTmcQbXZ8JWM2DUdRa6g31F1LyJ1/2wUfXpU9BSZkWw+m3Ao28M5d5hVSKLAF+hstGUC6AH
o5DSf+8rExloAJR7gQn6tdhIy/gz/yRKaAddwB5c91EvqcH6rPWusN/8QdCzxUnamsQmXM/r4+pt
bgl+Lhs+XIK2ToBQvtRMfD/40vkSkF97JLmcqu3lrbi6VGvKaX+U8BV1Ha1KIiDnH439TCS5BE8H
jXeDTEvgzeoFVRKW+qL63En13dFD08F3DUp9IRhQLmrGZZVYcURED+x59U7VTYnW96vx5QkS1TMa
r7LHzRXG3MeT0AJpKqjq7o6M8eAfm0CRwUBuKOI46C3SjbbPiaqPiHVVrxMHB1w4ogHGZcc9Vv+N
n1j2dUs+Mp64D/BeGCY1r49RJ6ifpR1FPpVYSnM3r18mnSmxu655qhhdQ+RPOlC75qSuwq6BR+ZV
7dilfoQQVQqJXJsv+ylmf8y7H5GPZi7M5nvXYAar2lfYuaxMAZrhDaNfIIl911Lm95I6HLn8tzRP
zTXfqugoCYyNeABJVuQ08oz/C68UrVWlZBCkeaLd/yX4dlBaFPGNc7GEJf9Zf4Kam5ZblIsFvxEQ
HH4jp5DuuYY5d3k6ZyDDPMGeZWMPHXbMVkgAroFS57nF9LCcfVu2Cbk0wmyzo5NisR73Lsoz6owq
h5oTnqmQOQ++ciH/2D6ygo+TenVPBc3X5bI6DK+R4xSZOKXiJ9M48WGdKjUOCDXjlr6Ed6qGbDkq
Pil2BjOTVdzEVaK12vJ+A8rqQe6UMDHT86Y8MqgEaepQi8JhbLPiLPCv54K4It31YwXY6gLpoCVT
ZewA1HLQy7ZERHh3znJq4qamg+pes64oxwO4I7pbYaO2mLk23B4thAYytYw/i2qazDO5kSnCX2Ge
F9BtVSBrsggyV+HR7rcRT7uTY950IGnaprFKOGtg4dG11oitdHsN2uGfTl9ubehGQbkGp0g5Pnvf
gONbJstDAfGqT8quj7Ov93Ljz2d3P0OSw6mmbLu3GQS6MnFTi6dtkeV5HS+Ung5X1EjmeKNwrBia
UF5Bd27/Dm0QZ5euIi/fKP2JzRiJ/VcfwmKpidSxYKOXdHaW5887TAOpR11heXFvk2p9PesrgK42
JwgiKdxr05wLeodgJX2OCjwFw0tX2/q1Df+o7VTDHdm0dWpxOyIRi5Xg/83/ow7GS5wjjxrk/K7L
DmPzBnt+KnP4YueXGXon09oVc0CpI7Sae1GqkcQo7q95IAPx+9y4KSBD419XOhLWBSkVdx3Fpam5
6jHguEARq9BC01JAfpmOJ4vQgznyWUDXywi3L5XRyHdnADGi2reVZJi8EyBgjjva61ml5nGkmpnD
Tt7EohNmLBMHnz4Qh0c1FYEKRT5EF6ni7qZ7/A8hhCz71pAMPd4CdjxPWpG1FPDyNUn/6WbxSkMB
quNck9ZMLk128rD0ndR2VLTwesvwAMSkPh56WYT3MEdmJumXOaasIHTYVHdY0TF/lmJYf9MmPgtn
d41Tjujker9zB446x7Ryfvo5kMaIMEd3IwD3TscX0VSp1S/KNGurozCGJR7ef9BRisBTh0k1Uzwi
7onG6Q3I0+KetRbRNqte9936ggPISlvvRMIut6oh057CizyFEQTy//kqaWMcsTmhinjcdzWA1ejw
H09BdS6ILYoPrzheSQN+08wf/kNGlZi3tIMYULKU+Z4MHXXAB1KVC7gHCrs5MI9e11IBQMzokUZk
+Qjt+PKOwNW9WT/N6AEuhZv2ikS6axv87zGihU4jmazF3W6LjKeJFlKdOlTLaKXHEFujqkBsh4gm
nwwTRmcN0241gdu8TflgcbLklApEUtYSRoAxfb/NPslOfFcje4qY1g/Jpy58glwrkCHGoPMg4QzJ
czYo1Q5Zad4C8vooEzfsBOwdokFS7vSeDJWtjMgJp2cYoqWRiVXs5bagudFGyRSq48OIxP6/bosn
hBLKKAnMFEX6KnBiqRc37u0SIkAzvfIa2d3DkfCJN3awqJJOk249+hgQIEDzY9QAJGSNc7B0i7mD
LsxbELL1n2aZZWncWro2ktA5ZE3O02YQQ0NBjnPN/wfiWvyWrF3PWPZvy5Z3cIidJmY6wNOKIbun
qJTqQZT6XX7POUCe286fg9e/HLXSxOhAkKoOqOmgFAiCBEipuLhNAgEmbegZyoUWE4zPewzRxdrH
WD9pgEraGwjAQDYppiLfwAeRG01yZ2ElB4vqtBz4To+gu4UYB+J0gWgu3fR5CRJW4PLEPEZZNs/a
+13ZqWrSTym+YgsQUcrCA9nJGFTZ8p1B4m3D3HCAoKUCxu1fLYDONmwLpwtjiP5vXWaHJBWX/rXH
bPj4V7HDuoDoGJAqNnomI8EAdZEoQS0tbN2AVUvririawQqMvpsP7MSCZF/9IRpgACr2yoPeRnev
JK25dG9NuTiTq9B6NNMkJfxR0GMQZ3Ragd4Ex3iUdH/mdUhznrEkwD62Ak5ciNMXwmXEFpVc3FGi
C1qGU5bI1zlk5CdiyIbWeUrbwt+Z6o+bdEuDOEE9yNt/zwaMveEKkUvi+GW7fCqBw9yR1YI19Yvc
YIyTxAYP3Wlhcr9PqATiVZ+hacF7ElH8RB43qPw1LE7IDqZtswGFCmBebB1bKrSRQcKLrT+adCc4
7pYk1ZgT79xgxpstImY/KpcIBDIbUiNQOyFMlx7utbtv/VYzz+npy5OQ5gD8N8GjP0SYeZ48qt/x
Z6mlcLO1/ghQO2Avsp3jsvKipv+rY3WtdB4dlUDItsMMTN/Ny/OqzjPkMQGOW6vdUsE2TEIyBucv
ZgHo40Ed2RQVa1ubTBfoOYFWnsD1sbhgSsKGl7xtml+F/1yEU7gHd39I8BVNA8dBNu077dD75LWz
vu4DGysQSLRnl93gGPLxWpOaP8UVJmVMj/SEFdH/UtO9AGXlhkqkteWHXIFhydZsXizRhA5eLdqt
e8FGDpv/H2baqbhIDtI4eqCAdejKaNvhHI25kpT34OvfQYboE3Ft7EFFOlRQCzYJ2q5sh3ZHeDOX
1/3K7ryw/s20szg5ERCEzJ2L0WS0Qec+uv4oPLAXRT4qmeLVPlScud7U2uEewf8cRcL6+OA0oPZT
SLjmagXaZ2XGpecziEiUqZXmhqDrvYml9tZYRG0o81DYA5AKZat52JxP7zWxvjanW7WhhdaHr0wV
buZF4Mkq/LabRuRnr9ORky1gDYdkh2/cKBGZTrmylL+E62zZCT+yGso0T6+429gXLnP6GxF+fGju
gdAhcTuOcfhk6dyEgrvbvp5RLrw6ckCT+9F6iWcwd0Rd3ULpVt/nATak1qv1z10K/NNxlBqb9vGd
+WR4+twIFgEqVP5pkMMYlPvJeJeG8S9JKTMCw+gq8TY+Wrvamo19Kljw/waYVm3Z2FS1G015YW55
H+uzFAmgz1hIEYK5GFvrvq0wRTzzjoxdalHh39SaHIpkzcobZJLeCRliH9Md79n14jcDIHie0hRM
psRo6Nv7bCgR7oMMTQk+XoiwzZmgnbOi/8xUVOAiGC8lo2h6ofzutHrkFZeGTlLOB7wypXBsJyaX
/P7Zo/hZe19DL90dTK4D1qlHmyWSQLdDYdRebq8XA4YWWD1lzEaon8p+M7mBlpnDIMlHCxl2sdPT
fRoKW2zLkD1LiUH4myI3QQet/SA8Uo0RNv/urTczGEkjVcmRE447mxj/sWeL8TxEmoFClU75YrnW
ucAW9lMmorZK5eXn97Q+1OzsPL5t4ncv97MGi/Vfz74465oPwAccaU5vV5SRLwAFAuKV0TaAirLf
WPTlflu9bBAW5Kfk03/FQT8m+D5V0gvFm7NYUh+NQD02/Mk+2C+BvTBuOvO1eEx5tY1BMBbGnp14
Iozzlg+GyYDX1HOvdlbdFEgo5zGxfcAtZ0p92LnoPzN5P65LMxcFMCA5T4kwthJN1Jd4mS2Slsa/
7wDqZ4dgW/mhOicbXZVaI6EM8j8lPtKwdg20+xGAFdTkcNJSCm4LD8WL0SMPIYQCsHh1hthxlyjC
p0GUGDcMPmrfWwvHvmSpNkX2pwj135YRvQepFXtIATr1DYHELwM7q0xO4yU4CqKlEOKTbvbmMiNr
pytLzLAzBp74WlxlTJtuHknBbUGhO2k9CP7ZRQQPBTNyMsPjOHDLg0adihiCaR/sgyfttwgULAl9
hCv9EhOoUlHTyYO3OBBWGLvCUxIdVfkSPR8TVwsgBmYT75tNBmoHlJmdU9SyN9t5u1iiDqa9pJcz
NUtePfR8mUJijM0Q/oTU6AOIqWIO2Ddx6zVweAeDIKNcMjaUyZ7GpjG/t30YPBQO/d2GrhpzllmG
DKKQALFm4JbA1qPJTlMoJ189LFrWCoRVu3i2WK1yOkTlgwatC3xmR8Wc+pAfmyNeDp8JGe55kZp1
lkE4oP4ChNcMb58mz83Lsgc5MVQEiI2aI6nYQZdT5P3AyYcMAykeh4zeopC9LIMLTQ6gUf/MPFrr
ADJdvzQjvlrtCN1oV6puLsC9DrkUgKfdYcgo+YLjUfMgOGqSckjwHCwFcJvmuoAjafAHiBFgekGY
YLFb7uJ/WaKeAEQTSTKgIGmV3uQT2W6SgfKVCBt+KSe2uc4X1Sn1Ifv7+GiM0JabwwbabJXnF+Gb
98Nry6+EikcAisszu9BHG53x2VV/d/dTbiSuazljYS2Hw7GWo5Hnvz0uFZiGRJED2ix7u5fl3m4U
NM58/VAHPJE9Y0hXUNv1vyi7MZMZQl6WF4ktW59XqT4Bln3X+TeT7Kpr16NjDgLbTHtaBr+HwSdN
uxGoDotuv9HzllQNW3hvSOt2oNfJgoLxpumhGEhEnJmHjSjmveOwsQ3wWToLTdEE+/lvvKHbr3z+
4RQ8D7sZ21cc9ykjPDzZpzKbL5ywbttcI+KAnpkShOf0m2cs8KjE6dY4MZ0A7NI8Sq8O/v/dJ/rQ
spTQjv5nOdnhGTTCVW5HIHhaxZcCPpJkdwSt4Qdjdiz5JUYCzSekKNnT74iH+YK15RC1qG9qIAr+
RSmFfgK6O1iLMJgxase2xbZMD8Cu5hVBJholFQFoyJvzbk6Dc94aiPrRZfommzoeACyu2zTAgZMg
uzqeTvfL2gTcBftBiEzjviz2NSgMZadapKgOmHgBRI0d6i3gZr1hbl5dflA8Hed04Skqa8ppGC+7
5UCZWOBk7SAT4GUUh+z6J0UO3lmI8CLf8tjHutWfsgtR/Qu9x4I5fFN9sitW6YIr8PRSsn9C9dxy
vIva4Ztct1VOvgxZY+qFvAtinrcvzIU8D9B3p9JLUCvmTTj7bfoXf41h9vpEkHqF42/wqwToRpgl
Breem0WGxStARYYNHKCEcoA0Y4nT1Px38f+JJPDEIRKwuReGiffJHH7BpkJiFm0iJ35yU8c4c5bb
c1yIHFtkAJk24aXqcwHYUIopvs3LjjPbxmj7XTS7OillErYJ7A2wdxpv3t2vewiR/tKFJwgy/zMA
RyX98VjQ+V/c8LPf81S5ZLgzEJ0fOQeEVhCxoAB93IwxxzCyzbBgOPQmPokY9azSW8FmRfq6/d0L
CEIhsAPXghlLxiGkS7BZcDKakJGL2rMHnN2Ae4iaxDDomQa5TLou7kbJXC/Zv5EVgK1YHV0sm7jT
tgLrXD9vu9gvwTOoHI+rwrf/dwp1ggpgtXVtgWd5mFm+OA/NhretZ6HrrX53bgxsLq4pKsX7n/eM
ciO1U8KdGf35PxKVPPtqOF4jWavbU4jrCjQXwvsIoV4cWtUpTEsNz4kmd2RKJ5JV4v4N+unJflJP
xpO8eaxN6IMMVzZvx+E4Qe3Cbf9P9bLdTnnYriGlNy5gl4HuYfO+6uDChz/RU/TTSnpJhE5JX3fg
Mrl1VHlTnKQyueg93fwyYEntz2AYXtm2ZKtIiJF7UZCOTi6Vy7PaodqsG0emIGdcd4d/jJkh9Z5U
5ILEb7ab5i01BGppPGA9d84SyMSqDhW+KEOIeEgue5CW6Zy8kqdBfnJu9o+0qS6reuhCeCZR9yEW
PfPR/kVoDvvT3qi4iFqWrob+xcHo/kwrhbbt7D9A9/4JlJmcyrtvs6oFGgs9jpWMeKN14lUXHrAs
iBwp0rwlqPexchDF+2R5cqjiqThQ+/7S7kiVwzO05a1DZ0CXu0SgDBxEUML1y44jxll6ht7kDbk1
JGcP8Y3/ciYvypuM0VWdBeREbQAKnmfN07EcFkdv4HZBx1DfOeoow8X2sXpZdbRbuwy2/wNm8FgV
EUEvS9VpVeodngtJSPtVLEIasGHe7WYZe59sYS8WMNR8ujZDqHWzr2mbOT57Mp8txMTtenR5jCqh
L+Sjsgb1UQgHbFHmKpCNQ8cRTg/z3jWDAVvI+CuzlymX+GMognGWEsOZBFSFDmjVGhRO+cgDXNDk
ooRkPtLDPnG8DKLc09pEnqwIyPmpPkEejz7TUF/l+yK/IKcD5BrBoexONmEniXqE0doJs6NIV35t
VlLuUgQnLcgODBZE17OyZPcbWOkf+/fLCnm7xFZep53FWyzqYz5YwKQwPh7sTUW2jIpNBGNJsTYV
P9CV+fZ/01WclR8U6brFmLg/2FwKv4CT2RUX6czlcgSYzzpMtGYZpd1mGWUxP69vxRVLU/KtcquR
Am2mAK824fKJQSh9ZiaBLMhgH8dVNyKaGiy3QtSQNS+ZpAj82H4xd/eNQwybUSFvCoacTngDb3t7
ObOs8+GqdkHABRc5biQG3VR33IpY1id84hY7HjsySNN3r8OF9WfLEDk3xNeV/bcAbB7S1A5QGZBy
DYmBOt8IfZjKPPHXpOLWhPPdLzhdikRJO06S61fhLEgHlqwqYEnxn6MddqKa3j6TxAj1THXSIfxT
ehm/nVUPDyylm5p5DYZO5xOpkv0ugCkZGxy/oAoeVi7ZDsHrRU8dpziGdaW6ExniwDQssQbyaq9c
226kH7b+Em0S7tuBKa0zLRB5GWMUsuFGJBBt41gLFBy1BfFqkGKUSguHpJmQPXOU0zziJLsddEig
AX8oyiQiHApQ+Jv+t5/BqCvqeLF48kQXFs94uW4fDfMS9yXaN/nydAHYAnJ9Njyc5NnRfaIDmTyj
PcYGIGaipizhALIDUhdaYqs3Kw7kT/Dq9j9m6gxvgiW5/1r1LuDOHbxcjGaDvcNyEKKMgMMNOp9k
Pu1qa/+Kz+lf0YdL43eXLccJDRcVs6TJWnfXGwGlXQ1kH9dsawlX7922uTBwW+Ek8dpMRrwUNZRB
3wxzypFO2EFrCBuu6/iLp3n1ddM0ZDwWk8OUFowRglWzl03htV/QX+YqWlBXSNd3urfwlqWvqNvj
UYbxYtsSoIauiQtqbAXqfF1SMHqyDgv8SSmiEitnPW5Cr4ephMJNdmg2cXKWVa8qMsvOsXRWcUWG
d2uQ+5Y9YJ2y5jUIJ5ZnElGda4BY3MSwEBMef7QfGpDMd5iwGkqyeezJfKBfiUas0kAQ39Kqr0/m
1r9Hksf3/BPlxEs9lOMm1MRgzm2O9ysTOb1CEtherfqgkZc+J3X/PwHlCYxrJ/s41zSMQnSPzAbP
+TsI19Oga7N7JmmUnb1I5Whzr4jlt+d4aA66eNHffYUKMEbhncnGCE3OtpAolm8mjSmAyRNOLMhV
QiBsZRQVMKNF8UiWUHbyzUlJufSvbl3fsU/aUO/u2Egv6ReK/VjAume/qa+0Wrkg9RU3v9C3IJqY
mLOly837iP52YbTJciHhmQzY4YmLkmJzhCVcW0Hz5H/KWFzDDQvdur/5mjaRTuSMnU+DClGgJfv7
K+w5nN9aJWm+/lLtvUk5ATfDVrAlpZoyzLxpJjAHMMvKpnm28suLrdWoXqxnMJTpudPKx/ZKUxYb
eu+/QzK3e0LlxnPWxKFJFUiqZC/hO1W4kpHemsgD6isgeD4tEnWo8xfiG/OY6CtFOPZHjR79qQe2
g9krAyHifltaisg8bykSMl3OGG0lKNR7d/2Ww7UwA/Uo9D9zlJWa+Q35l31hzEo+0UYlHSRi4eM+
QMsK81+WKkjDnSsArB5g95B405kr+JHt3O7YHhbjetq108O+8Fo3dGnNWOrgJ3JtqUMvG37RHWpt
8MfvEwHslqpIyOQtiCV5BS6PXQQ6WeQWBXk2lj8tKibQTVO3a+DAZ8JOeT4x4OrwlT0bqr7bmms9
NwryRbdWuX/ng3x2rT9in/+3VIC4xesjjn0S2m6ea7h0zVEa0YYCdWM8LJyFEXv4/jItPlZWROwg
6RsAgTghbj6WV9ZJw0+ffpaKhTI4uEua4Lxe0FNb5nw1oZJWgZJto0ixd9lWpJUfYjqY6XSky6bo
P1Lw+ul5x+dY8D4t0wXGZGal727weBeZqNhuIejRiHlS6NytplKwRSjE53+YhRUScO7HlHmNMC1w
yfN1VQFDsj8oIQ0ogUt/oFhILv08Fx8crRMOzeU9rRYSzXvH/WDJ+utxg141zdxJ94qz5Ot6zOEO
rC9DrexZz0TQo/CpDLlHD2cgL3vfZ9u1WohYAkh6RokBFDuyJ9D/N3O8fErSN2/6WYPTJsXS4ojI
d7+fGerK/OxLzjUjQFrMXnUmxMBQgfkqVM1DYzQug2s1ExTOqNTCYJ9Nma/3hNicQEG6xB9qr4qb
g5Vf9QuJh0njkyb3C9CzUMFi/fbcOGb2Q2H3nXa3DBwuy5a83ligAluOYzcpF2r4E2G5Ai19ADee
ABgmX4PfNzLnpBibcavls3UB7YOkaxAiWIS1PaGfOx/7GTongFaeqInYJ1XEOICRj3v89WNd+ZlY
0xUtW4fZTU7vXnEzcKzcsM7M5Q1SlnbHqWtO1oNCwjVl/RCcqwnO4s1vLA/c0U2DdLw5EbiiL2um
vQmRvbbzbEe2d6GP57PEtuUacP2k6N9zVOiNs1IAjN1tY4dRz0PWJVW+04JZfBQo2QIyX4kAmq4g
BQaqIxb4s/aAidS5VnDS8m9MlC4Rc+F2b6f0MUBJvmTud85tWd6+62mcXSVppmkmXNAoNmKIjh6T
iKPml1G1pjn4kvWtwji/MSZe/G8hLovK9H8eV2WQpPFyuy4ODkHVwrRq5kXpBhocHyJ1cOsKoGcl
Zot3RO7ui95/4H7fekxKyDMZ9jFHzaVRKdWGq/Vv0Mi1FhoH3VsL61KmfNIblTeygyyqGRge4Dxz
PJ2iSa89JKK3ksQlSOq7iHwL2WdpntPpzqcbT0IH+WGpt5cmCsoZOQ2CuomQpquNQSP3twuoOLff
iFS0YmuuRa4OIWq1h4z1vzyOdCifgRdcJ9RFKvUw9vdlCL5UwwD+Vt0ntCp1WiCeLapFqOAdT31E
awenwsoxxP/pnzNrpc/5qFNhNEg/fXVDjEx03V1FZcebAnMMWy0nWZGpcD/p1Pk5w8omT3YL1iHM
mR58vC4n3sjduThLOoc/oVgiII40WvLXKGYAa/P8MXa+c2rPz2oPybySU2wwd/OZL5fXwMpEK2G8
5c4XNUgjRmqkwzF4JvyxqsfoQVRoHnmhJhzSSbOT+ZSd87lnWwL39LcIou7c+7ReKDRHkcK+fegS
hBkQG4iyZVpuVOELKh4AGiWvm+dVCaaB7tK2gBgUij4xc1iuC1Ta68YWNUTWA6t43UEtasEwgo+S
1r+9mWUH5HtRgYVzO2Tt30tqJudu61L1gW5dJ/zEJ8xw8IoeMheOo1zYuY/uBL9piCmrj6vAuZTQ
ejkSx9hTqaoS9GLMd2Py3UA7fySSKzvPcQDKMIFVx4BFx7iV9SLZTkxyJSc6lIWDMeW+xwn9OiAW
dmbZ/qLuB+r/MulZyCOd8tX7hjayA/HNcSD09uGM+xMFSdWbOgflBOn0bn1O1q6Tc6fSHvsUmIJZ
1TiHjaQ0afFqWgX++vrQIe93KqbEOFo2nSWO8tXPEA1eqAhPYA39AePiQP0sxLe+E5TRx/dpoaqt
JT0fwqnl1O+ZUYRpNDzCFxUOt+I1uhYOh5REU5apKi42TBmANve6xYGPYycDETwiDEVlsYUm1flj
PZ8ap5nwBl9EG19vnudlLzsBXJIk+qxC2S2obZaK3mtzPt4YJUPbIHvotiUpFyb4RWcBXJ5MyTFV
V4vEdswCqz5rzNXsssdSJFwoR5E/8nv8HON4G+sWNprghmRT0ukRECW7U90FH2G2S/yyYPopbZ7+
U1JHr43EG6rbBB+Pps4s6564jKL5wHa88Q5De6bHxZJU3a9ZYtKJ4ZMvS9v2X4DLxUQ7yJ60/YeE
6TlePc3MdKUgbbMWhtbz2cKSsfXxhZg/nVp8wSiez/T2ndALNOU/NZoQJ/RDScIVoKcKA85Pi8Fm
AVVO5JGVTeRsYwyg5l8uYWSOZyAeyzhe9ZlIILjF7SYF61+71Y9LZRjVBqz/3nWXTu0Rs8bpJ5Ky
YRxZIPEZlaI8foHCd1qZAaIGzG39QYZ4k2zzizG2axdd5npJliKjwfhyEsS9ANm7JS/kMf2u4lnq
oJu8YutvmEN9tBzwky+y4AfNlsy2vOLiLPUYv2fS9TlIWEESVr+NxdcF+9a57FSGGhaehKCbs/Fc
QQp9jZAp0QRenaX+JI7JUPwT/fdR01NNhxtjlCEsT/SkA5C3o/YcD+Lh27Hb21LJ+23DdQ8Jg/We
TnxZ/TBGxuceqnJa203cVf4y5dGrg9bx9v+fqYRlT0JSuk5FJKPn0W4OIh6CnL3Uka0t66nCDe5N
pVo2UCJE6dSq8e89AMoiKzFtqNJ/NMp+oXlMA1S3P3UjrmB1vuyjmJBz1OMvkuD8MHcujt/MzQj7
y6hkgF7zgmI9ECfPENmDP0DojxVX75DI8LLHZ+yptTsFgp6JU6W38kVmrJ83nMxBVhAnsPCfSlOF
P2NUCk1NuWEF+oEytuNWB9RLs4lXfFTI38IxY/4fT/TClaQMz4e+pGU3AkFx4bnSUBnQWGn9xuYR
HpYZ3NVLBNdC8MzZk9XfqPsUdbKG45CMExZMzP0ydwC872wuCt6EWZ10OrVx/72m9dq/jkvxChkG
UkcqASofX2/uyhWfnBDjfuRHGpztn+5DxTA16FxNO5LodES3GhNeZk9uDZuAWu3UUqwB/NpmZdE0
5URICJsi2UG0A5bQk6R7QB6sX9G+7R33LDiJUVFvHsaAr32c0j3IwilCJJcTYraNugNSF1w/q2Ya
6UeID+5udvzWgKqGigVcG0QwlXRKku7xO2OTaKUBCMdf4/XD4nrYCZ1fJtxYczznoPfnyiRnrA8m
9+tr8k1RQt7ypJ5+sZ3FqIbDzAxjvUAnxypEuzALeRytGSfdVa5hVft/3/RXlrt2l9a0e3Ej0u2Y
zg2NRjtMSzYgjQpqKnJvM88Mfq/ZAfzUsoi06TSb2ECIP+w3iiJvXfXtm8uVaLmETrGVtyS9BIQK
WODVjoFUZX6UVdjLCNZVwXhyUS3p0l7Zh13uxN6qSh9wmB51YAXPbeKJpVKZ8L8brdkav2aOJkEX
FFXYaXp8evcJ0dHkEUj1nzU770F8juiU8gcDZQn87hME8oMxYUT1C+/GbktbeUA+qTB8JT+rhiI4
q4wnltbvBiS0lR7QBdEz0UhtTu2LLKDrh9vTjXIWk4NvGWS0aKhob22uSRyPHNgyQ/XXktmP69P+
mC96EhvOrHJVcaSeXkv6sC8GTF2fhx+2fm2sjELP2J5Zmul/AckmRaE7+mDuLeJn0VjfXMBxMBGv
KappHBE3zUQVWsft5M92azqgkNxRJaRVigLSUk7qWA5WYzzC+HjnMwFRN+anTWHt6mlhpixMfeaV
4tO4/+Obfy5RuSE4/VKhVwPfgIkGuxKiVphNRmRVpeTn6G8UteoDEg+NzDrX02NCbbAiGcB81VYX
5soD5j6BEjoT/PGkvBPp0GTujdxznU/9t8Ot1CdYjPfErWqRLW6GxyTjl3WYDBpODKFl3+cOXDQd
oktv6C/lIQHHowAfT4jvvjxtD0sd4OvnPC3wgWglCOtQoxbS5j7bj8rUKpFdgSmdLJq2gxlT+wjo
lchElq9ZV3HLU2q6AfyoXh7lxObAkIRFDZbETFoZsYEvVeiaMRVvnWECmTTDvxOUgy/n4CQSMZ5G
ZKD8sNOeePryMoeNq34sMMPtxDck8p7OAugiPh8y52+hNMBjLtID7MpsDUiEtN2e5tT6NcxcPQrl
GJhQTI5xpnqED4UeUVflFcgBVx6JN6ttBDTcuxsgiH9GgOj3RWUMFV9phCFmYvxswv6QfodBiNEN
I1OQ31DPRFhiwvJ5Fep66g4CDmmAk40mePXte/51E1t/uD4/pVTORYg2YD0WYvU5x1QBfi5Xy9xg
3SC9k6PRr/wt4UIZ3a402nsMQ4i3zoBOy2gukcRzGl5R1SWNMI/tDKPX5nWHayxuTQHrqAN04DjH
wgQ2z4CaLmErPC+oliT8tPHufG/0+7BodvR4nGbxmtH6MA2B6luqDJjrVCN5C52ZlFQicnESUSqb
kgpKM3fUwVA0xceN0V//E4H6LgZITdFH2qhJRxATONKEhq4PvNAvrFPS51VN+e1oTiNTzX5H23vf
8oX2HOuCmwQN06PCcljVDPuhagg2CqSer0cdK89mgckazXKugxGSFiac8LBHVyaAsqsYnVXOaGIN
vH/VdE1GCmPwZ4qQ4NJO9qm/Xw/Xnd9tpWLQc4ZnK4h3dOxcdgJQt4uUPacppquTJ78VMxWsOqDz
g0DXsic3XwW1GKh4/TSPOdGYzjmIydymwDbv2eD/lWmZN/rYdj3zjVIiGZkWfdA7XprSCxMKs5Kt
UnqDZ9hActTwYRMi8vJLPJSk7Hs0rUygmns6UgQFmLnEFMzC/zsmMFtfavhHcNrSq2M6RU0CBWtt
opKJs65ELWIKL/ZR+3AklcOBH0yjaV+Z5Oc40edr9MKIZHy4Zqzd5uhwNlSYRYX1NeQ2n7HlGwkX
FdDvdp0hHhta5QrI4izBxX4z/zdzSjxclP6piIofHJpZh3VMPt04SmMnBxjqIv/Cpy7a2R2dtx1i
c+efI+KuNelW4VItJpe2XW9wYQVuq5kT4JKleHQ7elkiUFhqv7sXNaARdhJmYE5pVBcbc6qtWHpP
/d1Q07MnX8jH2deYfgMHwDkLRHLqvX+Fv/0dFsne4bAZBuR5udMk1zaZIHo4htP8GOribnJoqOI4
2nvMdyH1RGe5i9wMeAg6aMGm88I8c1dGXlnk6u3BKnC48jkb3SjLY07hRNrOe0fHqdskKxfZjpEc
6IBecm0f2u6Io2fb3OnNCNaJYW8+faii0AyY8B920CayV0ukxBFbt0tkXMZ2LT5mfhL25NluXqXj
9q16lDRo+KWrY0Zzlg7iGqf5lMFlHer8sreWfJUkr0TVoMo1S3ngfjbjxcjfSJw4wulI88AvRScF
o3POEfdPj7NGe+17EbauOBKjpzuHQEzZve937F4l+M3qbHhHMOF9p/GceZdlMx3bLBpDIpXwhiHe
uQUeZrg749o2GZvTGqRE+pEYWafH0MuVi4OhSaqtaSwOX8WegsqYMQJzVkbdswn1T91M26UH6Voi
FVWkMGhzBx0X8uhp8XXx9IRHWcdgNmr8JeelO7OwGXbNjfSoKOLjG+ixA3PApmJJO9yFlvQRrtvG
Owc3SISvPd0e4dGXpOTrDpVzXOvdm+dgZD5qb/X5gwdqNk9qI/dxAQm37x6W4N7xEXWhMo6uSM87
SJvS5g2IZJAzw3ZaYBCs/wz+UGqNM7DB6OY4zhtpezIybv0V7ngXoroggBMSruTTsbukbUmldiaG
l1dkN1qUDQYwewBmn3ZtuTom+Iemk4p8gG4Xm8QF3CXMV83OIUJo+lXlvXJhfKmbrYZvBGNaQ1r+
Lqtc0FwUHTfP0KpPQNqexQ6/g29I0v4Qr6aPcHBOYKg26C3gV84CNMOkZFZ9wwrVbR89Rku2yaL3
xXF9JeBxO7SESvFyWebyavmRMG7RNnBwJvpdu3ssVLUUkOu5x64y5Xk8BxTvg5XRXw79ePrwGgeH
pcbvAX6VtlvhQ3erLf7g/WruR7iTOkTi7lBPNHgeYih2/BfX3C1ha9ecnzWo6zt2DUkMLbsesDHz
73/yWbYrO9WtkZbXph5KmMPhbJmhbOypLuXw/jbo1e4mJCPg8KO5PYUoUx94tHqRIBITFApk8hM6
HNhHNRmxz0N1y236JKMD/vgaT+my9cKkPHAkdaTWzOU6BMMqWBSc5CX4VK1f1iSwkkJE1v/T4cN4
fR2rPegW60Oe6mGk5dQgaWymldkJBc/42aUBXcU3i0D4NDonxmgD/OE9brrcxyMUassJK1pBaR26
CJs+Gre+9NK0pEkPAlkfNtztgD5wZ51ECCfaEhMI0leR8qTHzAA+c3S8Uyq1dbEcyqU8mBV9txPV
5ppQEsM+e9c0+GrnX+DZxKFDSljyQaNSNvG5cymE//GO8U6Orra5BJhZXrWz1tSFl9aic+QAh59s
L1OYZeXEO75oDtGGKiuHtUiFtUur54AdZ5iCbPMJzlb7rVkktVvyJvL8yzHPST7RlAa0JnfMLyf2
+C3j+qobkgQI/VL7nMffc072qW+3HNWjKZV+p3c8wFi5kXzmBG8lux1sNzk6dDNqM5XLb4zg+asX
aeE7gsuIbWPq8Q3Ywi7Y3ew1FGf6wrqhiq08vhU0Ceuo4TC/bpRhXwLgn1MxzmkMXrH5rMyHH3Yo
ryTRhM8QuQRMRh7JBaWMQ7MWaPx7gDAuSrDya32IDeoUSZ8nCjn2WPwvheC/Ufxs9kTdaA81KjsJ
H7pW5Qo2kq4/O2yg2VDk6nBeojmEz3BdojomFt2Vcao6svCIO4ucaRG1zWCX/NnaAboBHT0v8KyE
dh8oIWVm+Tgs/QA4BCNHNrxnNRxPPxvzzO7I/s0vP73hPBzOaJgsyER1NFV1lfFaG2zZo7hW1SRk
7wV13SZfp3W4lmp6B0Sp3eD0jRtVre6x/q88pSvrxKC6bGmQJhrh+zbYygurJqMVK4ODr1psYWnC
TsNrVpV1ucMV1p2hgE2wDCURZEzWzVp9x1wciXjknhyMwsYdGbIgtRz6sHVXIIvmdoYm0VaMzzEf
8ZqwQxNNMk/OT4rHqlAFH9JmTGUgK548L3IoaCPi1tCbcvPIyavXA6BSAysMkLJeTTvG5RQGb8Dg
vIp90bJ5qnXDyzFu1IQs1iGVZYch54qOfhImCk7q+kRLvBrIGTbOmW9EH2BA3puPcXTVl6xh8KL1
LIY7BZao4X6JklaJqrIBMZz2Bux4u9xCDHCvG1HtfWngmKlWaw2WIPXsuck3XvYRwKzBzO6HLcKa
FUiWO9WIMXBNLpLXzWZ3C7FUmv4xI5yOJaHo2U/49ZwISdubns31D3dbgNyXfiYl66BN3fy2jaRG
elNus1x/BcKuihaYnftV2Mk9PubPPaKgW0R9WaG+6ELuyKj1jtcq24bFOe0mtxe9b8mwn7E3z1wj
Hl2QV0aXTJ8Cn7q9x+2IJsDVv5J2IbeKkz2u5AwA8LKlMAGIleAlr+NHQmH9b6N6dM6g/VprDPPs
F81BFSC9lUzLT2ATqSrSanhgkErFkk5Ue1BPa1A8HnN7XLprDCvGlQX+UdQmeMe5kp3sBfVD982V
AaCqhe9Ol3RXSlGkccY6IRZi0uwvJBeQoupgoaWwzlM9y6Z8q/J5xnk0Wp7MdsEo3q0klvju3hR1
x6BV8yoDQHtNcUKLjVCD0PvMdvRBMcAf7ONUGSlqo1mGwJY+Z9Z5tkb1G/hYGxSOBNQI9LGSKh1X
cO0S3PC9R3ro2fj3nOTIOz5RQ62iVTqxOhAr70pVX15UjJDI2VRkfQxSAbN1VwNgZTyZjZNzhDch
gmZukr111zyXtcx5n9u9YTLQPxBxYKjJezmIJtcrPIIfPskK9zRzK5etZ1RhEbtWLWx0pGpleVOt
RZk2v9pTTe4FNhIG7E6dJ/Txg6GkKms9cMZSVgfk5rDfnM3pbS0WG2CmEOyN9ar/UJn1g4PUYJix
yOOkc6COramf6KrL+q59HO+uWhxwhdgQ9UgDgXIN9Ez+L5zK0WoE1v/zGyTRZ5r0ASD1n6MLyT4h
J0p34gf2HDS3HvnAH86vudU7m1Wz98hg3NWOOaeh/GdlxowbSu4ZgzLrbOGFhcpAMEgpfWrU0Mww
oBBDui8jmDixTHmGT6DDKK3/adCm7u67Ydqsh3gAGuxxLnm9e3Hn0RsSW3X9eCW3SJn9x7rbbjPk
yWo5H91gLW/xwpswKqvG2FudtsLiXP8IqzEJNYODlGX6v9lsQ8DcPoYAJO7+s/srS9fY4ojHcShh
X8CIHOJD8fURQ29/6D4Qu0VK/X4rp8VTEUbZItHbkh8T+29md6QPNa6ZO26uJ0LFdbrbJbZIau4d
3tbb8/3YApP5qPLRojNiXpTqKYJhBRLWeTa47S4+arrV4DfF9akkaW3ii090zh5hU4krY8eIi0o8
jdthASXECjmwEFz6NNNkVbXfm6wjiJ37eejIgUDKPXmlMJY8WNLsSFHYA8QsQ1bccMHarFLc13Hs
uGtcFqUO721N2j1GKScTMeKXhkd7AtNvL5wFbmhsPYivDHNor03aY19DW84JQVFslobCsTzN2NsH
sfjlVALYsFxLTha+q9dCMXXMHexnhV4RTEn9AFrmp5mSTqorctNIBocJCSyG/oWHMUW9ZG9x15v6
/OqnLQgcNF2Q6TAJbKx8sYK/ekLdcpPqttDK4Ox3bgoYId41pR7kYBVSiHObSAxxxN214CevdtC7
42q1Vdap6L6nRtOadDJcSThkTpcO/THUHzk8bvSYJdFm0zeMhzp/BqgCAjunurQwq9JtYR4VBrqs
SPqJ96qMMmbES2o53QY0opRjccMuXjD33M2L6M/8I3y6//sOuT66WaIcP8pszN8CYXeTZnzfBt+f
+6jyNfB9a+O1PphDNqiRIQfX1GBFbK3yAQ/39Co/nIGpbXQy+GvM/eKKg5PzUQb/+ChVq9jQNkSZ
wRNaE2AXt+/i/7giImSaOB1LH8phMor+T6cMUu3Pw94+uwW/oI2EOPMcKxXPunfGTMdACvh21tBf
3Du6A1sU4jWJtRRkPiaLqkXxJCeSYk6S46jtyfNN4IPoLpkxH0BwUMu7/CcP3jp5YgAZqEGjk78r
EMfgs51iaaunZ9VCp5D/ls4D8KwarL1snjuIT9V1h/pnhB7D0n+JGokZB56n5EwZbimlm63AVLEA
Dppj3bUYgghHtp2ZSKY4WIQkQGMOHPCmL20DAszKuvlBl814TisgVWJoZnT1Hli2/eOK/jX+TxvH
jwBSbtKYseIwoSgF/Pxttcg57HE99hkuSWje74XlTMRASMPtdhAXktso2lY+as8Zwq/k7pt4oOlN
KjAmMdh+z7rcOk1vEKSXa3huZ8WvS8CR0tMK5AD9NglJs/YJ4fGvoWtQc3nNjAgPqJKmwnjonk4C
gDr1fRGyyETtq/DCS+8551HDrKzr4io71NwlNZu8jMnptA+qQHU2uJrYLgE6E2TvJfnVd4IJXp9n
O1/ubq3VSA2go1UmOa4ucLLRnrddWNSmNjcrlnz5IuXY//rcwSTQW/ZnzEja2RSflLsW2Zvc/tKe
lU4/aJGfCWnckkdU2oqk0BzbejWEWzccpBpcTfOnj1suhflugz3DRRA2L+ZkLzShNW6LMM+ikjsc
2mipNFd+XPW2RRzCQUKgmp6qGU2GGfyzka828WOJ1uFAfT80EfDqld72ad00v9M+rsax/UDGZgoF
Q1wxItnGikwk7A1UWNq9//ATQqCkrev0aEtnRPQW16LrHaoGxjrSQFYeO+A/9AyRPc/Kqg4gTzaa
v+TQzGUz+YT6JE6vdP7+gdjKqsTg9pCwcCT5pLitscfUTbZZ5L6DKw23DzvNFGnzF2SXrgUCkyIz
aX8ygZKJdIHh5ydmK0RTDyfaXrGqCltxLDP+x4+LB3SwG2FIUgLP9Nkdxbq1OIue64QL3sTcl5mf
3JYA3oSwdJjjDby/dkRPVnkCRxljnqdj9b2bL4A9Dyu4YEK86hDnGPmGpDBDH5jlCL2etaU2kZB/
FrjKR+UgOSi/SHmP9SZ+U+5Ed1KaVxWruM681S4fiTxNexKAK9Q1qKdYOLY4H/TZuezWiQ/G4EW+
dON6iRw9Q67x8sdNXKpiKTQqnizdXT1gcpTm5FqepYcIyrJIe6RRbFSSGD4A46CuFjGBb9WL7iGB
sM6xc+aIL3mgQ4tPXu+VAK6QwOsHkSg3a7jlfZI9M/IJMfE7bmVpRKghiCgyGbvYLzfban1L8txQ
D7tUC63ft3NcuMrvFpCWjkocOjL9ULOCFoRiqMs0V+mNdZcFGrA8GygJh0hmuXK427i0caQtzr6M
XNcBvTL3RUfhEnjEkKlPLZQ7C/cfVajGKbpUKM1IycdVZgQe62yaoSWvMMPb0Bn/yEeL7YxBfUq1
wiD/2D/DvI+eWu7HOI+EKx8JM38JZllyG1VwTvXoo7z+1b7atyPzsy9thKtO/xYR7z5Mmtscmeyu
OL/V4TaGfLhvnhAzTx3/n1IO27lq1TEaq93cxP9bah+7XX4ibfORpj/iXHdceHDtGugATS05nWOZ
UGhtYjZMOqRd2rPS6R1L3th1FJrIRSLzdgTlxOlo6jLDhnsQAoUtXg7OXjkWELNKiYjPE4dj1ty9
G/bv/OyzL2IlmWzghgN5W5MgQcCJKhKRhEmUrMgNhwjCWXyhLIlFjcbCMZMwWm3/KmbnEMFKa3TN
ZL00aLC6twUcxySGykeVnLHJW6KqqpL2FfHZvdDWby1BLHBGruB/K7BVIxc3WkfXVNsJwWwV/GeZ
DLSaecOD0Pf3LpsvgHgA8AuoUc7Jl79NvAsaVZ+we4Uvjy8XBF+1wFMTnSBgxVDf2RztPb5TuMCH
owz4ST6oG1b778Zo9hNXFYiAUqhiDRmXEKXicIN9HMilI5goRSNudJfzFTi4FiJDM+Ks7hUlBj6e
36UnqbLp+pqxh+hw1nU4jmBA8wKe9/vLw9FJd6d76JFRbCr24mT76xZM13STUIjSeew97/wF6Rj/
QGF2X1dKcK9Swn4LqhawZJVO6CJNpHLGoUJRFNnrs3yEtgt8h2aSqicwgTqzfMfXuCY1BnxRzm6q
JQyyCpyFZvshzaHrlRk69w/3O93wgDVuqtJeDg8oAo1GeL9GwL4yOUX9FGDBtQ/J3fJoP4PSvq6u
kemfPyPaG1Dmfn0ehJ8B9end3aTEJOTKiC+6nJp7vaBDcsYG/Ad0GN1f/YJqdDfRe9SaqsAJXjwz
nI3gx/klpKKp7U+9oaVin42GeGWbROM9RVJQAi4+Mag/Krbm5b72StfiItizdVKjlEyrQCyyd1j6
5b1N4nHCneHTFfUaJCASv7kQ/TOwM6r2/V3z6bgcCgoh1kH9TBr/s++kcygtxSYd1o0yfFqiX1F6
lgzwREu/jdDccflpATJqQ+JqwPYLOVjAxvl/C77IzvyvDzWJI480srRGoR12yDuQY6UOn94MBApM
RY6lW7fy5bqiA0O/hLspcWngKaWnJtfarKb/LXPkmZgMaVL8AbMfyHLkW9GFL8Ao78wEdJhlGUfy
QI6jxxuQ1Ami+GlkLA+Rwdxu7755uycXnWS6XzDUt9WApe6pwxHN6Ra4SqDi0grfhxt/Gzg7OhaE
dOeosRaYaAWnGI7HRiuTruwg8Dms4ZyaqQYxEyyfpBoG603Fx3fCLYeKblG13Bif9b16VOuDU1ZS
tOVTYwHEVp398PBJKdmsw7U0SAtj3yN0dAeeUBQNH/m20nOmGxJYHxbaKVIjKHrrFvfv+Q6ah0Uy
k/Ydxf4J9Y1mbyGOIlD/se8JK6+JO0ZvBorsL1KjFifzXDLOesQH7WKXEvmZ8exTtkmJV+o/yqtF
08gYiyACVeE9WDFvCum0UYI7ezfhGWWlLDKtFYiXTMq7PnxZOpvr55YD+A+c+F0ZenaKSCknjcFu
dig17ncildJjNgbOKQj0fN8QzxE/ra2b84vkE9iFgxuV0DZmaVN1ovT8MA7Ky2xorQ7s3Pocgxsq
X4659C5XfIFVKJZdbuHpNTgxvi+HNXKk16rPeMyoEtJumxjgeWpcS6+Cz4H8acSVYwNS3Ub/ZOHv
kM1JtJCSrx8MgZ1AbT/4p3uc/BA3Yr/Mh0F6XhbaCx4Idticy1v4IEq/6QLX/PAbqaAcOBqrFLuP
q2bP/jzPgr6caOEl4WP5lCaS7opREjJyZMQ+qAmMJ6QhBUrLaHAeI8a0Li76Syn7SuG96W77YjNY
7JP/zDRaBkYp81ouUzlDI1vJTiy2YjcNwtEH3H0G5vjB6wz6qbAPHXPD7B6yk7CTwdBRqFCeXA8T
9pT0O56xS5GglP+Zdit6/rFy4XoQ4937T843kOmG68wNmshl89h3LPmjMFfRsbxC1MOqRLlTW5DI
d+XBDt8EVcOifFKCkzpw93wvgMptI9ckNPQSBpj1PaLFh+Fmw7KNN5Frq5nT+aFJaNojyD9cv8rg
DCdItGRpNPXRaaWfFzRgHQ8xGxTj7nmClYzOa1XJsN21J/g2RORGrVQHhXb+uBgsIEYNiJZatdWT
ZsaJsXNOkieiIKH7dpUILhQF6syZ9axNankvJgCdflCzwdEfEzl8KjyW8T2TTt6/8F5AQ4HOCSFq
R1158z81KRfww994LGH0YXQ28gAhFKEvMigQVHCAvjgtL9ZEEfa34dIxr2VZ/RvK/l88FMsJlQfk
lxIcYP8Zr1re8iGE3dhew7WSaM8QIG6bkhT79D1caaWKVqbupvhWEdMSd6OcIJhqJVA9xCVxfnAM
KcuSZHD0Qqth7O1wIc5eK4NUZx86IEJRLBPXO9toqJvHQqhTdUAI5dDhMMChnnT7Z2urssTGeNBx
si5qvn0AIjgq8FGDAM8Tq4tKbqVAXSUe5RXNV9omINguG9H+LDv9Sugju58++sgKiQXdOeo9x84Z
gGsDGRoZOgr1l8bmfbPbaYuA9+BAHubY64YiLfMdMkXHgB/bDKWQh/v7da6fnfeonyWjjnGqRyyO
uMkqKILGLxNLEFkeMDFe08Ka7kI59og37BdEqIvh+LkYpbUAHqKLxapDLB8GrNGsBHd7QeAffgxt
eBqtnT200VBLfl3qB9o78Rl77GSrxFQzNyiYuQUI3GeHQ3KAkl/qPtstEU/KNsTW1/qFlqipJKlp
gZJM3Anh5dOw8MIGAdFVutm0Bg1nx2QTDGZq51LlHUj30ducs+zueWCaTYwhMgr4C/t2egMrtnfg
CD1E9UCEGwnzw+iKaJwC1/ms650RKzStOhW5Rh0L6+Qj6kZDnkI1rxKYSbI8nVnYB8Qp/YvoqoMH
jIxrdFRpIBJBfAEMDGEaBrGPzOcfxVQiommfYk8cZUkE+r/SJXuSOTmcqp2JwpODGWs6ke/rGivm
38/MeZpJEzTseCHgP5Opu3+3EY5S9XHFxQW9/SIL++knlc4AFtiQr5+xFazZBmAETbD32Jj+QL+E
aJiZLpj04KU0emgsVXICFZMe8Q0CE+IHy2bW2I0TtRRZ6YcG+GPwxiQa9IUqqI3/c+QIlxC7zYR4
+BT0D/J86Z61t4+aXkzg3mG4QbQuAHvDICiRVEEx+O0Mnb0HjrMARQlfUV/iXL/4xP0IyImT6Lwp
WrJsCYMEQmzASnyS2XFW3wXl3S5OO9g+1mQ61ABMV2ejcWal2NGtwGB55GFcPa6+9Nc4BlEgGUtT
qLnUzKIQJ5dHOvfO6b0aFtRaiB1Q/ZWS8fkTRkrhEn0L8nsIQYt1qLAdGGoP3xbxl9GQOSLEgPLe
wS7T5kciy0ztcMC7Hzk/Nw26v0D0kUYtBQACfx7PTlveTnBeuSiaXu3xzhHNoatj8Vl2vfgTV6HJ
HraDmPbRXKzAHY+I0nkzazR5MzsiP8Y7epRXOEUfdr1aqYvIGi42Bvch0kcltQl+gWoQtE2nPZwj
YxiMmcmjsBisWg+XkuVxz3jbPh9/6yxNoJTCha9ghW7SCpfQxkx4lkD8Y/DvtXBdSgB2QWL/P5Ad
oL5WtluWZ3UlDJ8U7dIb51BdX2+Dw/txA3iSz2V5FQFfCyRn7ZbwPQiZEIaBmWGcEVv9qFI1mTns
jDE02oeN5m7c9kW8ECsjhvBOTKSfmiImPoJVPc0tjlt9417/b5YhZCVDwECyab01z4JcP4jwcCgm
LSMORkg1aRmY0tJblknADtNVsozDsUfjwTwceDk3IdCOVJHepKfmWJK/Ly8/V04NJkWfLLV58TqT
82vdaNvBkZg59sALJO5DyDfKa5kj7e516kEOSWqFG/mFTpTIbjWDJNdbwsXs8vhmSIm3yhUjqPh+
NjC+ThKvBtxkNf2yMv7kLxFOaFHFgRxZIl5q0yCOF6MAXT9L2YEEXPNyeIoGMiW1qD+L0kMkZ75w
fxDnRcLI/YG7RZiK9xrMZDuVcXHaNvDCsXsl4lUzkqV58FDYfH8S3XMemV/5qfeo49xZy5QMRe+a
5k7qfoeqkCOInEv+p/3b30OvrXzJqL5/zC4U0FNcROBUb9Y5Kvkrt7bp4cLJDZeuPYlbOrgfPqcF
GIrPMBmFEVL1i5Kskq8fC+OXEBZD5zMG5UNbhyfgG7/+nCN4rkJjCD6mCQpOGYwzHoczO79cAK9b
WDOu2/CC4gY0tRiOoaeLFVLjd8IqJ7eZsRsQTnsikMyPx6JHe4VxNwoY3qC10k6gdywM0BsW9Def
y3hEAO1O2RYygIqldkHWNjUqTOpzmWQ14DKcUmTIV88gBN/XF7nA1d7qOZT5kZk97VPImkA942LC
V3BWYaTs5RtH1dzUfMDcvezbi+qFW8+LD3CrNkn1S72BxAsMqvaTmLKBhtuH1SmpdCCZPC9Q868g
PoBe37y48XrA8CWSnXsD1VSOO4sRusBlN0pLU09ztJ6172C3bZbrIy2/WSZZg7hDnJcOsK907hc1
V1n4vobUjFrdieQ9dY6+HT9TnSTmJZK2b0fjQ2R4m5IYwpliwonvwQft8YdEYonzHeQfgmtRxZWI
KnePVRdTr/U4zCzwIH528cQyE6WCqeFhwbm7EausfXpdBFNLjJZgKPjTSBvkS1AbyX3ucjp99SDg
AVXl8cCML5UgktD0fLMG3OZ3reRcOy4bVwGbG8vIDNXem6dXVZe+HJAErnCFSXUOFMdRhs89Hwgn
ybgS4ZnTO15Jm6cHd6/G7TvzSgqfSzVSX3E7ybF0G+0fWUkvUeJOWS6MXHchzx/dxWxljUQZsDSp
WBHiQ+Bpw1+t66d0OhvfnAv1XAZiV+J3Va84kmStTY0bj+vwt2DRJZxVzm0a3ot4Dq/B8A5mM4n+
INkpN1sl/hcg85nX905bjseBIn6XFnUYbIbyssBXJBvMZ7x67TTeBF6sHCAobpBPk+XjxcK15OoE
yeBuznygrn631RtLlJsCkSJ+PEHHQ6AZTkdo2g/afZm9dQsvhNeqMSRulNvVsKmrVQ7r3QMaIZs3
No4yAy/TsyB0z1AVtW5ntXnAilNDDaqes0mnbJLt3LQj4ywG4b+6OmRifSNXwqW9mcw8KosIEM47
Nyj1F61jWLXcMZMRe1t8q07nW2RPuA39RMfXT4uGbgzRr2Fs+IdVTTUa8XmkgKaAcJWC+SaMX6ig
J8zWGyfR7ryxdpeDkW7SU4faLIwf3WmhLy8MO0Dsl91ug5dycntYKa68ZZEbP43INODYWQS9NBcB
1fG0xJ4dQPZnjONSChROaGJCxsLDQN1vvsagv7FJiJoSijEYqujg6uvN+88qGJoRhavGupMiHBpy
0u0n/4zkvrJBUyEZ8q+7HCxAjzQo7+gyMFy2Xmo1+nxAAlvp4WDc7wPSl6DIG0XRDadSarHAvQaO
VjL8aCRuPUhCn7/9p6EhwWvvuBRLsopLrsDm4e5o1G6VQ+T0UTFRvffq+H2OTyqRrOsHK20IAHmE
tT1LtowcNCol1DRp+iZ7vPRC1CZtrtgrjxjhoDwFqy2lyOY6KHQclDPe6tasHWMWrf+K/JUwhL2w
K4M3sXI3ol+Iug74TY+VNaWtavYbEUwGJqloLAj8dUGLIt+YBSSZ9kqBGJpTaf6xJR6BW4kfpzNZ
yBdw1G3lC0brvJdpvxyvsNXMh3iuydTsW7nGOLwlS0cfI5UjoAS6lFOgpCwR7dr30b1Y91SwCQH7
JAROb4e1lijzVesnSZ5FYlFHwLW/jTF/M3Z9ABDvza2KGt6D248Mac+V9EMINixSPjccElPRK60R
G2HvRJRfvG81lrN/+eljVYwtDFhbYVUT+ieUFImaqMxORRyMajmw880QS5+1s3DSfbHkcvg8cPli
5PHVBLJUd2H8liFjdW4h6Kmw63mabO0XKd7DUY0tSj/CIOelDt7n1lUN3QwdgjcKxEleI0F991U1
yl9IfR9j8Z56zfmHm9tU0r4qzWwsMu4A8h1muGkYR4Qng0uxClXLlGDfS0rxsZi7GX8mSH/pdK3d
omLhODVRbduW/wM/e4z0NH3jm69BmLRNeB6Ah/x4FbyLJj0C3LbV/tXN3wBfiFphXaFOJkFSseNz
GClkEx7NnURHtLH6H5gAQtIDjTEQFZC5mtQQvGenSrn2DXysLCnw0lNr07Cxplt3hHnItpT8jY99
cI/aWGBsoTuM6RVqJpxpl1cXM1EgM2zH3OvhOZa/Jl/GK9kZ8+/ql6/OnY57a6A2HtOYZ+6CBb7P
nNnGz1pbhQNYFvVaqGrgFovwjR4yj36Bcm5cC8JrMIhOJEMzh+QdVpt0p1NOb8q1/An0wnsugGo9
MsOWUZii1MLuikR8Kv3f0SqLbckGpbj6RmV2f8LfF09L9TCWcrEhHGGS+DV8tK7Ce2fBpgjRdQ7Q
WYx8bYSqDy+Cbu6DWlnElV9MqBMPXVnTSMq5q18CQSmuBQdoxaGpNU0BwpWSWg26j0lmzP36xfSF
/aVeNGa5ZyQu+J3L1mHtH+bYtxYRhRdX/LslQTR5ph9Xj0TsEMVYSZIONsNOgSAtNAre0wDfcfYr
xBkcgDqbMNTRGfqjAH6HJ7+2v5wyJQledtIjHaDDSvybH9n5GKrj7UsnGRKAcXUji9Z9ztw3WULB
FH1A42mGbAM3XrqUZ4k5shHMTXI8gVQlRdMlJsJ9idT3DZPhC32mt27rpMfAmW/tjN01IhykbEhG
wUdptONhlJ1sIxvmp+4i7f6snF7y/yeaMC0kqY/XPSTFw6DZuk9LVFeSz3VpT7zHkDcHyXcCC2ki
UWQbdFEcWnUI02ci5rmoS6hjbyjwr4ssjlElifoleqw0rp1ExCNghGX9TVnZ6MT8IUjkmIC6oNbh
H8hNB6mkAGoojRoo5/qsZY+nlbqYjGrYq8SlaSvDImq1r2q+yLHwqMUHSYKY9m1wBIh4dJZZVxBe
AtSm0XJM1nWZU94+DoYJweO3cfP89ek+nIAyd0amXx+FAukY4TeWfqPFqrrB/oE45frGRShLrt+c
vVWXUUsqnTZ8Ic+9f6oG/RiyBg3jqN0ISvTuCiGJque2HMcrBZ4BBGUoFvyD7nSjdVhwsAixxROo
1hzu/Z6KvvP9bzb8lUf8OGLwBRjSKMrZUx6r9Zq+QXgUhLv3UAxa9TNsy3MtNtuy6/+F1yQjnNKh
9M+NwN2udTM/+c1VCVVR0NkZEhcBznmMWoM7a5LB7lKLLWEGq8d5TxOtB6fqyDdnYu4Gk6WkiCdF
n4KFn01VANmBkC+zXVXpTb7eZJ9sbRWz3FPDLmFMJwNehm3XzMRJDQFSvJQIErJtW85Uatf5J6eY
hFCHvLHxYT0zOHJCDp5WFW72dJ8mHpESBBguBaP6GGsyCsW//l6qzkrIuszGO/2mhJuXEfOXldBX
hVdSE/hrbFnR5esWHH229lnggbHrQo5lK+p/HnBIdaOcxE5v3O+sSakKk+XzdHtvAPXjB4DO8X0+
1fwngZ3C5/HsUU0Z1TbBKn0YcMi86sscgYk0BfwFkUxd4weRTvint/q2HUmZleFCb16vjWymbx74
9lLVftevyD4Ex2wQa6KYJh2lnkUeNAvJGA8L+mWXYV8wCoY5l1YSTxbtSwvqIVIbErtMInZmm4GF
LAV97CmNqm2UOd2c/SkoinULiWvPxS6qtEkSwvJ0qgVzOAeLf8rOGEWSP1RMonW5n+OuGM2uDRV7
ujluftntFTlH5VNV5sRccoGqU3p2G1fVwPyQR0bcQx/oANbm6VzEfTLx3Lijm/qb/pQ8VTO1VF6z
VWuVkAdAkp2TLwZ84IYQStgyXgDDz3jZbCrqYUedYj5zMcRAFEAdESW/rmri47HXKX+oH7qdeM8U
kbb9kWmiYdwxk/qdgi+3yS79U5cgobH4oLtkxqIfvwH/NaM1+9UVksnWC0r++4TIB0aBi+ejPo2n
Ux6YgYpbRqsNwGwNPxo3UccauUd0kN8nQU5eW4wc2KHU5+qn7NM6dABnW5QHNcHR/Je58fnQtkl1
vOibz6PLw31W8L4Dl4PcwE84ZhqiG5aV9tUh9dSd6sa8sXh5AH9yorQb8//QRjwa1Ya2TY/39Doc
91u0VG6tIAwFfABK9XUk8AdZ9DOQYVhtSgsBLdPElQKLlivT47/6r8QquVFzYLEPjbY+Po13WgAX
HAU4O4e8DJaZvqwtkLEyKpLTxB7EyXMIDmeVpgRqIbMTfvTxSoI/jIUwhWGEE4Y0E3Ps4tJTW9Pu
k9rEf85L5ldkluPHdis+7zOyC7mWBLElscmbmu3Xrdr5NN0HMiGacQWvt40gTQKYTRMGyxyXVxsH
nL2UUckalUPBTVMuGscpMIV5biasgsLCEt3obPuMlx4sHwn9srZsfPLjMrO4LGmu8qYDqwF+JRpA
6FJQDwrxyvZ6r83fneQbjE3LqELLFXehZJNpEmbhh9iYJyfFfHn41j/O1qxJpGsUfHNXMmC2Nmit
mWfndsDKpYmy0WJPkS+kH12hbzGuuzhP0+Mow8Sw4L+Dhd3FJpdOos5FigPkOXSWt5hbYP6ceU3i
e+pap1oYcjYVeYBp71I9rP9SCMV+sC42gL607TLjs7U/9QBDkDRo67mKu6fnjO11avK6Abk/k8n/
ty2lFEfz4L9bN2nrijoZCjUglyvK0Q1Bl7cEffYeK6K61po2d8Skb2Zkn2pRJF1cfG06DBfeeuDg
vRYjmNxO81Df5dijM2onvz8FG/7+0SUUBI/zV5DDYHl8prDmUMHyQmi7ik0GqlUEW0lmhxZOUxqF
VA0jkJ5iDtwJfOE/hFtJiBr6yKA1xBBDJYxN/AGjydwzLARgU6Ay2DA81GBHcVpoltFVupN8qiPu
uLaBb5+hhe3xGU3HFqUqAXd6kTNW77GZNYptg6uG8wEr1qMzoiv4gI03rpQeWsQw3BKxdUelq7eI
kk55CMphP4cKMtlc0RR+xO3U9VshRM6arw5kxYbYHCP3qaAoFKmSzabVovtuaEzpABSkZcg83KZB
ZrLL0ww9TN2h5dylQqcgeKrA4Sz3tzF4azl+VSOO5WyA4HB4YrsRx1hMUkWoR/ja4k+qq4o9SQdK
fi5f0CTNA10teC+YXPYb7DoA2s2qWJt79I90gK48/mIqf5PkBlVqnWVJ5V6UbR953sLdJA4VF/Qy
FH5UkkRu3a59Hfb6u7s1yGGxUgpLNGGwZUJckpGR6aDLSfyyEoXhuktYEdSv08kGKRR170omPaFP
OLmjrrBZcM8Dv3QmzrhxncyWYLxy+ICA0IlHawyAC9XrnPNz9aE0R/2LsoV8/JpNL29TVEbZ6oOX
XLJMOawVxw9e2SE5bcg3rfBu9tBniB64ni2hAgXoq/xnT5QWOrAgi2qhLX2BDXn9Z6ZJWTA86sLI
q68pLkZZGfPV5XaMdRBqvkqhVqLU8u0Dq3RoBK2Uv7rAdkwyGMreBvca8uWdaUCOJ5owVgaAHdo8
rFRtBYJfMuhOh4hU/6Q8ySg0BPyXLIbd2U3/qAoEmAO9xJWajVTTH1Nju/DaSFdjDVvyDPp/aLbc
K0T7xJGjkfgqpLT7NE8eJlh/DjrART6f8bI6bX3V7JJ6kaOdAAS8dZADFeRRF9rucqL8A9L/Afs8
J4YNJa+b8/PPWxYcPxWgpRrc2vnyXtVy/9+umDAMVrFYERRvRD1XCqQSUokGTziGwDrTgt2sMlpx
m2f72MNiW/Bt0V8Was55DgXqWlC0B1fbvRDyvmJxIqIXZ+3NcUOHumK654595IH7JuENI2IYd/vb
s6xavH+W/5T6MZWP7ZeeYyw8oS18HALNbxlYWSHm+1bjepwDRhe3GvrXD/XM4HEz9kBswty74w+c
UE54lJyMZ3ymZoFMuGkCSO1oyQK1HdBMiQ3abks4azMbhMUcgrMbCkBPvUMjKgVyMG2o8uFGsF1h
CnOLqpZg0IrcnqNabT+1ZPfVItRZr+MLPGw5UIOAia6fBg32BBRscRUfNXUCwuaPk6b0qPzhEHIy
BpKOrcYbOgHQT52Dz8PW9RG+ZABTCLg2RaeJ8obZOzONAcvE73l21+vpwQRvOWZeBX2XNLOJUbAl
tyH4zkALPxmWhXROrV8ObRArOx0/Cs2yO42rM5N4Fxb+nOaqNV6c5tOlFMfv+Yal5N/5O1qmvj+6
7yFOUDrO0OecpKw+IDRyImVzADUXG0pR/oC4gLVG88B/sKj/phCxYkkt5jUvYvgH0TGoRwf56lu8
gvt64XPMbPJL0fx1p9hXlnzExC6HbFEv1gZScUDjbYn/tt6vFkx9483o1JVoDVcEzyaV+jHcr8c+
dVguBnuFSOjbUoWt6nBdAw5CxQN9GXQEUzRRIIv9TiU8vc2Qefvz74+SxYPMdmVQ4t5B+e/R8Ggd
4Y9HgNYLr1yxDsUyI+y2fKBqPih/rLVgX+KYonIo9z1Td+YNGgTBHZbYH1l5zrVkhZ2dXD2BRpuQ
btZKm0sE0rDrZND/7lmYQW8UeMKtsQ6IgW1CHxQxk1f2FnEkLdrB4qTVzI8z3BCq58QwPlX77Bas
9UWJ0J7XD+5PxMNzEbCBPMTbqKann03vq01gHAM/SZECEe6n5F3jIZYItI2w8u9M7kWCfvp31t/I
huckSOP4OO9BbjWmqMjgVHDlUYlq9qSWQ1dCD4Kc18w6V5c3ifjVKmxlHQ/1Facso3khCGOYd1mB
/w5r+/AgXEJn4CD2UVbxuJ4j/Fs9e5kNNHJoHTQvFxdFyD3PusA1ubn0WVndngPALktdYfSqn7ng
AOoCUahkgZXzdKh5o+sQAH/NPdW0ZP/6wncsNbrXzz9UvT9NYUAyk02R2fViBqcm7aBn2YEAwsb5
gNDYShpXjroW6hDyKg41Q0qbQud3fYGGJeDS9Xhs/+Z1Z51/VRzIU81PY3mzAyNbrv1hg2OvGyNU
I1k16MlYBfAgGS8d2+dNvbYUauBi0q8a0xJi5K5P1t6dWevsuqR2rgAbd6CXtmItxExb6e2zxgog
mq8zzuoDjUOKt8gNZiKRFTf0OaK/e7Ar9yzMpSQyk2z5sjgNx2IAx2d43fB6+zzqDWZinrThEvxV
ebJnj8TwZ/b9aRYNTZjlZCzfkkm42GaDWqqtvMFpqmksLqxc7xJ/kfz1AkyrBMZgyOBrs66Xa0ai
Sb8DyWyVoCjfO+LLnRLUtiTABG5na8lrt2/wLfuTWriGjxVZ3yzxY0DX7lTsceIbMhE/pjD7ee8u
3Bgd2hIxzkRgmo5wQB4VKoGJ9eSPLZMUhwlQL31XxThLK/PbFjBfYegL89aEsB1/IJ054xOrGe4/
TzhkHHqjGiJNSWdsIzyPwr20L+63nimSQi7hmIeQNtkjwr3fvjVkldOue8INTC3qwBFDrFpIo3C0
LAK6z1M2rT/W3nTwUBXLmREgdsaeKgs6WpSyiF5zri6b4u/ozGKkYPwsOXQU7cGBIuKaZy1BjN9M
4QrJmtZUaavulZ5Ghn+tbMoP7WBN3oIX6e2L6TQOE5v6CIYwcdjPdC5Q5VpAI3gKvnst9/UzGBcE
Tgbys5IYd2OetoW9OFX3vJDJiFjJstrMCfOW72w20ZMsCVMcDYW+6u6GzXrRBZP0lbC5i7185gKv
l98nAEM0I22bVb/lKBCEaxFe2qE19DOfMgZGa/1jzKgEVOiTLNCBawHP3DhbgdR/4yrBFUMWSK+x
cIMaDLwI8ctRIXFbvrJcPoNyXAq08a19wQdgE79RdtcTasH1o/KrUGk4m0UYOCoDKEq/xCs5Ryr/
PGvc6bQ1vk2XOBoY1sSonMXvAgCRrAGGguGgpAAxMUaLK+/QjzR3Tis0WBkMjaN8c5g+BYNrC2Hn
8VU/JhdQaLQhHsp34eYK+pqG2FMC6PxRHZGAa5tnA+qSr38dq+Zxj4y5r9A6mSd5+fqiGK8boEHc
Uf4vyfgxnSOg0d72Ex7GlmSuzgpcLJ6a51x1quTc+UZwUz2mLDAMmXn9RDUD0mxMJC68XDG4UrfX
+4A+LcVz98+VICue7TkBxxGgxdSSVgXQDspc4ZYB+V3YCeuzapmNO72lqPjyUddk526lLgqYhrys
/Jjg3xM58K1C1+hh5+bHjVTjH6XpJpcdnJpgqrHunmdUqarDDv+QY9PWtluRlAq9O/NgioNqB1V1
zW8+DhrbBfLUQLJnl/96FgE94VQTPdCKyNCA/nf0Vo92jId5AiLdUR94HJlt5Jvz9mcXsgNd/lT4
t+WCjftt+gxmYw/xcn3wuvSs3yvJPFcphxeJ7tg94n9lz2pKb+W0GzDgT9UcqPcvoQc1PZ4Wxyf+
0Je+Kf4wvLbv4G7mfrXKOcX7lFwfVkf4xMkPc7up0hao24ClVfeJlZ7RyHUlm44aagRbB0Ugn8tz
93ZGJqzx499m5xvoIQd/H3yYExZUT2tABB2cXIrurLYz8gXF2N2vkOaxNao1f109MG8Jq6eHdhCP
k7FbP6An58eta64aTgbHR2cNRTWe69YBnkEz7WN0NNAUNl1VMo28nBxFr9hehFND+XWE2V51ddsc
by00lm80gF9/M8AoS2SkXDbPdcYx99hDp220f2r7flOEGVqUkoRgidd1AruHM1HP9rEo4uw8fXkr
ZJR01WEVtcXMB/z/oZPadNid6i/2V3Hld4IkMM/ovAUYtZCfXctBb6MHcIHcVaRjB/ATDGV/mkG9
D1OqFOLJn+9aCfGFftzrtq+Vhx0J8f3T/wqPpfZ7gVl/CzTbU6YTWXBDtA0cKxrtK61xRD4NJ9hH
PE1HjDL+vakf64us1hlv1tg7ji7HzTlUW1exOZoGC+MjTjIPSi0MagG+eot6Y+yBC/DN27q8/D+B
nj0PQXakTc4MFZXn1pR+uyGBZ33zJdA/o0jBSKIwqdksRTzUc8WRr8PxzRhWqfiQKKUWsTvwwBNO
NDLhBjjZrZ6OnAmKvMXskNiv1NLtkKVP56uTR/Hltx0QW6K4SnGwRfMACdpRwlQNnA3oR+B9MPVq
csyXTIdLJDIq000OMvx4GxOsvqyc+u/CQ/ip7qN0AU1NbUFStygzeurwikj8V4ubXEpOnOdseiXW
WQQvrWDmQ5yio6B/W7jaEYwTXZuuQWDgj/jRT/kVrZ62cJRfxkAYkuHqoqcwa1Bw9nqOonyCWaDm
dzA4s3YFw24OVxatKHc820fzHAApFkcbVKga3gwwnufd44dIntwMHIqIT2/ekQWWcPpMOllwOk/q
Tf/ik67HpwWui4MR9SotS1bTJCVhutlUaYii3n+2lyjNFiXKfQ66HiGAfFyQaxRqCgpCaKhW1emp
6MR9AENLw9nmf7Tvdyq/1dwjuydo7keq/RDjzUygz2NglfGTUw22qozl9Ei2HV7cJ/mSthMQiAt6
1IZccLTowChm5QrmGfH0h8dSFTexo4ck0i11PC/R3XbITbdAL61rHegICSaQxVlY6ZI2RMUUaUKa
XvzI1ZT8493gs5ow1iYTNFFF+zL5Ka8xJQKFXj0+aKWg0ee0qWNboNsJx/immCNZCKBG53Kz0MzS
ShUDsaduTzPuqrlwWLeaeEo51vL87QEnC77TrqP2P2cKLssToGgkzqtB/f/Oj6c8gOrQLP55EwCa
s8o4DizhC9LkvMxiDxUA1OPpxsnir2ZpyzveVxwThY3TqhHln3f8fORlfiYTsFv4QTlwnax929Qb
DshJH7rTkojO8NFDQwIYlzgGFABTdKh3848kor3namXEPWw2hj+ZqNILIjQEH7OUuzbl95U5fuce
D3Jf8RrIO36xpNIkuC0Em7hsgvVh2H/C6y7WYUTvBbB8DB8KjRPxZy+TAGMjmVY7c+lrCVF7FHV8
P7+0B5lK84szrW6Kp5J6wseFJ3iJyDTWfOCQlR110FYqWOHrETRO8sHpVW3Pyga2/UVaNBJDG6mK
/0PY3Qbshmsza69rncmUUF99cVtBdTkz73wrceeip+WmPWMuQVl7tCSsb9m7tOp+fz7Rqs5NUmsy
0+bPddDoupWQJpiXom6/L3kZvR2uXMT9X9WNZuEulKZbZpzpa7hqYEEJExkksiSHbbugueumnBAK
cE6+7yzGLQZftWlZ68KntBmuDpG12BCLPGCK2OdjrKI2qhnU4n19ABAsmVbQo/Ph5fpOAGQiL23f
uSV5rfUt2FdWKOaZgIj7S50HbIZf77vkt21AeW6DCevj+DIZWYtQWpJnoat0P+ToIiowURn4qGxu
ZWE0ImIgNJtOOXNDGlfuMaxpLzyjYqQR2vFIlbYl+Ni2Tk/89qqABemxPZGRGMkikfpFPVnh0vKC
yhihBqqHkG+uf1oi5u/TGJi1lNJ4jTra3tQJhsBqVYjaaifuJ4RfcUP72KjtEw4akiljnZ/oahAD
FVs+Cw/VLcFgAJnWIkv3M2CivqjXJQdU/OD5cqP4CWulIQTDATi7Jgu84trhyEtZc2Rh6wVcn2PH
Mhzc+TLeNYEChlyWbij2GhPRQZIKftD9J1/EZQXOjpoY2sMMYVYOLPMHUT8U/siQzFBQl4Fz6kYZ
QIRwXHBKO98CPebStBbVY5Or6BwAUjsYCSk0mMkRLKj0hee3TrZ2Qtsz05HeaH5GCd0vaXRA2yNL
++UQrWssdG071g4+Jjvl1QvJa1G9Xul9BxbL5B7SOYr9Ovx+SD10ZnjgrhEuWYE8rvrO7sbjYxmL
ZsO3lEBR/zqXy1Yzz5IhDABTF4CAdyZvrALsDu+Nx5Q/2MWyje0GupJOvNg8kzG2UqVHLlu8sRfc
GokMscbGAh7VcfgXp2t7SihXXij2uJ6Vbnz7a4Ok+lPfkfoYCGxUP7obS7VICIlj/WMb1lxUCoRn
KV8fNI1XZHQaXPr/oy5TBk73W9rpDjF9Ari1dk/2/kPIAsU+1zkFmWYDdf7WH+Ed7Mw9brVTel58
Q5R5GTdzsM8dWmhNzpI3v+EX/2xckDaEBZsB4VcQp3VHya8Dw52YQ/tmQQGwo9lFejyp/6NCvmJu
MDIFTIjGTAxhpLppECO9nQtKUUn73NLoez+PuAXL6A54eUx6yJ3DJlgis9gZ7D1lHocFv3w5e0WV
u7dNygc2MUDLGuZXQjW4a8ifrWo9Dylrq5zd3YMpb+5tpU+eqsx7xeyqYhmhbOUs7t3JsjEii+h6
nEzW4g+2HnUepGs06ShD8leWqFD6CBcMWBE0vzHzsXY0ZQT4qGoyysaq1WCpPhXI5QykMf0+qCwg
uk+e3Lh18Z3Av6HT+Fz02Tf0olhLkWeVvMNzyqg6QfdMwxOUVatdeB7mTHMwayuX34ub7aImEZdC
aAJo9YqPfNE2YcWkOMRaTRS52ql0zHI9uKN6IPCVU8/qeOaLLowhqzZF9tm03yLhQf9oq4VREXWa
z1oCvFSS3h6ysAs0XB7FsQNc+moyCUL4jDeUxdj07P0i4OLnR7y6v2TQnkp+D39GDIuqJijDNmiL
eEfZPfm1T4qIN6YHANLNtQQs7SSUfpt4RzX1ae3a4Q2bSeCEVffawIIuq71tTj+8IT+X6wDfcsJe
T69coVJJTMFRWJcSCVyhCkP8CGEEx+MtKlpdac7vVSNSObX/pv+iQ3BWXyN4GxIvOxwQFVsWlQQ7
IpJ5tWQTflILjI26VQ3uFsMJ7i6pTOBsskdeaE21QQ2nmNgpg4QEgK5XAMAO/+RF0uDMqniBxXx1
RgIOoD5acMRG8VnJV5UnlKifSLfHxflCsSlUfxdh2eeGQ81iqzq0A5I/wYy75NVY5IPSDdwkqAoy
rLrPcd3B4k8n6K0Dr0FpTFlKUSFnEbJGwnoMKL8RTvS3Xqbdp1BybbP9Z4vzbxlIQvD2XfHmPY/3
8nxKavUnt812jnZ/3VAKu09UEFrk8MloS7e2p6dTrFqL4CuBawFfWZHC5lG84jC5psdIEk6fXk9u
VfgBmn+hIXcnlh2aOU77NdrIArOEv88l2/OGPML+qrLNEiGqE91oV4mPllkRzsyUG9rNIpRzNKVq
XnqpDpAnZkCrsRY2xTio472mdBJWa7bQw9A3jFJoVnGtWVGXpZwIyCSM7qkILl1UcA8RadrSW7u3
q3sgclUi8LFMIveFAl/IlgdILCRVulu+5tf+RKUcZPLJLORWyjFT78ALWYyDqTbZecVCaemebhcc
WfYjgUKaitkPcrNzgwCsLlJ5W5TsFG1Cz3CCBsXZC/tfEJrB4sosL8jIu6NmcZ5pnNKNvpLGYcCR
6Hd4ydowReHqJGs7tGJ6aGRxdhyg1OVElDJ+GlsYdsatThG/VDD8S057ptJkl9Z8UITl/3NFbTPT
Q3cl+nn9qP0LTIntlz11B+PFLqq5TEFTfHz7YiV33UUsEHbdNWjFxhCl+NdC98ijKsGSALzVAS4g
IW1zlp/xBPt52Fq9JJNjAdLjnZkkXM4EwS58DOZaIaEhROvcrZBHkWnZnLWBtv5GyBilgQJea/Er
zc78mqAvdqUk6qB1tcqEaJfVVBNWZAkIf4SFMzhTjE1DwYJ8KUWI6KKvCAXK2REMPm7JpHvXlRBS
t9O/wDMBwNnzcN/cKz9hq+N5ZktcIIhKhoQN5/skvZyGFA5r6AEn8VZye3DN5lUHKS5Kfb6h5HvH
Ga/EKnL09/Gy9txJtTFTtfJIO97FrDiieyby6wF1yAmkLCHGowy/7SAPBQO+CJglr3vmOq5mnmT0
AQCRjem2Ool1TU8QuMBEI6PEC+JBX/SR/uj7EfwQbnWb7UX9/Vu+myrAboj0Uj361wcOBfx0sc88
oyduRtvO+4JfkTQoNXh/RhvhtxTDxPlXtisJ1KUWVBTL89MbCp3HKaGs4Jw0/nubz0KiEeB4tgSl
V7O7+m7ZaxSPETFCS9QdImGPpCNxXr4PO/YoLAoj3siOsUk/L4JF6CZev1q/9PFO8NUaFQuoHna2
Wo2O9bjbhPMLF51fCvOx9++W6FnvuY6cTz0y2xWybmFD+ojPvucNTliru+Hluts7g10iEGBC2mfF
COkB3ZDqV0OdKbOFv3Uw+kuPXvu/4IvZKA+M3oaLyS2fDhX+5M07fFlRuRTOxd5IaqEwTXfyasc7
CNzT1N979aaOz8tbn2CayBdsnShUlP3vDWHY+ZFfOxLOKk4nphE2GQ1k2RvtUcsLxZYVmdmzEi90
KjLhp382+42XhpA9vddynhsi0561/KWG8i6UJnJQiGe4cFjsIaylrPJeF910l3xXL7xcJZZiCA0L
L3lL/zpFyx3b/qZMd9OCYzgFn/dQxBdUnclpOOxCnFlyOYoZ0P3mAQqZajnDvPL3OW/F1zJzNoaX
P2JVF5kzi2X88BwccCcjygRox0t3agH707CQMwcb98nq/V7xXUW82/CX7/t+3V2w+BewYSXn3zfG
TpBrqKiTP9z1smf2zg+0g4TCmSgsObQzlyShVql94iHz+bN9eP4b+bnyWy3V2zyVJJcA7ZGXi/zG
9PXUkH38gJdolVflvxtuZsYCqc5fwhXKZOdHOrPhOT04HP8WbJO3dEyrCXOk/NUv1sAZ9Jr/amzF
vRhBgT+NgUYNfso+5Tppm/rxRLJT9vPtxk+0r6KSfNvWc+6V8t/NtJlH7wRKRWgYT/ozPiFHrwj5
uXclGLnmbLN/HzvQigWwrZaSQ7owc4usEntBPiZvP1GoJRf+/zygVvG3+2PIVNCZwWCBOGA2rZc0
tvwZGgVk9SsNBwwuuCePlHNwlg0vODqNwX5b61cf+s088qDBWHa1h8pwtwDZRrah3Kl/kW3Brif0
3vPv0RCCZEmqnW7D9h7PZiUo3sYZqYTL90wPqkGHmpE+oxF80kePq4FcYPmBG6jJCDQA34iN6dqK
pGfaN09d2J6qlx0a9PYPzLmn0ZmDuiG3XgA2qmU4fIxg8uOPPdtUCSbNiP2Jf2JHwD5yl6rOZuxb
/6YCmF9fXHHPCvQlRNm2WOpn+ajBDZhgztg/Nfd/p/yhq5/FdtuxYpVmFXFrbCpRN7SJou/XwIb5
qaaTYME4qDeB1dpRVDkyHucurOLasRHFtmGCSrppKW8H3qIaM48MLQw+FvNfw5yl4HickQ+ZvUdu
zrsqQIS3A9zaYx+ZZ+zFN/ACdeJ42BL/A9eckQ3w9W5P3bv1ezfjx2fknlqcJveaq4MukrVqUMMd
cggukzyhK4Z5rHU0E8fxo4u6+ZlzWQJ/exmw+8tChc7hpSXYNyM/Opu7BsTuSop1I1gqOP6M6CfM
7mvGH0ooPYbebqeEWqMf69gxidFSPJ16vInJV7YbbFUmceHDxREs/yvJESENrUvsQODtlR7+JP0l
0pZQRXGoFEpr6dzBYejRP+Qqe9XQE5LFzIboCGIZIoyStnKrM6agVYqV/efUkEVrGROmMh1SEEtZ
r+KBQmudYgO7gSqBU6wuV+xiAf5wjrmtdCiQXyEZLeA27ymtnafBt4vMNxGErRglA/K2+5M0b1UL
FUiIISxZTi7FBHDflNMIErhE7LxILY7OzVWBQksJFeD4bxq7B/r+mC1FjZR3xaRI9zYqtvOHGfJ+
6HzmMKhA8qTO/Yw+H9fMzResBSwLMcT63XBoGyHSx4uDek5NjAnfgJKoXID+BaIfVdZS7EH6mOQw
F8nKdmNZ3yFer/TYvE38zBS35ci8MUmFqS+zOQo10yopTP+5VgyRV+rWTx9U9vawxoZZDVKU4xj1
+W+/9LaYvyq2F3q2o0nNLphprX3bEuKr5sadOSjoZnh2CgS3ZfzgFG4nmywd95Pyz8ySoVave5HX
A/hHIJ9J2NPNIxUhzuUhVFIiOkQNcrfMK6Q7zpVuWTvJB6fhSoqw61cWRU/PHTIvNS1xT7Wvp/o5
XD0u98vDrRHzeEdfBM1Sk2Aj6QYrad23dVlH0U48pVZPD5CdEmu++sjvCXbWk8Nrrr7/Iyc1k/ne
KEXXtN9EYO+T1F7hxcvajTgfPpJ/CF9Bv9zs+LKxskp4913krwEVRSTqn9/3r5LSFCta0gTItxNs
vD7oqD63GYLTN9Dp+Wzrg8l7U9CrtHyldLQj5cphBgbBD1OinH5n77b9lqOHKvMyx2UId6YKl4lw
hF4XUaucO4Lrd7diIN+UFt0CnZhyGZ/cHOyjmVmgch7qKyOcgFnOHtBOt72bV+t350Us+MOy5lRF
iFsQ2nbErc63Yr2JB4n+YyXl/nECZe/Gynud/IQAtuwaPT080eq0NMa90X0F9Au9rBB7XMHyE8LI
8aJeTZuX14ztNUv41DIql0zzBLRDK1OCJoIDUKc4C73lDoE0HWZafjoaOayGkULHpz3l72wYmrrq
aQYviqGHMqMmL2lQGvah6/2NOjNghH9OsHZzCc29iOHSy5M8dQ2WYvls4ilGv1bfuIIcOEErXfw8
Yq/XOTAHrcHMFWLSnaggOzxlWTvbpTrTKwE9dnMk9NW38YsOg9pJJe60OrCrScgWUq/OZjMq3mSm
tFHRXkVzUUFARAW++B8NWLRURKp5A0dAtqZGMscUDdLQnCu/umfockxmQdMJgp6lN4KJr1VT9aR9
Ynh88qlWU5YPW69W/EoOoY5KTSVqrsfZz9ozKtV1btCItJ9EFRmq8X1xs+/f8pIK2p8b+dA8Wcew
JnpVa7QiIkzWQIqXzg3OzBakEZ9hUJyTL2UaMndek6oQT2MDDdVyX91R7XSpTtj35cZ3Cctt8mcK
KfOyHUA1BSv3puANYG8jv5pJezSd1gNFP7CawLKqhbHaHz8SFQGywbEcPfCGKB0BvtrW3Ut+z7gD
cpnwkHnEhYF7UhvFYquL838JjAV06+2+kWMSHsZb5T2jq4nFYS+SFdc1JlkGWgXrUkVZBymvL9Fp
bdSmUOJn+iJ4bMR4ijXm7vEjLefXbIcakZZjQmHQn9OQ0eIdAnqcdYhqstUb+iMMSLsq5JUDIpkO
6a7313DYfeGGqSX+MkSyEAsEJHl2mTq5JpVZGBDLwgeK7/If7RJOuvieWjauGS/PAHTy8h02Ujw6
ZkDwlVYeTuzXXW3m97jTAw6B0pThfzAVH5Tc3YlfocOLNhXO5hXMyK626N4KOnquEpSMtjvV4Cqk
IEhsPB7tQG/k7yoZhc4rRfLBe5Gdv/BqHNYTvPE6Efy74ni/r1XObdKSA0ALus8HIXMaB6poKmvd
qG863cJVJfcyG8lrEi7UZS2glheAOS1LNpMR8kCQk9GfkyjIa7P97Nn1XjuJhOi7iZKYkaySuUz/
g09dj6uChoLlqxwXu1HOrRcVSidxakdXLdjldfUkQHOiaxpsgvgOFGwlvl18jsiHnC59hgNWjAuC
C+ETmj+1IiTUZ7Da0YaK6rLHgvOal0UdnF+XjMUyp3FH2d7fVOPy4UyXjTfC/zcXsO9mE3fNHQaU
0q5m6mCDPgkvUEACU1VRDqdB95xh+rQSLZcIRc/lORRQ6/XGYXQxxEnn6EMaUoT0xjUe17BXNlSa
zrfDdSSJZYq4U+NwCvCO+wDfjWkCPaf+UMtLpPNWlHeKtvpf/lVKa9y2WRaQyxNdJ90FcDL9XSM9
OSM7Sf1G9wVJxj5gZuzRIu9R9H6vNw/nEH0Tj3dy+uvLT80CppADqFybMNWEISq38492gZfmCWvT
b6nEefI/0LrOBzrN9DPILQv8sknc5Yv+Bq+0r9pQHa8LLVjSf40dO38uh07YYIFQMwi6rbqiaowQ
Yup7vsk/K/CxJ/qgEKWsEfPuIaW6LcS4eqLV4GBspaeIOc38eaGZUC+JpmCUf/6UqiSwFqdj2t8N
TqctkZB2HS3aijGs8yT4ePqIE9TC65Vzy8UAXRw7NJxEdmzGv9l2GGe0lEQREgUj+iJjIDe9ukSg
gPs9o7edAFj/ygbxeWIf8rZcvqKZvAEmkyn9eU+4Gf68CtgSNnfQiCl2RUCs4YBXgA47inN3Ohc6
u6XAvUOyHuFI6wukQmx8wHabK9j7ZWNZs2f6jVGEJ71VDlJ9yyfYUspb20LSTFEwIKIudbPA3L/n
1Ex0CvvHqvKcTOhg3NT8ew/nr1TubbwYRWCbuWW2Xa4qx8g4zHbWv/8cY7GivdIXbLSZYLOJVtHN
ZdxeJ/N4GGnQQg1/zpWJyuVZdfwSEv8/P/hbhYAa5/wD6B0UROBstqkLJULf5HWujLKND3xKoQ6m
1kxfWva6NZgdkyj9uXz1X0H757wz33eH+L88T/oGmJ3BGlb+QMmpkLGC2RXEE0mrqPKYch+c8yFW
940NJKYssO71onFPc6BrHcRWiPT/zp68mix7vosAgw50KvlJY9BkCZlkOv9SjoXIiqyK3LyVmdhW
rPqOrKVASM9U69v3iB4f32Nf0hq3fJ4D9w0hsjhoQWIaWY8+c94akT5drUm/4tQQBamaNCjinQMk
/YnGpFUET4sp/NBGY3YQ30OWQie0gDYDcEa39mO854t870xlMJVQ69PrIxXdTP7oonuQj/C4Mupe
r+S9120rkMZC/SYUGrit8Q0oam943nHeOYMEp8vAySIgiUy0XQotZ3eun8n3DV/4p3TDBQOa8E37
L2OE8XFQqBKV8y9UYSk/00t7x9ia5vtZe5XS5KvXsTs+2ps/CdVW7S/AFy3LnOQFqmSKTEb2vEtM
KalX3JZMWuDkSuLBd3JSQdfzIzAbvx1USHbuPj2AUKX4nVLG+kbk4vXLDCsOUO84syoyR988CqlE
I6CxnZJV6ilESftyFUMTZNOeL+p9jwkqwPXcH9+Y698KTsQy4JFNWY5P3I/WXthFsB08OJehA78Q
86QbH3QUSdb+NTnmN4SfSdx2whH5WQgaNxCNvZv6A3+9IT/4izG7C6AbVpMVuj3onSkya9JjOcKm
XSSY8WIY9FYkyO+W4JRCOanhjDzwU2GZ6o9A9H9RGUBC/vDUWbMK4KaSy7CVem1gUzbWbh6frwDV
pLvIBiG7GLYhxIwME43bUzT4l6q9wstnXjQ3TymRtvYNjZsKILqwFEkiOVfbDaiB/CE1vSmbh9rl
WWd1lUH99YdLOfPgYe8cxirMXvIy2lyeOqdcuEygQk0p10qe0dlPZks1GK3S04RIrQIiMvEOKYuS
ru/3yFljejRQW6qXy96bVorE+41P45JoYG4Gh3gq28jpuCG5+RC0ePAL8fwqazSWT4akSMC7w4tg
PGMrOrWnNm/5VvcU2w96+HdZ4f1ISWCrSM76cCPkeOFTOZ+3lqq4kKYCQ7ICdSXmgAg++lI37Q9f
AM/qMIc44gAWH8fYYphXEhhJXS1/YAwA2TszxF0SFhmY7Ecr14ReWshBj93IV+l7PD6OvqZv4Sia
vD6t7jOwytpgAaCK2JH4QvEEh/A6U0IjaEba2KkA3oqfuwarhcWcYRbG4XYmEelbaKrrpI8TQSd6
9h3u2CfpEqiW0bhnPutkZnc6c97eWa/lrLzPtk9yXEyaVjKjqDx7LajQuLpjZqPIaBsDwX36rkgn
Gz5te9fBALnq3X6ex+aetJegyA1jO+3ZTawTvO6oHwstYJLebIeSLEtheJUj5ZC0u4UHqqbMxZPm
yIZGezlzefiEWtegyhfwTmRzV2WoRsroO2FsuwqrYLp6L1D58xRxSQCzKwTYqEPTzVIlvlWj6iHa
2G2pKdVPqqMSPeVbATBhcBkB2WJtSBDEXfWyvUrH7HJc7IQyyH0D8Tuq5oRtQyYGaZoEsH/dZmak
mmsUB2X8Ip0O/Wjpy+8hGv7ynWIRw7+fETCCXKCZaeegMeoLUtRG6SmiBdwmdP9YZvM346bz30uA
DAIWVLIvkt8JZAgkY3LN7gmLpIT3t+CtQ8VRT4Any+FyMHBaTLKDm2zURRoQdJkE+3EtcQswW1Bo
RoOMSk5cAqK7ko0FsemTSYdJw6KBhLu1tB55A/33zayyMNsrkJ62wCPvBUNASJo7/ImT3z1oXvZ+
NSqwc8pw+uxB+m5ql0pCebk6Gx/MTMeLyYiIiXoppHog/xIyUOr25A49LcUawLesQRa4YM4p9rTt
Zur1/9fk7s+1yQPKngjQaVAEQjLlTZW7KOhk/XSTvLnvcmqjSV41oMsuxIXd2bUfGZGCtAirSEOT
f/zmqp5UPc+ueIe9aRq7bqxyZQC8bJ7Fn/XlU95XXGU4OO4zb9UbBtn0g+/wgowoXzSdxwVqyerd
Aort4VWX9GctgKmF0K+2P2RFaimVeahGPBZCWHnd3exmApNYL+jiL1ZeufKDyW5nMGQsJR5zuQG+
uddLae72UD9k061XQKccrfzU4NDjf+tiA4R/2KiJegOV4bBMNhU6SNeKZbnKnv8oskOL5hcTJfHf
8OHJUcM1O0Jghol+9UXhpiYmh5OcgARyV8e7okDOuFNUXjr4VisCwlaSB0EMp0I0AEm5HSagP9zN
s8oIlDTpaIptujfOiwjdki+ySjHKXT30sPDM9/GuIucFQA020uNxes77jXP00ILWQFnEJZpPYHA6
vjsghVEEKeiefnhM8hRDjlT5kp2fWnE3MXe/l9DGCqiviZjneUp2W95FJHX1K9WQLdOj8bkvNyRV
uY2qakyXvCSDIhC7M08M6irg0wB6+YWfuNKygKYzpaq52G7gcXJp6necpZv9JWsyKSAaAZ85bMt0
bgX9rxitZuZLs9AeG6XfNRcKctvCw7k491qwLzGE1d59B6Zp1GuT5x6A2CWzJ0mY+xtb1AYZAvad
g3D6ysf4hiKF91fmCIqmoA7DSQxeifaA5cjDC76r7IjD8he98jiuFUye/sEx5iuHFHM8Ig9ZT3vC
NM3MT6TXfFMxG1v/6ywvKBSjxmKb7U0Oe67aT67ikDvQnema56pkcskaTFMA49K0J5lNY+MAehZS
CUjnIipY0A1vKsUGtRM7f3lFFwQ1XAVHIv9sHMT1o0R6+vydUL/mbdVbwK1OItAXKFdk+h3bvDlG
D/LNbL/hpR+gnyoGHx3kStAvbFkME44pY0T02AkhDLnfbrydz9aZUnNCs4b2S7LyD9vCFNOiV5Hg
Se5K+huVsUv2N6qcshzm2mKz1SB+GhkcpYnQ7qsohArG1NS9vWRT5HGYsqj0eZb6Q9Dv/KqBIpgz
ugYN93AMKMQMyU5Sv/50j+2AhXjewThyFp99YdU7LTKVAgljrvmvi/ExDzkz0KRCJSOSh9m3SFMk
u58spHXjH5ikTS0+3ZRFUPMv9cdzDbyNtz714y4CaUAKRj8novgVklox9nPV4vKZbOndT//vdGcI
oDCjP2AsWnA9V9McnZdchf/xaG54EwSolG8jR7viEgXAZPzWHNdQG7Sa6zzvRdzSlFBT1otdXO5N
h3YcF8H9doebJHp9OrhtPb9KcFx0Gu2pfTFODFvgFndEhW6JvNyHAPFTApwhNMrALmpF9Y3jwbyR
6Yx0MJ5gFTv8mEqOsyT0VJVqG29+9BmsD/DUmw8OpjmqyBurGm7BmkbHt+Gr/B6+MQQ0S8lLQzL1
s0ADVqk1Jvacy00lwSmLbIlMaRhoR1ea0JtNVTC39gD2SQjmYfbqIP+SkdDyEvRzavNxBMXoVxlH
sEEcFloTjUd4C7RMiB2+8vWOVuebps4oDboOICScVLDHMptk4ptuFQYkJMHtVSglo0vUiSpXdNVw
0xIuHTVh8x1jsuNWh0fa+dHXOTBCXAHU7viaWv1z6Z6dkxAT2fbPLQLqDiBqkGqJhxVAljUNW4nk
JQv1pkVXJNDVbm/Bv6CeJw7QBXZNysP0cmgOcFvOOdpgaxpJzMrexibF5UCSJdl3LSDwEsmpcrl7
rdInDfRbtuiTx/U6ahVeghoo/h159r8yXJ4yv+CUGXaYzdkx4Mk7L3eD+/9WFdxED2rKHwPtK1yK
k3zT5Sq2aHy/gQ6hv0gSA3cmw4Us8WmChNE+BqECiFqpLeF+IYK8htEaMjw3yr17TMM6yCXvM5iO
gTN1dho8k6cSznCiFVoaEIrrYiXfGXo8petXXYptg207nKxpoj87SDqBA/npCtzCLDzJ83L+13E3
fEuTxOgA9QozMF1J30OLs4jNK9ggnQZ+wRs/WH0dmSwvlttedzzLcXuhvHKgK+PuqzaAUvKNEtv6
9JehkAGgxm8HwSd4ODDhf/c9V87Ho/Vbx+PtbGNueAVuBqSafslAZSY927/LNuLsRgxT+phH5o8h
CVbUpGUE66Ye12eglZ1THsmWEFtujJtKH58BLSVeRBmc8Vr/94202Mst2shXNXHKW6bAQWc7XRgE
QV67KUSoqvRI6GsPk2yKQDhpZWbke95hBe7uPt+hCvyHIo8wlmP8H10ixPI7h1ss6Z4shZd0O6G9
8i6DC3TxMF/lBKZqvAwG4UE/bmgMd9O1tuC3MLH44aVTsiLGGyZgpzEeTYwxrzBCiNvtSQggExfC
qUMRviB9Bpfvr8OfGBYp3dqpkd4yZ+pDReHd0JK9DZ5ZEQqO5p9TRF3dXOGGAXBgQBZMgE0k6Ci8
xHN2FUQE+4cyKd/5inQ9oxOsd1uxz0+nuUxNk1tsr9PD2l10IzyNSolqqkM+Tykqmy1xJSi46xq5
K9INunbb2UgfROR9+xsRdXSA2wLcBFe0DTkPDd0dPQxWPcbw3n1iIE/6Cw/uEtZm8s8gY21af8Xo
YmJsBoxRsnkIjC7CF/LGurEEwdQP16kyOytnkARdgA0ZrI9MXn83VpL0EnJTTWWrnjshMjRMg8dE
J+ZI43VQdCH9gc0YjqGMcuuxNYrj3LamYNBXo91CXJe3Bicsv/Z9UfebDgmw8crlcwiAOAS+pN4o
Vp3Y58hMjIOCm5P6xtKUkcNxBivnpE/8rlq3esLXqXyNq3clUWZitU3m4DKG8Qs8LYShPzPMIC72
j7H94kfpg9W9vZ3Ndkbd85canLyN9nMzZ8Q812qRhASoQWRCHbBOjnbUPo/z1VWMV8Z896XIPYTM
BteAdG7StE5aBFUgX1MN8kD0T6SkiWQ4+zO8LYMdI3QNNhReSzEGV/I4ILMMqaFRmQ1RBYktM8lx
HeNBsQm+g7qBEq1Lk5unBwePqbFr0zQP/+PE6D7G/K8q4Ht62LAtMOHsVa1vx3d34E5O9o5aOxFN
1mf80if8RDZZDUMAfra9c5bdOldoIbLffrZadZXwt1LY86Q0tuZTjCgf87mGPi+6snAm2inNwFji
VmxR+sPA6ukV/jmdF8tkKZmdQtXJgKsV0u7p6RZ21YKD1Qz6QCc2rNufQWAhx63KA0Y/VOWtetz5
bnsi8V8SfEhIjwMgfCu66WkSw7JBk9IJZvWOuo6xAlGLnlrTIk/r0mAherV/joM1jawqWIQSyfsb
/5aiRSZL7E41k7LBMseu8m6q47yLL6ygN1K53mNd+afg5ViKVIbrRMfFwaH6ihduul7+0z/COmKf
MJ1sy0fest9Hkorhf4kKFrRKtLwFqpAMenBdzqrMXJTc3W+6qv0+ru3YrU95SriII9jYUN/l9Iw4
yMaes61Yd4+f8AHLiN2dUPVZW1BNScaJP5bi8bJZHJG71uzJSE8672OZJTuEfcg6i7Gj2IyTow9l
8pwIbsyYruOml0l/Ftyib/dev3oKH0ZVF02ZaR4OBKocmaoMwPs4RoFmBTu6DOtRxtRsB+DI0wwB
BWH2xyTiXETsoiqj4XAYBxq9J5vMrprzxDUK4pO8zf9sokgRBNURDnk+V7Co0E87LbVaeJVq9HHC
34RnJhQGlWGxKytXoWcLu8jEB2q6Scal5+DoDNDZfnmNIheO5YiRZJTFmMLX5w+n4qLhzaWfzCbr
XGzJY89wuozVgT8n0dEOpMtAzIrDzOdwzKsE0L2OpeBQdb7KuXWRYduuvxfsmXxNm8sa1Cxo0MUC
rTkknUu887W78JGqaRkEgyM90YPONzF1TFJDeIWPLAcFw+rRCEAv0eoSLuV24hyD2Wqa2yjIunSh
0BKT2AI4Er2YOuDCNmR9re+G1QsLG+9sxFdNhAwQI5RolX6x0vyPKFpiufMsXR4v4xow6fPa4MiH
BYxQJozYnpDHNea6NutEjUkDkFVMEDqwntygoTBItwyzxKK6a0zADF8jbZ2wgWrZiEkuUN0EjhuK
/AUMEqj7R/YmLwvw6rn3tNhJOkAMKGC0K35gwGLJrlrNDbplm/tlBmIqHsK3LMZ+pdKRObZkdQXl
dPPzmzczQKsg1Uj44jQB5bJZrT+0uq4B2mMIPDjt/TGMc2+y0/cMd5y6PBtWVX0/9cqgKa1fdkEN
jsRQhLuOdJBPn3Gu7NlGfTG4jGxB1CEJQw6cOK2eurTuC07UzUYcW8RAsqq267GZMpx0PM6HfSio
KhYFh+imMkOVP2Vi0ZQYMNUe+go2KM2L9b7vvAfxn1vq7xBmol7pCfzFyqUs4d6i+cm+I4fcBJq7
YD+FQWRwtrSMdYUJPJJa5GSyXmz7fUgOihiQNlsV01AEuPiOxczIaeXHjECK2EHR+FoCqww8uICg
4dRb5/1b1zVQHmd8unyola3PYMtrBAtWqVm0IfTZV/Kfku3M04LsjhuU2WxDZXMr3d48JyZiN736
o9Nfxs6jn8GJUQUXwx3aQUk2SMsCGHtF/9pGXuzZmI4/SNlqjSSktP1dAtwEOnAVA09bi9+Zv2nj
zMhHiYT5JqqNr1Xu9LjoTSXFiOp0wO8tvMPSuN2wRTm97qeqeGuYjnTsNocgnxYZGoh16IL6Oe7n
wPQ1nw7WK88ZKh3B8/bOlSG04D8Dvy3yUVcBmKvRcy7PqR1gmQGyBWlCBMkifANLQuXO1c/zFqgQ
ccJRSKr7QyQU82DM9i7a6Eq0rPxSsvEymxHNkUlAsfHfBEZx64Siearwwtf7myaOVcOy19UEpTHL
qGq+Dx+4iSPYERVG1XozlR+HbFSlJRho1+FqnGl74bDtPma3DxhdW7OFQwigsQIzTx1ivpsA4FQT
wJwkWQIlxZ0Hl+2JGQJrJ9gClzMlz9GgfNmfkXFZhPuZMPmcESfpOrmgbWKVFe9ImLSjTwvkW4ag
EOmjaeSWoYo/CEcOxa0Y3A8ti0nXo7NAcTaQIcV0+gcAC9o0M+O2ZqNFS/auelku6r7mGgO8rBSI
UuwRb+brXAjd+EG3FHleyOMD1MG37sGkwUT8MV7FslETxETHegDdLPknrXJZc6mXBzeCnxX0sH+6
wAYaemMbbEXIgxsxne2d743BzYtkIkA7u4Muls3fjeqoIXQzgp+Y93MaUfj/Kbjvmuc45wJE6YD6
04mLfMmsThdpr+nAwMNlsGePBv+83/xyz5PZDKUi/fRq07GhDaONeJBEFplLd3VHSZz+zI8QdHCL
DCJzWJr5/+Zy2amF8D5JOKmOtKfKUZ0rWJDYGwp7x//Kix/X2lih0AMl6WN8LdIWmeD7RALg/FpH
H9iqknRvkxyguWeJ1xaGjMrkglFPEYZHCkH7cvjAvz7GMIjaEbrPY5nKobnt9dUA+mtktyZNTmBR
cSZXj/lJGfi8RFwZPjGhO3ujSDkY6Q0aFVXOeymCiABhTvLJv8ZUEXDTPPKdDEntF6W9pD49WAbb
OkoyJnXEHxBjCkhG4RVTPIMnsrVAOODPw+znisNZBO3lcLyKZFUOzc4I8x1kbq48MSVqYLIxUYmD
z+SCdUdZKw6DoeasdTs67hJj9A2YxR3M+SYxbLC13I74aXALJIeLaKY6veSA19J0vNrlEV2skG01
qJFO8yz/jO79MldJNFyFWsuxfk9M/CUQyxHCzWLU8AaCYKhLfXi4DlCQkgdltOhGW6ip3GoWI0xj
tq7C2qJhY0x1Y00gKqSXTJxMiCGJfB8myoNNb0pETOydlfttR/wbPKw5SwLDYvUAfsAH0bB747YW
0/ili/89GBHNjxexzlKGxiOUbuIs9vR9ufBplVA56URaiW5hqBB6JSxJvujEVGRWPMb9jih/4kE9
13Nk/Z2gvX23UeRuGabWCPErw6UiKV8TcKsEBgfpuXPS/L0ih9tuhDNfCRAHh3gGzJzB7vbTNNVy
ttLvB6TEcW8ARQmR4xcZdm2bzCjcGuTcy6AGHGFf1X2lkovT+sfWi2vYzLJwGGH0QNbvwb4Q747O
SRFA+cHfP5qrYaPWZkKpVjew056F9d16L3N2MwKasDu0NJuhhIsuxlebmRF86fxEOBPQXmJRTw9x
qyV1tV8W9507U31pemHLRT0Pm0htNTkSUKCJvOU2xdAe9pqAdcEyrtzApi8HXGrCbfXEyhAaD6sM
2Oq5NAJrJhm+BSYPvutuSppxibWlz4xS7NeDa+zlp07jMIHS8W2z4jTy/ZrN4Ua8OjdqZeqmoVYV
wa8aJmL23hF7o6Cs3cfxumzILwjxQy1WK3WDlhh1XG89KFUZ8dYjXlO8l0FdR0chYn2umM0sZI+H
+pcHHcHzJaz2LRelm210FUt3VBQ9Uuqwmiwho57pfuX2hMea1DIMT1722G7kDhXRzAGExfEmTLGq
InwhWQcgkWmVxUIxAPc1ajAP3f3OhjXBb+RkpSZiXypPPXGvU7DbIMWZcoDCVVC/124krII0esdq
0IIX+wv0nJMkGOniR0EL1PudahCm8gDlegCCC4UrG/Y3YkoKytPyDkgPdPiBHenljkzzf0BZi80M
ijSyR3PedCppbBsW27WMzx3kgjLk11Da9egQ8uNH9nbklcWEbOVHauNqpeaDwdGtLm1mF84hGc8+
KWUS/iRNsYdxhcfswTH18dy5MSMlrh35IFmmxcFa9SN7WFrGEeiRovuhib0SCclhKGChzyMCL0Bw
o+mVGtXMh/DAIT8oYFpOxIjCREwcnjX+6HuAIHLhUdHukDUm8ubY4TRH0Hyv4D1fU/fLN6jU/8ts
FPzyx+8YEsZOWOzCNVQWiAErWk7gZMIGXIlRdJiJlt1U1dojKmMuty5vGSUXVS8Z/Ied1nJxwKTG
GkuQIZwS/KcdtnJQpmogUK0h/YiSOME+WVa+chcSLk7Ap3hFylBgIaWnxlPsQupFJmRKFofFcPN5
B42OA5Ur4M16oxbLhx3lfa8LFVo/wtRUNENyanhMiOagJNmO+D/cXsJ+URFwwhFm+i50nKTFLlsk
3sT/OR/tQyOKnwSBdNXRlZ68yd7uBM6bGi/x3bV2UBMAORfc1d7HrQflwbW0zQ5wZbULaTH64ZFv
rKbTEz8SmstDgpX9xsjlF/DE8/FTYdHLH2mJ1bsGvtictE6h97kmCOl7n1HKXR1MwBTXOc70ihPD
BqG70gaZ+EtMMAnQaaie07PIrP6HxNctuL2l8eIj+vtTp3ktWT5I7N19oo/KTQe0x7qW4FjARPLb
UwHLfxIr8gVlhAZBiU502l2iWW78z0dyW9dXFKnUnmQSJOA2PolWeECaMyxiD3t72Xn+8lnGz1Zj
i+CADZAjznRSQnFU0tLLJQxeptdG5nK9aG9l2wESYfVngsyAIRcthO8VX4TmQ7eI0gq06Ymtt6M8
yXDOemBv/qUvI8MjR+AV5/MXJuIw4zyjwDrVuskiCOScACCIO9VfdPWXs0mmxlN8NyNrcwHYiY7H
vD3lFFhztvVFzDXbgzWSOkvQFuLpbNCEBURoXdupphZiSB3Cn8elxvKXy2pjOtFYQwgMZn4qMwy8
CsY5Vx96Jhzoh6Q1hsfK+itYTLgJ1HSeqLZNxtgkxeIavTla5jfEaA3jiXDuQPYbDxgrJrlZ6xXm
GjbRKNPbJ9QLJoPV+q31A4HBzETLvvqq9/FTUiPpbMSBg6ysUA63J7TTjBempjghuq9/MGC8eCEC
fzL2TSlyuD/71VvjJ4mPZY4PPtilWSPux5jqQECdrLA1smsDd+zPCkhzsBlYd0RJmcypnICrjEvP
TaEL2Uo1cCeDeqd1Mbk+cxfQuK2iBaCduV1u3yzJ9ZAVt3m4kXVQuyskrHaDNXDWbF2xIHHgSIuf
LMoHSUOrnzrgRGLrs2zIvIgQstc4WfyFjvnHDo/pja6mTJnmNQCOa8YkdRHMdZks/vDa1vWedP08
kNSG5/bCAw8hKNz8VXAHvMqr3g1lhcje6Um9zjhuJfa8hja1/0C4wpTJ+OMkjq5OEhWt+11zEojw
O2Ij1pMs52pBB4EsM1W/4tZG2VRMlQaoruVF8rBdrh2dYqvse88cV1ZDrhfrJN1gykAx6PTd/hsW
h2JdEgm0wUY55FvRGlEaInyoX8MQFddvajrGY4IcO6o238ULk5aRkqu7rdzSakhSe5MVNY58MGb7
Aiq5l75INtaKDjw2uW88ImM/8SVxyL0Bq5ABaxPSF4gZVMAF1CKq2phCw1DMT2XpBM71RZRcKjP3
2WhjZEJ9yNgDOIxVyFsMGgloRWxZK+u9kxjia/1RJaleFWaGfgWO/SBu4jS0G6eiz8NQ/2bAqnrr
aIhf48zNe5Qi/ztzU213hkfv58mJ6w56x5730GpnwRuxhJsASzKB1xJ0oMJm+4foPTKPfVO/Fp/S
Tz6HL2UA//KmY2Of8SyqMAsaHyKm8Vqjsq26MhrMQ8Cfu6CimaplOeLIxzHj1R5cqkzDfPiMW50g
N6kIzvtfQ2TLKFs+2/zfpa6tkEcE288Lg7RIKGfA8xE1V0sRzO94dgDO5czOajTF1rMzAf9eHJLP
ekoOfqQ75OMcjvAd3gqoEJZIhwRCbefxlcQmqa3ugP3U2KH9OROhGtXA5do7+u0cqLkIMct0MpbX
ccqw5BIXBiyXFjucat4KNa9ewTMzpNXgcwTL8IjSt4LFha2iOHSL509ZhwQ6ckTrDXGnto41lqRW
bPhEXctdbYtcqsjDxmdbYsLA44MkGVKD39iqahjiIXcYDacbUPdVTeR2uVRP0L7+37yYcD3IvV4K
RIfAOkWRHbLnHnLmLhHodKBoHgugdu2IUKIE9d1eqFRMojDKHPp6HdAcIs2RAcYq8dgZlTkYMtZW
68ktMLFw8HG4qk4p4OeFF/TB3hC96CB3dBb9dLPv735lHFCl4tivQNus3zlbzJlOjdBhaXmcdx6J
rxHwKq1DdxbA9DhNQ0+c712NZMAfxG3A37SphtcgTEBwx3ihkvR6dqk0fd57qasRn4DuSWDEWsbM
zMNbIumE2C53jtOYnX2urOb5rPJrDCSJmargx5iJXEtSnqJvi+Fp9lG7SkIR+7JwScD6cFMsmLHz
mmRDjpzSL2nM0XyYb6dTztp5s/5n2f5OYteJH+en3DO/HIE4xoivSmp3iscyOxT7VFQCUMdimye8
NTxEOTOs+j4H5rTvVLQxDUPovAPBmzjhSSkn9NWvvlO05hdyjrjGPqTWSWSr6vkEs/PAYHHcGyhX
ql5CsSZhCNZn5xClslCsp+b/utkPxFwOt0I1VIn3OlF2t+SmObg9++SNj778ha8JOk2idPm00PQY
Y2tZOKSomDEs2H92zWN0gDPhP3ZcIP5fYc64EhNdUMBwr5XQl2dE1qX7RQVeXQzR6JDLktzqYX+4
v5Z/doVI7w5EWlDx6Xt3l6rZ+NW03QCXhUivBDF+IFcNIWZG36/kptDin0k6yUORhOew9Zb9v+9x
ZiQIR63DiybXLai1BPx7qEeJjNXvLvyWG9o3i2Ii0NE1WNZl7r5gqbiTySwzzZcx11JTk/MRxp7I
2zlcJqkR+s8uh4NBGCBxJ/jNrcAux721Vxj1I3IryQFBMLc0sTrO/CztcvgIlAtvFDU5Si+O4QoB
ypj/oofOXu7tKcLN47WOsWM0QfKgCbV2kUpnOzATn41vBUfQbJOwyvZe2rxlpCX0f99VdA5mTOag
glqwR4PHr0H2Fan11iyuUY1fBsNFJa3+RjXMrj28j5oMyvq6jsO9Sz8747FMjgRx/2GIm1Yxvfx3
WaUELs51suMNeq+fRfUGnLuHiAvsskz6EDo+AuOs1jX8Anb3ot3sarspBvlQ97NSoiDywUBDu1bj
2w5f4nK5ksU27Q8FugeVPCiv1VrIgoNwBJzMNDrgfrqq1SGScPYN1rPkHch6QlKgCvBxmv+xzRep
58+YLP57yRWNndgzbacSJtG8E8vxbA96NzkgOf2oD4ze5sn76TteLg+in+cvGlpKMZ4mitDRJ7kk
z0JV0kSV+CV86gylNEDz+Rc3yaaYAqH+9rXkSXqQ02w0XfI79/D3hIsyjor8ITEY/vllqyEMZaZH
5tfQifixOAvP3gF4CvDjJSEj6J5FOqUi/zKFRYu18MIJoy0J2z+KaDgqpfppPzGxH+elY26QPCv0
OKOTFzNjT/Cgs+fb3ArEmN6VMa9FlfpdsziPWe5HBaInBBZdLlVr42b+GhLRc0YaLe2EpWEaqQHD
Dj/8cmDpZsjUvuMRpd6nErrj1t6onwI+W1SKE+SZCi12IWM+ATTuVfq4xDJq9YI4QBqzzUcXjACv
dccWWoymT7ehWf4kXWQnQk1AKxlARhPzsqdxzlyZE7EqNUFIw5m843M4PCOhpnVawQoGLkURejyS
gi1+vN98vexoTOS+6R/ez+A1pz8P3fswgoNHi71Pal0ByRUQYOwFZWgPb22OmBx8cIPkASTj9EdN
/LBeJoa9gz7ROto7QGwFHnb45NDXgyQc96d9W/b3ZBVkNaOLC27USreFplActF1viBYyzJdMYLvj
/ebEXwG2iyyGfJb2iz9ofULyyThWNsYbozS+f3OvXLbJqCUERLLXR2han+ck1VZ2Dap9ZPaz1UAr
vzZriDoBYeJe4Pl6baKYw12CC6w69yVQSxEGaUtdLsB1fobTj4bbcRGwZwKyGHEdce9ZCWOQqj0j
Gwz3weVWRCrVe9EAXFgX79bT4BF3jAYn6yxerr8fIK/RT+5L2Izq3x+3365l6AUyVSFWY5ABvmo9
PE4ZcEDBrsSfHwod7sfMIFG/AcSAySctAWHt6zTYfpJNflApWdf0Ccw0CruQv4kdVKNli6IXQiww
sRgVQksd6yg499bwcNF9uewxkapkWayv8UYg9eq/T3uPUjgK51qDfs7nE3VN+3uovXwK/HOW8ovi
tzFB311+6F4IxCJf2HK/EMd+/7Co3Mbvt9tBLDyssh9fhO5SYELCC3vo0ebAq2PAcCVMuh77kBGF
RX1KTegMlTmGzusNgIjSD5gqRIuZOlh3xPJ+HTMALstRVszak1CMpoSdQyFo9S42s0K6bEzaGldx
leLi+7NjL80TMD5hL51x52wVhxEmJrYttjAy3BTq8SiZJ+QWm2LSpUeQltRuA319fqr1gad2C67P
iS19z1UGyPrq4mzi2ezY2w1UlZRAdJSEz+Q+HwfrbzWGVdo0Q//lWAOPJixBStrd6z/jPfY6MDaV
Io8S5f60NTTWAsH+gPzhYHHXTRNMh0yteBIfphprY54uVTOaTY/tj3BFLyLxpICjFTUaEfih1zlR
56zwkH+CtPnSsALtzUt05FKAFdRrUKuMpluxvX1GPpx2BwNVNjF9Ms4vfgDmF/4/HOojnDJ3kyqL
NICcjBnmDW54u2Rhs1IW1iVWRtYUXRxVSz5qV0hWAs3KPmj139vi2/x57q63jwYpnwuvcQMm9mLn
H7kuag5fxmlhR5yAdFvlTlWzoRPXP8HtVfaXyvRGHWO2s1HrEIUOGblnt7e9dTyaGpuVmxbhDNjr
cE5xH7pne7VMAyasDwtlmupgHlvBcYhK+q27qhmT9Fi+jKJ+jrhPNgNIMQq1CUCHHEUf5pSLGyS8
SUaIqMprn+nhCKRXoPN92gAMXE5ejcY3ki6CIy35RAxUNkn219+C14HSCaAbW7c3kr9uk3vdRIdp
pKX4D4kJvGG3+uyxdBHoUBUTJNsvq847wLj/qIivvPtx3peDc4HppRXvmHbm+2BJBOpJmLU25GRW
gygOSKmjXblrEVUr8zDbJCKyVfyPOtA3ZIM4W0KTo6eRQPeqkKcH2QNV6M0grwTAhq1hQhHyvCQE
8uXVQwwgL3639dFlQ+hTvO9cz6v3NDI7qpLXOBIs0IETElHORDbnsQdeLHzCH0fmZW+kH97NgtCr
46luw4IuZMMnxXZ4Ys8mf2GIyRuw3MtCQVdPJq6NsWJnLM3R95fclW9mXDNlieHXL5QLfjhRdNEx
P04g7buU+qaLFzNI8F3RU5/uMoaZv9zZmvbCByI6iVJ/2PdB+/gbsFqKAhOdvomgtRew+r7oH/J7
ID0k/UiSeRH4k8qqaQlwW2ACbzIRUWOIceRhVFOaXK8SuzKoUz5DJtk4zsUaD5MORlImsI1WAGoV
XjY/sAb8CFccQGhWbevTjZxl4rrNH27IUgRcJrTqwi+EzddY0mTGhQqVsXjMtiy2p06nHhWYLgTM
ZuKRBWSv/exr50wbkkmhgMDqOKBrmFklxNSYus2FjYwWvXfX84g3LWnVR510MdpD9gG0pdfvkZ4C
0+G1OqlRoBvt1Vrd9iXyyJJma2SAtLZFXD8AQNssUwK8CrtjI77XriQ/sc155lUr/0Z7z4sgiowN
zwMKHn4gHUTaVZ7SfpepyRLls7GV6Nfj2azA9eS74af7mAKqc6xHMa2bpb7qqjMA6xmPVVbUfZqs
6xZtvJp6z38c3YE0e/hQknQHZr90ONPRpMmMbSgzCMGvGtldQFb5jcczPKHLNcD0q3HCZdQEif5z
r+W3ApRF+PxpgeWWw1SsYj0eIOShnYh5aq/bfEmDV5I0uWS9693/HXU8ikGm0MHpekG0cSGW67xx
IUN0qYYjPdi4+xTXT79gj1er0HzaxKFwYZbMpXM+ydW6dqsW4ykdHhODe6nRj0e1ZhyObYTtWGqR
VmJz02A5CvyG1ENOw0pQpxdVfg5VxZpa9zCYDMj8DhCb1LrHndqP4BBIzAh9+9Lka/YziwXMZ2mv
qj1eFYnGLugSlptwhVt2FL4KK0p4tZ51o3gV0Cs45yKOFEkwnY3ZaF4lEjk6pmCkGCYBJepXwNPT
0Q8i5U/JL6B7T5ypPeKTvbA0QTc1SkFaBgx7yyrvZta3XzDFBE1uKOoueHdvYroMPxQVs0Z5N7hg
ySmJC5ItI6AMSBvmKk9kxq9aCBNI/vDlRGdMMob9InYKOoBJgetUjOvXc2cU7ONnoNwqv73N5lah
ZBwpk5OIhFc7r1jV6URiUNj3zIyp+L5BNevyreH6Q1y7eWuoiw1DKijJUMj3hJvDbKe1NdGM0f7Z
15hTXh3owXt3iNMViOU5Chd4PqiePuHOl+RNqYYi84ECdKqMTdPsmWodlJX9phtlVMwv3fTfIbuP
usCWpcnjjoQ24YQ0x73YmwwFgA3G7lmjT3l7bpnGj7rAyVSszqQJywOT1guYcOwWFieRSHmt5MRw
4QeV44MojBtG0CmfD6db5zibkdXFUdiRi5rizszMjufHM77EsKqiUq+CPwCxNyYt32icZLCDFwdI
xK2NrvTvjMX7LlKc7sdSWskHUjjX7ifvf9yr9b3+4Ach24mU38KfzG/OyqC3b3A5CNTjsYNTiNAv
eJ7E4Ey7r8M5xklmIveLV4L6wxkPmbf1iDmVwkP7OQpPVnTpoNyMWK++lmrWoOEvI7aBlmrgaJ/m
L2d7nSF+/RGFoJSYfdPokUbMpxEjfmbvQqaZfHJFAjbM3807wtmyDNCwnrE3KHy7dD2Q9u/Xs33i
D26F2mRYMiAGTnvmKufZ3G2j7MpMGxouHE2NMOvdnzYD3E4NgvdBBDKw5iCr8HS1NRuMtst/jnNv
IfWB6Y8kSptxKtVkF9i1+y/bWuzQ/IWYQk3LnEkgMeSb7Rbo3BBZOLgPoe50PnB/uYL9a11v4Bd6
TS9SzOUMkb8Un7TQ5XXobvPTSwRlcSa9B164fT2YPrt+uQcNRr5PSwaXa5fGXRuzsdQZcwUHP6v6
uJ5BhZ8IsSB0/BCGanxvmwh6I1tRxohGMpBDoecXQOukIVtOO53zl/rtyaC2TP8/uJbNcN2AHWAp
j+z8ezLidPpLVTiNIHrjLNte1ruC86YSB6+7y4XrDg/S9392ii9fJtTC96noohj7unhu5mGeLvUr
qhXABf7/W/e9hK4ShZ8/28sJp/LgXXPVUlRKKwpWNu+KoCqbSS5rwQp/IyzixLX1GE2N+UtDwvTz
89146U65fWJuJuYH1hpu5BcocEG+I5/Pvhcp403d4aXJjNDTUPwinsc3DCSEMbbBMTJwry+fTuhX
yQshQjT9Zg/qHERXjey02bsh57zp5DrDrJRTW3HBr2k6F6NYoS0zItd4LVmTV6+kN1ldxJnHKciu
VgUNcuzFx+0mZMG+Q9cG22yLG0gzBQrnq8081V2dHIxGtAQxBXcskru52zG4g6Q6oCpGl8DRfFhH
MZ2dqKxFe+MDf4qBc+cR3WNb60xIo8rNLVUf6fHfpDqoR7g320Wx+IQ2B4rn0I4R/Au673fo0w2a
28BCoa/i5iB6UgIO8o/0jAoxOV9PktX9RqCSAqgSvI4zwYwIwvqnGiDoeen0o8sXh+CA8c7wRbyO
FrT5GsXrq12zhMO6RXyQfMpHfHBMxjdgTsgtfhdF3y+CF1ZRyREZDIK9OpyTroOSQAdguJ/jCz4x
smRqr4+RSinTnAv6Hb1doDlBvUFXRrPQa9GfNKS8MboDHjrZ+iXRSWdmC2QSkcyEKYP7vC7pCPvc
qhUleaSBKG7eCv7TfLnMac5mwYjFMhzb5L1c57ZGAcakCd5RQvlF6aeevzMZS45lyCgH4JVf9ggi
r0yUW7Ypl8RznfR2DiuDcqmKAnbw/m4V+a8MB7S8A34ZmR0ZxrrBwZjckwA96llrgVOh4vWu9AKz
9xTiabpWb08bleOFjTtInb8bgjl+mTo5QB2DqsTa/UEENjlIQ3/nZhcNLkfGc9ijW9ReCmWWOhBG
cAaitD0XBhlpi3ZJXJwSxky+iNRKDyTxpbpDCzR0zbu7AJcA2zU1i5ElRkP7k03+3tv8VCF5wkye
WW6p8blukq3scN9HiDjIRXY/J53DcDVFTvYJ+ycejD/LUg9wRaTfhFQoU8kNd8g178iK9kbMNMtY
Tqbr3D7/yLFDavnpRNmhp7zlguf1VGhCVG8NgWv/JK1VjflHWJLD0vGVWuUwIPBwOMfYO+J+PSLQ
TlRdbGFmrPWENj3te0I+afa4e6ub8mhmv/Jr2OnOixD8UQsySoTDwOwv8byCcIXpjRqgqLXAOfgT
cjCshwVXHLxwKJlD3FigqWhPeSprHIYnlW64wtQmAk9iTuxfCVVBFX5PVv8sT/1LBxG/E2xYmVS3
33PsuWjinmROhN7UT3Oj98wYPrpDnQrsmxjy4mnrC+ufENa0EnuB4kQ7pKHYaqoODxr6/kzyIuzk
d5Gv11Bpzme3+bdKSaRFJpqnUyd2zNZNje6Y7FvrlUnddCHjkyCy6D/TNnfQHTvsIY9q05tjMYIy
QGuRUo/+ZNjkufViqtCrs03v4iN2fxxkiZhTn4bSRLT/DyqIKaoVkSYBWtW4Qa7Poi4iE3x6kZFv
ulZZA9UYa4sAe8Tqu845MTAMuVS22+lc7A/VYAO1NOTt7LRuvIOpAlujEG4Wt3pCrT8FPdaB1Dqd
q4LXeJ0aOuxoXKb7u1W2TAkExo8XJQqHUeloLhmNgi6ymq3wqFByFOrqYcok09fu4Exb+gFDMstk
Yr/LCU10FbQwU5DYDKhtQjaI58AuCrB9Tzmiu24Ue5MQu0dxk9BUObmRk7VMM8qg4jxCsfhbZnHQ
4ikRKc6bS3hRqvvKy+gdQkoWpm7YxgOsJF10AOAufbqg5JmbzesRm0kLwZbJatBHme4Ji5j5+yQ6
8Vp9MeMWTZGU1g6dl+wVVg2ssd6+XHl8K+/CNKlo/waDJKMZUpp4TrYsmaGVnrKP1evZQ5G4JEGN
lHtFjGSzyfXcUQPDL5t8zdFm4Mbp+cn7zBhnuDrXm1LUJpRaIebSyMvCYYCKCf0w83SNWiMhv7eS
aT0h9x/u0jiG2RITglFtMwCFcNV7q8ZETfk3MFmjmDhrFBiIIjKcTKed1uti9nB2IYypJTXriJVx
F/MUT+Z0fsJpS2PkVrDT7o70fJtQYEqQ2qAre+wn/LfHnINJ9X1gzM+oELlUMTwqPbOSFWiP5VKm
BoZB2X1L9tuIcFVIopIkC5OftSPe7ySNyOPiJwgpKw2Ktd2ONeiwFIY9W9SFyKJtYLdEAtlZul6L
9BAEZnPl1veQYvN89y67AJzFNHoU/PiksCIBYOBocULxD8xSLcMo+d3J/V8ETjhjiez+yTwlyAhf
qpEDySERr9448eT7Mwz/sx9H8f2Q/goMnhAZCiwVhoWj9TgUbOrIt/WYc3cGv36IcoLvX22edINl
a3XotHpafgugm9aJldHNnwGeRCGnRu0ZyTdvyfWGjcLqeDnvO9PdOcpxsjZJbg2m4xyKUoqRvnBn
EjR5QV5XHzfmzckGsGjMehgMCeeHrN54ZXuIIW8dGvLwuCpOzjbQx25GRINRJgtnOHuJvBz8Anfc
0PMqHNWyXhmkXDUYMPhSIhJN9Wkk6fW7YMtl/kPdUJkuG4/oKFWr4DligkDCVOvGKVS2egyqSwJn
1IFhKd9qI3Ocuoj/mrejG5isWjsS/iAr7ABj+4pRffuX8ihlEAnNlhsDQFdRf4JMh8qtZk749ciD
mwZYdHbRfQ38/QmPfjlarhUCmTK1BfaZfwZYqU784tdjf070hIaumjxYSHQJiDoObHOCVUys79IN
q7cn8vbdWyQdVIlZSuliQdvY9WVnbrvWwSIPNwhf2wI/CrbpdO+acn/y2HKbfLuAeyaSHnmnb2YO
bDDRBSRqIucyy9MUv0pTYhSv5kcK1i7asywOXzoRIcWTTHdZ1jgsdrznLqDQRXAT8TZJG29KFRce
jh4QGgZ3l6eSiZY3x1wmAGi5vnSoj3umwGvCCfgZ3d/btroSbK5kYRpLT5It+JgVyX/fuJGTfXet
cqIDFv6iop6+cYdKpHq8edQsHDQ+1rwVzaag889T/M4/x/O98kyhudgy09JxjzppBC0c4HT0Fwaa
PCKYm63mAS2kZ0tbszjMkJWn639l3KuoGK/czqHuHY5fl1MR7hagfwc8b+8YfDclFAI10zsYF500
EAfuzW+LrRX9ExWOVgI4K1SxssSl0LTFG35YAdFW8U5gLb/gae9Rdx2fhpQrPmUEysAc0wnBuHxd
7xArmFt0LHLDDD/5vlKI2jfRBoBM3mGoCRxPR0z+xXlgJ6sEwzsCRtLN7VPWxey8iyFzwaP8q7Xh
xQTr8iIV7VmkaQvFZ2TTAdJZQJ/lL1ujAjeHzaMD5VeJTT9i3v2JhdUWojZlEQdmZRA82nl7En4S
wny22orcCvYZrtcwcrqJvqjCxaPdTUy9nG+IgrOniSHB1LCy8CUXak60bbxRs9Pzdqw9eeFR24gu
2BCCpEICN/9yshn/e6BwKF3xST+YA3HvYmsALhugDskqvm8Pvxa9+bGevJRXNhTC35YlPdpDk/Bx
l0awIvUAm5V+tr0kk2sk6OuIncGlNRY2WncFm54p78l3//E3iaMuh4iOHqamC9WSRxLw+ZZKvxn+
C0YBw9LlfLzfcF501RLbpxDnkbUECv4ded5cYtvKuV4d4HQjqb5DFOW5sSkEDeG5rbfvmoAOthQ4
zdHytvQRL39CEORvLLFn5IN2aJESuo5bFTHih4EOU0CBS+X1G675HJxf7lASLSnI5V9/YJo8vdoO
dqCQ/1mnUe8dLKXu7lx+kW3TFKrzF2nU+mld3yo0tJP/idlNpkaIHPldDj/YIN5cxjdVPHoGvxUm
K6XIyFlslvNtNWm+RmobbQuJ0biYcfeU7y3AmlqzhiOIm6VXyy4JGggUbYjng+NKPIGa9eQjv5eq
1/SCzMkjTsJMQwF3dYk1ufXRCFEHJCr7F0RXvxAvaUMHbDLhi/0POhIWorA9P+xKblQjON4y4fMB
JvVDDqj/pDGIhFNxQMqNMsiqKIAAyjrofKuAvrL42CGQBrT0DFgO+T4mrOTqN9/2GTyIEnw5UBTF
BZggy+vw45Ac4aNGoLLsFrVMeGuCwJSPuV0fYelttO1AVtSL4q0XZM/3fLxYHarTszKHBUfxuvHj
Z+e63bS+bU227AlwFsYug2RnU8/MBDuYZOaRtSf0dk/GqLU/mLC3iw31IDUWA9iz1nGVeHVcsN77
fVWTrS1WO/lLu2/85wFEI0X/pONfpsrt5uVCfsjZDW61Qe/yFkuT8xHRKbH4wUDUoZbWOgpXARVQ
HODeTO3MNET/QxXQ5F+AQTgS311oJmoB8NnQAxxbw3lMXHu3qLXlLQY6MJNv4MAQm4c3mfdH2a4Y
rY05MVgyXDZPBdi5sXqCpAYdAS2r/nUUnidOa6BrsSI6d/fGr46gliqILm/6Xkufv9HPw+sgIhav
MTcXggfCHhp8Ek6VaIV4xbheAVE1HVuoieQII4LdY5sY4MzvIkipHPq4IaSi6vKMuq0MusEti6fh
loXUhwjjFhvUN1hCI3JzpBYAlnxfLf48FS0FUAbY6RXieKpKa3mK1yxIZOEL9Q4oX8RaZ6h3/HNJ
DByqUZhoon5x1H6JLK3QRd6adagJZcpP+7ZI8KL1ePTv3u7/rQcqkEZsZQdcPBzV0NCIGoVoorFB
W0WrgzRSnpHj22/g9k3BEa+F+JF6CERF4UEK4OKT0fA6jIprgRoYsj/c2E/5Cy5pCp9/CoBdomXk
E2CNsFwyHx7JYKiztDH2ISW+XHqmFXaeiIcH4SmP8SsuOP4jkwP4o93DGuKC4lT8CMmkCE2Mlk6Q
QQAhfGjjaAGiUz4+lvQ+s4cryeuIrNG9uz2XGbhuK5p/1kqwJNmQVlmYailX82ZEgkd/Nxlm4MHr
oYwiQ7C6c7CMPpAlCYc0qH28O5cXfuLzqSMXx8Ge++wiBBFx9j6A0RKMV6mfllTT7WxbzqbQOlVe
pDILwZ6gBMRnYy8RGKkLQ9NLYHgT2PGSxl8Hf+jwxLTCVEWY7iXvBWITJINv5U428BEYCqaD5GfQ
+LOVysi5Z4FJBfsyh1qtduJiF/ZntXIIIWe/732Mf1p7qEi/5TxyuWp3Ehnu+9QTp75t5L2nwbM9
EQIkzSBOPGLDlbdIi4STmXL2Y1J9e3+U8r4TZBiqHcaxP5KeEQhFpdilIO6aQeyeguXfustu0BLB
Op+x6NBppA+qn3PLFd9ywW+ZQ0iqxzvVXFIQebYfSjOSgSfY3uy+iqfodoygF/PvSrck+bolFy/B
hoTTis3y3uQkNkXIt3UG9L3t+uflDf6L5QVp7oeiCwUA9+de8rc8gtoCaItVJEzsEGNbJc2nIdqx
3lnMJrb89jGKUcCs6sgnKYLg4sZ2Vq+ICOwIlUfCzw85EDImUFwKLrKTdg3586qaCjzIyGvUYa10
05v6pTkQde0bROBhbm+fNYFAZk7d3Q405SWgUHS73b7j0GGRbk8isaFQO8tTPnyn4UXNZxrLYR9W
rsysLc30Bp06Cn9q/SHf1G4NQ/eT/4+jLQJ1T/b8hAw1jZqkuHV5204jDJKdYuPLGkEqfiri/cdp
TdduTKCj1raEwzVSGhVEcKVsWm1ynM/VNv72Qk/wGcSRz5JHuQ1M2L047KwIc0jta9jrAX8a/SYb
WpB40TPbFW81MncBgPW/7OfPclb0WN4jrIy0oddLwwB1teVo1maUS8mUQg4JyXQS07JxSPfuqcIA
D7A54WtzhiZwWg+yusH/Ws6CyTHmfaZnUSyCMcckyCDEj43ph1AuOXnQ7wGlO0PDNJJ1+HoJACQ8
llxJaESBAWe4De2ilt3BkfWnK0dilWxavxY6eHXQXXR6DcFe/i/SZosQjNEp5jd/pJ3wS6LXhQX7
CM0/Fgu6b2LsCrCcbeaDF0pDgqqpsTUIOVlPASo11G2hje4OlSklPk/s7c6Hse95WPggZ88DY2YG
/kdhqn7DMgrR+e94hK517VVVa3mKH/C72gPx2+IA10pUc7hb+NaBEltN/BtpTPOs3mUVlfhRBhT1
Bg8MNIarg1NTJz+4yhalJ61DGkRc9lXelsO4GVE1uU6MBfN1cmXN9xI+LxwoHJSzZqW7oEkx8SFX
n0mE1eKGVAM47Na7fhjo5lpqCrA2NzRU4E5+SX2iy5EuXXXh1MSLCjsB4QVlYBGZ76Kd2u+PpzHV
xFk0swVLYg00puKTr8j1z2DM2Eb4hPtlmFoWLvnLYn33Pj3I3b2U7cR3AjRmkOWxcS0XUUzpbTms
hEXzkZPN6qjk7pvG+7bnRR9HblbYc429WlK4w+rEi/XuteBohp41+0aGVPquwV8EThLKa9kzd9Rb
zCgZ/Bjy07UVgHrhdy0H91zJ4OqFC8fGL78fIsmMLjc/IX/MFmZ2B3Funee9ja8Mrf6kdY5+tO7q
/t22X2zbovcYjvQbdtMXtvZQZvnBkLzVhPCcHKPXv5/vnRpKgS8cycXXyiWIxve3E8ZHddd/t6Aq
Nc5B8sA3hd22fhc0wb63HFsSRag5DgOwNV7/Uvtp9NNYgSIpi8LkPguAYborlDEYtaZ4C1dRMhbf
v6oujHLJZ6/TZOvX6ewaoQrUMr+mas1TJ+ic1pSrn9m0zM4An+fNMVFr2P03iQkvOZYKvGZOlktX
3gwt66YQoiZrlxavyR1Y5k7RalF+x45iyYxrgd5e+TFpwYcGwwM5AvyhkAzHaP7m97Zd7c47AxzB
dfaDsL6sHqEu3RgIMyUtODLrz9SFcijP6kjHpi5HdYXmKtU2167ZpKY67c+yi9E4aoADYTEh3ZSE
0NtSkh65roDQUrLi+DsK8Ps7lHF5oXrWfl6LUDW7yngqUlEpAAP9ZFTHDDeEpVQJYKb6qeOC08Ie
8BO2vQSJman1uoXZj2bQrTBrPlD6ftFAJPbgUmx0Y/tvWM6z2G8po+vovGQZoRvgMlZiibyAt9BL
x1OnrfdIPN8tXoGCtG6+4hvHQBnLogRL+vXejwf3TNm5CUAj1JV7Qk8my9A2CH1CfOqQ9m+V1q3Q
FMo6YdEkib8k2jWzAOmz6al7hhQcxbvqkIYg6jrA0CxuOc+PQK5H/AXDLAjEzShgUbjI16hwTA4E
cMcuSMv4sOVZNeFQr6S/XI1oorBQmFePREU4GY6rECf/QTSD0AD1oVWGufx0dq8RHEtcYVVDhz6Y
aCMJR2O6hXhoosYeasuLw2Hy/yV9l0BWk0imysSPvgc4ivfGimvQQIAPbwpHLV9Xq60BJEqmOFTl
sMAiZrnieIjXwbs+zSpt2nwcg+dOgubbLC68FZrQoOXLyM5oQ+0CMEzX1rnAFdirgGKPLlB0cNQH
4rDHYUjrHvDR1lOdzU6EijBoBAfcJw+wHWrNUjt7j8sZDtzQRiudVGOf85golghG3+Hm+gqpL3uX
GyEv8xvyiGlZq3jEdZKl/YD606/jFSZk1HAYS2e7gGp3+kPOYhEXw3Zcg9Wzomn40U7SXX8vebDs
H61nCIrHQeRpbGCvgu1wt1cSpXdopKumLS9v2a81cKMdVwJ7NpnbjQuOOUoF29n2d2XATMGVne/1
1zg2hwHuHxrnLqvQfolTgvj1LEdTPHny0rdsjaAOLQSoSZYXX8dwz6Cq2WqCLStm2CsQ1icWvWTR
yBVCKjhPifA2u1/pNmi/gDyPgoApbKCdoxVJuPPshusveMsfwBRDllNoeO/KUIZh+rHPCC+JS0p0
RqCFmIwh9Eq8fEys4w4NLbeqWp1mXxEh74l6PmKauebobJqv11AQyUDVSPi2h27wZVyPQeez771/
JyLwzzY5gw27MXamaHHcQldGBgPbs1kxA5xOvjZOMpyYicCA9y1qOalpdRRXQrdBhM7xnbhOtHfc
bn4xLXxZ7zrrX37dBy88++zeKiWetVjNlY81TmUSMAmEtdBJ8n/ca3Yc6V/5P1esLdSxvL37XIUz
lfcT0Z0TxHSL4Bh13Y3H8ML8G7ONI/2vlH6k9PAIMNmu9ilJtjrkL8yRGfQDzeH7GjVxV1RO+znj
wJX/2ipRCxFVfHehCNZKMkZjoxDMSQg/YPTdt2+QQeH5mavvthNlJ6niqnYHKJFf69q2Bh1pTK0G
qWE7V018xmao+2QeEgXtGgpuU4+mGK3lStoyJS0qvO9hnNbgzjciDrxQlbbM5rFtq/dnPJV+AOzU
ACsNyYYoaWPXhef1PSl8PEqC6N9w9Eqd2b7zlkPB9p198hsvx654r37KrikkvDK5BmBCUzU8aM9o
chjgJBAmsX6dmbnVbfJbMlLAXllEO8auOsMS8SkSg7T289ag9YnTgeVPOdjS+yYfAMQ6L6p5s90l
YJ3hJpj/7SWmtXafQihUhondz8Rf48LzvfMLEoaqEk00WXNGiDjiC06sdfiTNmbyxl3gtsyJ+S/p
I0vI9tH8/S3dIG0Qs8HhuYIPTjuA5UA6zWNiFKBg5ZpOPvNyoAGJ13SWDhoHcWmbNG/dpMHShT4D
045uXjR3puXhL5gCyhT7DjAnVC4wUALv7fPVq2BLNIQLHpnMiA1JbmRWVI+sNWER3tn/tXm9bqOf
OlJwb3P1LdruTcwU45iWrRmxjBsgbtq2lOZWne6KqWRmLdjoiy5MCv6Bg7ECTYO9GteszhJOSYWP
sc63sTP6HGrEX7PJQWqVXoPwDgIsP+Esw8G4PLBWB6ZyxarPpx2UGXweMkdniwmO2e4ELhfuUL8z
SNh4t6kf/O8VrLc4fuo6z6n4ZqSNf7EPIoorKqYdaxQyz1VRlRQsyLjMsn8kiiK32lVUsAgL/bHM
1AVWXQ8VPwi3YbvRu4ZZ7KBAIxuU/2bxMqDfeR0iAZIK3Xptmw1rFPFM9wiGhZudrjTM0NxIkHG7
eLxNOrjScoX+0JDCuzf3NKMfHzs/Ygdv62wgHpbANuzqoAOTZcBP5i9xq4zMq5/7JNfxZm9W4VRV
duYOX920ZaxC9rveCyBHhFsNoxY9ic+6sBjxxOX5Xq5IicIQk/uHykw/2fUjBc53ujeMGorEJhYC
koBNCJk9D2XtRLGOhEVtCqFeWZ3VnL/iJvHQZEH/pI8/dcb0pEgfS43t+qBrbnDvSsC2hmNxkaA7
MiEh0CtpmGY5XoNUU/dn6FyHGjhGhRiqFJRBFl5sVE0Xof0B8Pqlu2zT8TgUr4n/cDjGbKC0YJXT
dv0MUS1bscFj+uM/ZJmYsNJTm+QIaJVvFR3f38uZZnxzvpaenpppgx6szUS5TKZFOEL8mCYQRUGm
GiS/CqVSUA6T+NGyatho6Yw//NBeACr2sOjdbrXE/06cKljtTTNoK1y2xUXDd/WYE2CtLbZrKO9z
YAT02i2zxYnCp7LR7nFKOcWMFBi5fTLX9lxGZF6ieUZezgH6KIwC2qhRjcC2fyrhgkAlSSzY6Nks
k29eShF9C7EKiXCLLcXoBTF/VfxX0rRcyVluHGRTb7hRV5GX7wJBbTdzyowjWqYfwdSXYnySmqja
FkJ+D3bs23ueZE81eRLNzza0WsXfV+tEeHXjH+/TeUzgQRFoBmdJ1Pdryn5g5wRf8hDT1aRQIM+T
X+XsuWoIfYgZCvyfBldQVSANIFCDc2GDzP6Amz4yMgTuKEA8V7MIkoWxwmnVIpO3xj6ieHERBrk5
TpXCXvJK28VCR/mdQJ8KKUryf9/CwQGrjYBPfn78g3duuzzK99hME3zvQ7LHFG+0w0sOPxI5mZBg
HtBQy/h9mMD9J3y1ReDtrQ8lImxYZ91xW+D10H87G15RRQgRB52UEKEdN+lrhxQro5FVGOb+Hyk4
07JlWmsDkkA+HAmcHhn4c/mEagXksEo/uRacFIuYegS33RdUUbt0mnpDGaE7qffdTH4IzS4muixO
UcxjfrfP47r7SDqvYkuCqJqKhsuWYvQIIqb9F9Sp2jRtPlKzfHN/ze3vRIZCszWlDSVw3J2M++XW
G7G8hHLLQFh/rhpjNPltL9DMeUcxVr8buDuolAkqYsbjZV//FYne5jyZQolDKNa22jvMGRcRjKuR
Xmkhr7GCbjDjxRGg+XIucmAKN5WqZnYGJmmCaeFOFilonJNJlP/anWeqlDIdPmLThTo67vbQs0Xu
1tdjgWu5/mgBWTJOsa0BMFuHMsbE4YKBT88eSYrmtoy6DRryoYvWFXSqVxdtDLQ/XTwV9XG1y6lX
fuisvqD2V/kD9HE9BYUfATWmN6Y1qKi6BouvVB/mIElh8ahihRXXKQ1JKF74uYQZFSJUu4m/5u6W
KN2jJXtJJpfwPo8NMqCbcuT3+CVVlA+gVxJb+Vl2SdmJ1P7kq3PFJ8OrGg5ITWl6N+VBvSnsII2L
fDkFr0sSma/vbNE+i3e72LrAa/E8XfP7yVvWppMqtUptFWM+GUtwJdHWpH43nZYdflQBkmVqePzJ
55OcOx37WIJYOsWtWytDHxRqRr9YSo1MazM3exdExP0NauB/Y8VBcghlRejk3lSLrr9spwMpNGBI
bUEJ56MIySkOHIu8FZG5aYnq53VMOshhj7MCw/yIkBTwRPTabBUtuOQ5Zu7EVSzKmSeOlczUGRWu
p/30ecm+hnUM0lglekJn0bP7oJV12drqVnfTQp6/oIMOSyDohTwmHoCW8gy+xNsAlVHFVEe1kpAY
6xapJHaowv/usNKitXVNBZkrZl2/ajdJ+njhMnj1vGFE/TE+UkBMaWJ1VUvjAwbCzpZPEE5crPQM
rmSJcyzXpTxxfaDS4qhyqkkNXgCtGmq0oWZR/ihjwHRHbzo95XAkp4bRmDAtupeXUwu/lx7oM4PL
4Z79hiFdPsJ+a1i/UF+XCpjeSFTUIgWyBCS0U/zRTqPZVIYlenym2PbhdhCTDE2kQdPeedSwK5h1
oC20dMecAdb6pALyJptDKin6ltazdvB/daWUyNfsYTR9I7xSJf1CFOSMecScBRAXDWdz8GwRXcXw
S4opmQJlbaqRQkNYY1YBZ+zUZsN1duWFt9izP9vU+UYOICrKlclS4WPmBwiyQxcdu7WPkhqpP0qg
cjSxkAWypmbj2E44QMZOUOQWedIe9W0wn/RbYfeEHYHSDSQQrWclva5ytBN9uRyiTOBPa8ZuBNFP
moswAKkxQKTuP488CnOBsOdQxQ8CxYeiGWjhtvl8OS+ZkIvu9Ai6pspp+5pmT6igLRA8bLzqs8r+
wSlPI2DdHNZooylsGj2srUA3cN/FmlD/u30XGW/i9B3FLIm4gZLnqgIf2M1uGUG22WkTTkqU510X
oxC1YJyWnbY5kcmnkJaww/BLXTWzjkj2QHdgfjxPDU8aG1NcYBzB9LjdfyWVnAG6gC+Uf3lrlfcR
nGg0TNsh4zICrnxGW4iHQ48xccICWD0q55e1A12cpwf2EJuigFJz9AoH3fAAOV1ZLPvXagtgB18O
FKdB4RSFxe+WpUm8dc0c5l5gKc18rRqCkutKkACQBGwoVEBewiblKoMnnqDZSAnsf9L3lpq4aXsU
ozp0ciwjlPboMCr0520YaAr+M1WYluxKVd353lNJioGeBQPucGUBo4FGWmML3Fmox9++Um1ZZP6C
49SnwiSuWH3/g34u+KVX5EGh/p2UargpuEIgRxxp9rGV9bLs+756ffB8UIuvvlQE+ijytUc5vVe6
7pI8swrsoFdaQKInKAHA+KVGZ4VUNsFy2ZDDvVKYaktfEa893nb35eo+OGah7NpdSvbMqP4CdkI3
QubFxGG1udgD7ggonhIj7uKiypknEPuJHTU8qB3Hm2V71iqK6eSRUXRLf6ZVPgaSrpcT4ZAt9JdF
4CUxd/bcv+EnbxSNuRqbO59eGRT0BuZRNKAJUW1STT3eGsNPagD1NF7P6y4l/wwepC8JCbJQ7/zj
dfbd0b1EA6/umkLxY1HU5KYZWD0v8VT+7iiOUoPjT0yx/ocN4NEidSQHsLcCu2p6YoDJ7x+iZzyZ
F9nLgZMv/cVNxcLOlRFrIMX8X/nQelwWoQk+56E3iT3hLbWN+Lsa49zXy9QhdkHLczvO1VvLyYr4
cXgCH8/1J8D2iQBK3VqB8mwrPkRQd0Xf/oFarocUlF9Q1kx62DdUL918r8XxTFPrhoNlSjgjLOSx
izyyIb6TfRGLV7eWcwX0PuOySAKBiGQTYkcY2ytbeMDmb50x43idySytEDk79bkCTbHEPHK16IQz
rJ9UKjs2UAJWkDzwFkLsB0ZTA5729m4UREDYcgPJdik7/x5ADhpUN9htNtK5SvHxJfrHJDIIyLEW
+A5JIAIJIlBanEHalhhaS+s1T8WAjahGpVZtowo9liK+tcBV3Q0Zx5bqyKvktgs/cVWG8yzdaQWO
5F9ejer0KdL7pS/iO4a7YgPBxiXhNbhIgTylLkKLBqU2xkNp8ByPHsQYL0BuJCwXkLOrdrcmi/ZS
oX1m0/U2sRTiCtbCGQAUZeykxSQoD6BcP10G7yjAB9elN55qjo4vRfLZ/tI0PxVwX323LwUe3PDS
Ky4bBN7KsRp6AhhgO81vel5o46FfXA1ea4MbrQhMASUU4duS5+y5e1AAJHcqeoKcvY/iI8Kkqp7q
53/4aGleZmP5VaupgRo/KifcnNuNz+/c7NOTtP8XBD+rdmgn2MIaXQhzIyIHXpbeb4Ptzu6O1Cp7
nFBxSYzctSTGRJtf4SbicnKm+YWwEFZGFcQK5xQ2uOauwAKwN78Z1uY23NtwMNjQV84yxy57FezW
DVDn7TNGki6xTWEJbTL1nJb3uLTg8RVbkQSngN+v7JsDIeYB0p+NqEmKLqw2ytF8MR5OI0M1eImA
Nx17UMLd6w72GIfRWj9rv96TspdIg8cBixUym6uKhgzaWAKBHMaTA0RgmEx/kecX8qOWudGIoKz9
SgrdCNB6BEc2VI0M52xKZ6zeUCOTAAirSsaXMkq19yPfhLpd0WTvQ/iWMZcHfo5QyVUWoK3wpSA+
FUwPxJQsUWId8LxPxT3xXEJWBPN7Hz80vP5GRDINoxMRhJfOOV0CUOjAdst5xp9fDjtemFNgbhx2
paWKjROH3nA2k7dgAyrIE9e9iFkI9wwGJyQ5fEs10XAOMa82jf0vv0csCP5dnwZkVdW6xnK3jjD6
EoRGMAjROApFag2f/ph+5RN6LUk7UDZSG/3bMsmr0N9LlRpQkgvkamWKVYOTwznkKv2eCnz4/+iI
i/mdrGHw1b4c0HT1AhjBk2RaPDEQaCVL7ZKaoJgTXRuFgjlCckWxdHZhruIwPIRjv4/e4QNkyt+Y
wJcDz8Xq/lcSTUESrGFWhOsx5nUW1IvN6/zp/d34w3b1dQclWd6mSaYn38mX9LMhiPM6SVeY8CbQ
+TC58lDFYZnf8kedpcPNh80l1+/ABPEOvD899BZjbVm/lz+a3R59sfFxgPFrYyeJtIkjyzdx2oBD
vaqmzhc6ziamo2MdSjDmYj5jufLPFGRYQwWjYKnTXhBer0S2HMcBMiAHiA74BzTvvSpvjtGLSHxA
IxEjfeSO7PybCTBG1m1AgrvULHnfjGkIIbtpsjLIlEYHPdKrJpHxWdqTRhbyq4Z0ER2UW7k0D4t1
YFdmTaC2q/w1nNyuyiILYQoEFCTGAdqa/Lr3ZGPGyM7FU//9pejoJR4bMBwmH38hjfC2Jh81iEgS
R+GI6HX6J5P1aHLOqnFZ7RU5j7cKIPlNxIzg/4b1GUdvK30cglJWODobieLloWTI3a3VwBnxlGnx
GY91CqFFnjn0d82woQGmvXqtfto7jHHCLK47GgryYcGnbyjmClcIAZda/pNlkkKZnlJtCzYmFjhx
WGeockaSKBGtW0a7ro+od9cZtz+KclDNHEi1TdvDRRwBZNkB2n3bj5v8tSoo2m5gOoyU88te4dEv
fXoRG8qR+Q/cFLUJgEwtUPlogeggIv7YcHW/gBygHNfT3p7QCyyS9cga//qrTNCGxPNMnCzn4CJq
+4V2RmrA6QNoa78Ge8Yn/0xFrzqX9CMbL898FoCdaQEnF6rr6D5IAiR02yFPbUWtbijYgWcfpXC1
p4l3BLsetz6zq1xUllnLG+hC8EfJwxAoBHLa5hdzxzsimhBen0RLlrByYfTQZcFyo0d6dfpnwqiE
DFaB0/NdtBk00zNlMFxZOQ/TKtaBU+9Qxke2650SBOua/RxNbG8BQoUFgiwaAkKGLH0FTslL83kO
wDO5L4RWXdsla0zi8ZMR41Gj7EIa6PV8qUamxjhLvB+ESvTx1yJ0rUNaRmW5nq2Q41pk6pACTs0r
uhgNTSJ586QhIjhwQlxgNAiT+DwhQx4kHih53r+F4lgreemRgVxGYDunaCv0rlVyh03ELtHK2K56
Jc+XFgszddx4wVOiWr1A+SZr5+jY+qI57mTMIu02Y4y4X3T0CvdsOjBXbX6Gr8H/1IKyFDpN5NLe
AVcBit2fGZPov9rn3kWsdwdiBovHloWtprxAyVgj2Vv74Ip403eKK0fsBgG4TIb+l1tKb/w8T/GK
hr6J+0X5V5UcDOFN1EA9TYLXeFNCZrN/NXr1I5noyul8/S+WIrCTjcA1FISWyBlj3A4rXHbXrdiK
gMIEw5mM6uNjE+ED52X2mH19ynV/E1mDSIG5M4b4c24JTN0wu4+or4l4mHPmvn2P94haIa+WIwND
EXsLasX2tM4sAxM1yc0Lkipro1ohTReavu+HdpRVRCj2m0Vzt6kfAswSI3AF8D2fS9xAuDXQ80YE
0whynpz7hdEP5pg6WlKbfUNpcsxVhR0kLeTgh43KIW7WIQEy891PhHiHApB8xZzz8TVtVHQGKpZG
Ho9/N4cNjPa/NhOLLqo3VqzgfBsGQq5jX2SmxR6T0jI5SxIIR/CQOOqJKX31jKvqz7y7CV7Yzpuo
wzjQm2TUqkDIi0Zqu/Q/lxpcCVlS90c0v2+Df3BPN9bVBJlQr1sHTTiAmyNeVxHn1Q5Ky48fNWxU
29Z3Zy5GoAAXVobs6A4t8IosffJx3bp8tFPGGF0ZnHz589584ABLd8uUw5/jiY7nJkGZo7ib7p24
8Fsu/F4kLW7zibJbnYaLjlxQ8pE/gzFnbYHf9uou2apG20rv85EiZySmt2ccH1I0WCHg7sUKhGxo
UtLuW8gs6CgdVVEcCKrxDpItRt+2iQe6ILRPdYk27Kx89l796D1DEanZkt+68+Psj08O3t/OLPtp
4EGOHJMhU6a35BohwErstniDttS4QoJKRJ7LEGeXzRcsQk6v+WnGCCVcV+Ul+C+m309QpiZkGq95
y0dgZyP6oXFmi7c5UkbXrXoA5O6tmoSTUFYGa8ERjVtg8VpJtRHvq70ZTyAz6n4Lknwcz8/0ZMsJ
krjRkHmRId1SE1yBu/LHVBi8oeGwlqPw4LdNXsu/4POAaemBfYnfyrkqobULIV+xVGne4IrHwsgf
1xcH3Hl5HJRdScvZ3HqPwzrmF25H6Vx09aDcLbLUaQumuVNsTvQ8NyjUPjzuZXqGpW+8M/KmJxnE
bVjIfEW5S8ILnfSqEEMNKI1dhYTkVQEI3/NxW+TxoZ9Q5gl335o/hjU2hdk56XUkG+Dq1hOgEbFM
K+CExpk5Ua3LP7joqLY7jQ42/LbqmaVlCHQ5fXztJU6n3pNL4tPyF/0oxLG/WPxigLUOOCKWpS/i
kFfz56ZAkYZyIvdz2pn3iWPGf/2SVjI+7+Hu1DRz9NAdVTShYpuORFv+SV60Qe/xfj62yAsw7riG
c6oX4WOpSCBjMN+VEFTNC4e/0WgiS9QTZWg2nkK2u9dQWuZLl3rawSLtRaz1oe/3v0W61JY4tbTy
Et4zv2vT4ZSbbI4Y/k5+TLSw44xNR77KBkNky45hiZ96cbUpnYFo71YObuTjo3xvnzETgZZD114i
N4+eGNw07ssbseu5PMeK14rrG7bjkDWMfv9TiUeAqgd+3zRYNsSSsgWPKXu2tn+miDYlxBINBmPX
fURqNkG0qVDGNoJU/zdYRBaZm5szygOQ/Fezc6VKDCVy4k1LnqF/vYAyLM6OE6+03ptZYYJu8kxR
IfglAVshbGvkJPMG8sc6CuqLgT6ziXIpX0pVCczl0AUgH9/C8aq0kh9Q1KdmUM2YyQkWHd8CISPF
ug2iJHZ2ZOOTCBlcU0/FtwRGIaagjTKhagiH31rcvgmLw/CoaGhQ28y8HaLsIP2ngMsS/gu6WM2K
Q9nps4do6RtHyeV0wnwtSR/RGp8DFc+8svpnk1Vdy7yRdnON59jxuMTnTyNLTx+7184gpw5pBJ4j
jg7NzgU3WC/LsyDdT9nC9oIXPOK0hOkUxkwR3Xhak3R21HA3dYk0z6xs5IctAE2V4k0OAVCFYSQo
4bHQKmOOzS08imlgBtD52LPjJh1LA/fIeP3Tll52d/NXJVAh+h/emCaSCVO1oE4iQmsea5qlhZnp
sOqA1h2LzMTN9KAZL6sv/BrlJH5G23B96a6Ij774bEmp1f1ru0UkOLlPUi7HJ+Ot6QE2WgW2KKga
Rh+LTco0Kf3Eu3Vg6pjOjjr2gj7mYfEpZd2wHL6MNvK6JqK0pjtLLmuFXCrprHxP7I95clrRhi2A
xV4EQ8SdiWvF28+vhdbmjd+TVU1GB9zHx5UkGDoP1Ft/Lhf56O8Y8vOjLzTtNgo1w0dqeJuYm5bl
jhkxNW3qNWkadxcIHVlCq+0kYVdjGcyVUuKVg4cI7a875IjU3P5UNG3KxT2wF9wNu3J0oXXPfnE7
J+lp1ODqWVFldyZcCQtw/2vNjvKycPgJAdaXDFTv/f3Pv2bMfYQ1KPChqxG9D1Ufm9gBGrYH2zZp
rZbfevZkC42Ul1iQiC5SfwjTlCxDyPdl9Wh2hKYBGWaEKk1No+v/U0wRTq7W6B9uztq2TQdi3OHJ
kSergXb4+0ftdl2fqhvBzyljIp985UshPWtVpwfYM7eXfxa4VomiXHf9nGGhm0FNnRT/SbkZ8Ipv
fR6SxV9NWZZjN9MpvZPT7DFSSHlXYy7YYy8kqFGRZK8pLcgMcKXuCoFbnHf9xGjfnp06KfRMQCMu
GA5feuSnSwHFV+uLf8CWz0RksOmWeUrEpIzPRywmAAVFbMRMIiFSjpBw9fcv3WKubOBwI4SbEhju
xcKFwWOSNxrXCkcOKN52Kuo+99/wDCZA0K5hcC6MMc9Oee76N/TphLONcXjGlqHhlTetG/l9k7FX
U2FS5Fx1XHKiXctoBIi4T+6uIJNksmXZh9ZCfTNsSh+Sq+ES8TAc2RNCufb/5PU+9p+pNoklve91
RoCoCbTPFAb/1KcQ53z98a7bJomZIRWwQRCIxbTTtKSnzfMe7CXHtMLLv7mm+cvBxsLPLBmGvDqw
JPeMxlA5vt8z+ibtcl+N+DGWCEgQK+5UgSVdF4YVbq05NulGiRFo4OtLeXwbTaf3ur9YJza33PLM
mpm23UL3S7tKOt8I83Fa/EUbyoYpHYm4gLCLhNospQHojVrKzBTOlLWTQUkf7jBBzSpKy0yUoMd0
ZRxitF0J15oSWm2Fo4d9ohhPBtlrxPsGWV6rYQPXwVLcS69aObqmGUUwgU2Joftv/CQx4Y8jFK/3
pxTZT0oTq+yiAWi1GZfu6NjbKK7v3eH+EyMBARRfTN2SRmqlmR7xwW9DImk4ZUSV6vFrYQ0OYLIj
OTp7/mrh5+k5tM1+OmrcbdDO8VN7cc+nLzJuPI4Di4UB6dTpzDSsMS/Z9fCl84obgq+kMvHoleH1
T/5/K2g4UlAIUfLWSu4APiwrD+BsE5fYhijBlqJFEg6JHEFOplH0ZoKeJy2M6x3WO2pjopzr9eYM
BvV/nkEYaQQlwulYhteXEGAC+0z0IsjAmFbaHSIGQ5wTTFza8j8j3ALhQX4dEPysbxpuhcuu8zWq
mbqGeoJ3bcQq63DRG6lCs+ZXLKUEtRGWZqU1gHqoEVRUfPpUP30ADMirc8wHNNHXoojCZMN+Pse1
1l2rQksX0wn43weV3mr+lSQNnMmhAcNdfYKiNsQZ0tjNn5gPGQLQVmnz92bEKjo8uH/+Wr1/uhrA
kX5l7fMhqvRbU3QR05ZObWD+u1jIdcNwxkK0deqS/S9RFb0XosVt51Ci8mBRchIY0jl4OS55/VoM
FH+vzcYdasPwOSCqZYV9KXXJGR2OTap/d5vVpXbDiqdhhOWQA2v1IyCEvQ53eatt0HHUKOw0GSkE
/MwzOU77VMJGaGyxxKdIkUCJ+bKUleX/GsV0DXfhjIKHn6JsyiDRitqTwfNO+Z3ijMK4+jVLGaHp
nzOFd5jIFNdP5tnnwfFiegTxX3Up+4yrLPjpIJ3MfXpZr2OtMixeqrnGFf/uS6f9gea8U4TDGdI2
Rfyzwya361oNZw4+lPODCrDTqYRtGth8mBTt3jJe0E89nlPl0eTh9Gj0zOhzsV0efq3NoPHmf+RL
dblTvnrcudu44IQl8l6CMx1MVeJp2a2Bd9p3ww5QxrIAhfm/uqT4YmtZnizyaNdQIz8Xj7bMcUno
jNu/ej4spS5pH5nteMm9jIh33AiafEK3f1XAEPCzn7Biu717lzDdasYv+FngOKGvcNKj/l3FVD0x
ZaaCPGCqhCVtJAGEV9dFMOTLNLADW8dp+O7fkjFzoaFlGKHUik4RDd+BYmG+9pczAW2gUwVHA38V
UPq0enTRRwDEyG3kh2gl/ZJcuWVzyKNRNnMHfZtLv5RCjtRk48jBcotH0V5faxrpJWqqS3ZLGk+5
88GBHt4jTR8xdAlmVo/VlJtX1NPph5fzidIA8D9GesagUKehXq25qIASemBfGb0oN9A1VzHVoSKM
UFsyC9mOxv/aO4h+PP/pSXY4I+cVMHWyMfQ9tl2HnNas2IBK+rfMJx+ztY9mR8R/bIT6B8Md5oSi
uQsn8FhL6u+2xZI4PUi57ROZKfCBdUP1jL3AgyxsVoy9oj7ivQ6fXxjfoHY+q3yAtKHcRXc9JVm1
rvVd8SYTIlGN5klJVYL4ORS4GlNQOzTM33Gjl0Zf8xN0HY7+6Y72fOSo1o4gHIwfActSVubY1u3L
06XuQjZnMt32URksbV+daq7bUH++yAECNbW1OFHoQUzuAPEF4DeXsfdtzlsKXYWhptfxgNjA8AxQ
hoD13dYYHCkWu9UZI9q+wyE4rKK9CN9ainbVFW9aO2NPXt1qr9+2Fcik3JTV8uVxbN0L7NZNGJoj
Tk5LxX3ZNiZ3MI0i/+L9FQsiFxrk6kvQ5OfCLxvR+seP+RJ3/hydNbsPZHmuL7y13Xy6ksaGoaL5
jUwN7+rMMmaWcKwxGYuYna8qhoAG+vD4bp4K4nLt7yO5l+F1+8H9jdD82HIYT1UBijjzhWtbP0tm
HQ/0jEtjojuANOqZdQXviFWLLrkjk0iwIKSgaoS31gD18rUgrzcvlSlqt1VrQyjRNVb3BREbrpU0
VluHMTaSx/PigfO5hs3bpT6oMOcHki4Wt+bhOfvCuVFzaRTR+lvXetGSSEBjxRwQ6YzVCcmL47gQ
BWVFJyISQurAht0n2HxAvV3Eg6kkjefTc23DBn5e6EdaBXIpLU8S6dpMKQBnpU18LpSZFQJOyK4P
9EMOq1D2DN8GJl01W6XW8YgBaDaqy2qFA8LroL2+zdBbHV2dnNsM26KS4VrxZw760CzaeHoRF5HK
2jBf9C8r/A8UkFHMyGAiEZeC5luCj061Ukq1QCIM9wR0wEhLyEUpVWDiUoEnpP8nC5f4WW4RKAR3
N1pF/2akf0lr3e5PhFY3PaCqIidVMcTt/td3xweU6/D4zyimaTHgPVKBtjLXIWuV/VMMS7ygg6Yi
Un+X1IYEaYp8jj/idSOdteg0Pq4bCzl1lHuOGzFHT5xGz5WginNJwbpi4qL/SNuMXz7PajxkHArL
ZsTivPh+A+/1TlvtjqNW84KUfAmJIS3xrjSQGQSRI7Ag00vghLhBnqM4xr0Y5uRvFb7YLrhrR4Nc
gINnDIyfH4tmIuJX5GSPQHRwPmo7kBQW1vaJitPo6yqbWq5TU0ENerJEg2x65wFzqd7xwc8WNCJS
eXZ7AA9+ZCX+lk6sSLkWPlbpq7kvcnj1sC2F1ydAxpxA16iz6OdBeVo7WtUOb/6tR+m+Nv/8Ks7b
g/LraK88UT+fMKA/G9ka+NUxTx01dDZBTY80w0lYcyPc9La/VpFmMY6XR5srg/tpk3S+kxZLKWmV
+BzN0Mvv41DX9vGmRKoXDbaZC+FYxqOt7KM5+oTtL3iGd+/SSGCsJlOxKlCwE6SQyL4PRwXpAys/
Aob4yqcgFmEMw58TDpi5Kr8t6ClxjSFFR6vWYDQ1PJH2h3ooCh/Y3tjViNC4ZKgyjyXu31n4H+et
sX9QIe3hu5k9be9qZER2lYIbU1LxaifFXOKlJ83d/kr6a8cNLpMbUlqm+P2lVIXX8pWRG5cEz7iT
U+vqAfbqhOrFvlZiX0QEHiHkaXhD5ZRFLdAYEVBcs5WBc9JPpqKIfvv6KSeFMBNXrAQX1uv+TLfE
sSG++FrMC7tHrEmpwEO3SuA8S8uvrG/BQHnpRNk2hm5MnVmH9mgId6VEUTdAEAuM5Sfu5pK6DApH
b2zRFFEXRrmNHJIVGr8VVdgWndyEWKz1fpWwvnOxPDPvQe8mGZGX//u/b0ZGTQaqeALOX/7ksbaz
pOiNt2SFfOqBqWmQTPDAM7+HW5Bd0EjEQqar/BxMI8lQgSwIxRz++dGxLSF8o2Zn3mlFeaURVMw1
Ic7M73JAPQU/jriWILzxN3fDLyx2KV283FEBkn8iHPX3CFpXTEMH/E2STEfZF2kWUNeOZKUYlyMM
LGVoaMx/gwiFMT/724GWO5OAUwEA0imVmToFmt2apx/AvV0zDQ5Bg2BwpA6TWh5umi7SifM6IY9P
cviZ5+t+mp38ftU3Hl3KwyYOaauqM3Kw/AkbJ268HNFj/DLjJSll4zWDrBKfef7WiPqx0a0ZBRLn
qav+iEu+CTtHRQZ8DtgZV8Z3f6U3RTh6e9CF3VsTa9RANSLQ0W+t795w4SQeA+dULKMZt7NXKbEC
q18RuNaDHTOHXsF/r+3Z9/mTSMTbj9RaD4dbysPKXsduwIDHsq/8vSDsNvRNAH1C6pCfjrfP75gQ
ryJVvS5/5sOjAedlcojRiEejyGnFGzlcDSXah0zsgwvU7BGro39Pj8IGcaj8zBnPB65Oi2IHiYia
4D2NtiyFpVakGxKMiTg41dwoRaPF5gRMNRaM6amHve26cozyGlcpb064ETS/paqvICAXEdXlb8XV
12FNIlpjxh6LJXZRnn1Gbd1QKyGcOraMlORoQHoG2SIbmf+7mnRgt95l4CFicUTamNHQtx4qI6Tj
2iew8GIztkQfjvwHUDNRMS94Z0EG2jboJjwO0Y+TZVMn4XBguQZJJ2kjkCzBQswx5wHmOH45LFup
h/C44ughrSbr9UiSwLqCx2QcFhIyLVijiGLBvFidn2fyQ4g+XPYMPYNyDWY+WBDgnkm6Onf0BD2x
8D5s0p/WYFmgI/srl6iihvOGvaokk6XxHjy1jozTtH1P4JwrRzNfqz+8O4wqPnNT+jd8opB5rEbw
FR3xbrVs3Zl+FgvpCwkFLbFn3FwvbiU54YrGsKdvWx0eejrbe+ZTMfrY2u7sqso3S0L9Mred2kNk
mtLTHwQhwiySIGwyUb0DIXKZV7WoE7jQ2Q7rj1OuHzWRix39KDwQHcYrjn6+o6r4RSPjHf4Z23Cf
KBlS6uSP9edD9cRSQSr4IDgEqxp9i6w3oBoNkK7z7spfL0xE8QZCvXdQxYrkb9rpiDpPGzLwCAou
V65K6kJ4jSN+3tD2l2NEpNQYp53UZhcdxqPJKS8+tykOg3BxzGGsRHAc4q6WqBVt12e4kq3B9Yyr
oOvG23r4+N8kDJ5nNT07YdjnHRpa4utfVkiw0+jZGoxe56mHvrOeypbktKsDgFEcnkHnFdyvrJ3q
V3+3wFkx8DPPaLV5z8xgpeuWXI+XfaNNdqhxXnHvQS/mS4xE7R9iXa4Y/EnzNGDqsF5+lPPY3oWU
CdgIfTJrnvGlMm3cyh66r42uXSia9jqhQYD/hl2cu/scOu63d+Zb/kuQRpnfR80LZTf125DHxXlK
3qLZ8EHe810didEwFmc4CAWz54dUw1kBd4qzozi1CjaCD3wRCrW5DMu2zFyl7D/vK8QZ1gU6D6ul
iV4/BT7pkTMfnJ1uDULoTlc4ok7FsRywij2nFw6dIOtYnModDIwX3XV3XtZ6ykw6Yqzq2VSEA0gU
uPwqOM9zJXpkuSoE/1AF9kTGvlQdprxAobPK1OJeVAW9yYuy+1z67WRTIJIMRbJMH+6tuGZPCS53
dLimtnPqCaqN9JoudQypuYPF3kn23Ib1R0HSxD0zWVTOgRbLHND8x2qyv6Jp/9PJbkjFijrUubGF
J5U1xQ6CY/2UzXSm9db8gLtmsFRFTcjfU8R66XZjl58Rz6Yd0Lj16wKs0TZw6vB4hNq6BIdfTndi
KDpfVGCT1OUC376e3IiOhZDV/D2PvooK6g0CFVZ8zPI2ztqJLE/fAsJjGejkfgUt0QY8ZaPw//5L
obRkk9J8mVCbeugM82GoeShkwO48oMVnjPmPkudt7PSMF+qUhi55k+nRX0hvGO34d/JV0XLla3WQ
7JRFGOuBggcFs24RldQNYGK5COwqv4ZBWj/Jh8vLuWo1NGQAtWvWKk5DbuFNeS0Gd0Vm0d/UhZI0
q/nlAdI6gR2M6eZisIjBD/Oqg8RhweDEvd+u+l0/6PATrJ/KJmlB31zodQY+F6Is0oCXKuSrXv5j
UG9DZVX0+3xLEa7dYI0WAHOFApAQ/ZoomKtYXWhDzwFQmzLvF8SnHRUShZiyAh4IG9YoAN2/Iy2j
YAZiN8oY0tjDrJaxQ6Nk/H/YIPG0oZ3r4IUlwLU58MqkeFh7/cYQm494r2IayJqXniAdSff4jxsD
9b0j+rgIeI6v5uVwVR1shAQupSZ3ZRm2MXgM7ioYOwz3jzvGucvCaQXIRITn5VMdz2mYfgIjak0I
33SdNfq/7ZgipnNmtEPT4AhXu29XBCDLM7R6MYcsffN8XR99RM0URE7XaOlri1HnL0HBQzQAhcB+
bz/OXazod69jiDJZafCcqRtIAK5pMM4b4w67T7FLgmXlFY+U76yDPFJtj/IoT2m5pTCkC1MsvLBm
Vy2gKBv9FMCPjridX5AkcVlSMHMYMpD7CPTiHScoSRmkQfBGk/szrQ1ggioo2GY71UqXEhskfENQ
j6FAX4sRSo8Odu0YN3+4NphDJIGcTss+i93jKB5/L4dfYDAAZrEQ/Gxs0RaWezgmIUKRHX1Q97sl
2ihCzYsyuCy3JGJCuNDj2b16VmuHva87TyeBWOk2ZMSSnnHejTnXeM7Q5hmjHfHp+DTn92/bvjXU
iaYs4JdKO+zzXd8zmsZdS0nVd1PCaXcoxlyMuCGt6yG+jd6McTp2R+g+zvZb9/3G7wGMRyKMabuM
UBShVeIlIrSbxQyKMktqw5ZVCoTeGbqx7Yd4ESxN1dRpJOaMvATpolLROX75Uj9ebQfZabpcNg0D
QHXvUWK/nyduGk1vExjPEUdZuh0jO6KqzvLZTq+tIix3wCeM6FDd0kF12ncIMkLvT3U4UlxUL1fX
GKyVeA1faU5dfYVuZA1zQOIcXQ5rozp7uAKObunIweUoKM7yjGSxNpb4Vc+QeUigK7KhTn3q5p1i
yKtxwcZj2VIWMuEjyts3dhNMRgAp+Y+772kfVEHBqvZOQ7L3EGJafUMbzbjAWJopP778NFOx8Fvb
u2QgHwDjdCDVwlV+obvB1ucnFjqOrjymZb0fcaULAX57Nkp3KlNEQs9C5xhyptRFcDBtj9Bxzjqq
jfrqs8vMZyPoz1mw1JCJR+XSlsffSbuwZVTKL4nEdD4Tk+GlS4xpOWWVhFp3hA3r2HtqDPHidFv7
z9BhKlimebz21dHUN+VRxtwND4Qx4pGOQsChCplxecUfrkRuWni6KdCuT/sFsyrCvMSGCROvRQx1
vshLcrl1RvRWKe2dxFYuOHoXtV4z4slaazEdnTZF6dhjGgw36RNXR10l8EFrbGMOW5uucUeLl6yX
QiSBlHyVIQLnzhW4B9q7ocdFseROSaLjtrrWQVJe0iy0WNAvfFSjWOxf6CCKDJz8dduCchgBRzJS
qPcbBgjbYTametJG2HWtHRh/b2TjjReAMzouOgmfoZkM782BHUMyXLM7PfUVv4l0riV3mkwmPt12
CBe7oUAfFhtAfxzGhEcXhkhnIyk50X25FdsseQ+xvLcD4xGtqv86rp4349EtijPoMLexm1RYJ7sQ
NCO9Z6AlaDhGZbZReHKyTUEYQsWu1Htipv/naPdtZqtwWbDUy5BsIs6HCS7H0COvzyxP6vCcyuQn
PWqjC/DohFs65u/KOQbjQkDLOt1ZnMTNgWpstskDIwVh5DgXJydUTDOurgaH5KZMWzF/oKpHv0XF
S1EZJAyqxURHSWIKinSbnLVBSycxYPdYaLN2yKvt+tIBuT0WSRpceACbOfF628Ull1Uw6sgYmh1m
ws0aRmHtzQMpjtbgWa/3ZnYmGCOvnHphEHQHVEDYH6t2U3hh5c1SiPXQygoYqPUiUtYMHLk//LjJ
fiytgzHFJjyaNH/HufuZdtfD7W7VspU/znpg/J9jR0Tbdc4IOcPyX9b8WFUoxPQjSMGqQHU8/4WJ
6w+2HLzfWW8baqnfvv2QBUO+/1OOX3sMYPnM4FKT6Wd0I1cJ9SYSzbb7eippxqYPTQ3Unz0xsPMZ
BIgQLfi8D7lVZeH/BX/ZchSJaBGN9Q8Ra14vKD/E0f7D2/mlKZOiZiOFEN1bUkeptvR8kaV0ihX4
pV/iVQnWwFf6VHf3LozHPCE00HkSpfs7uxjPFZk3RDVcLrOCRz0ZewaaWvlqNn83N+VYwqOlhrHy
liXO4iND9QEYIqM8SrXK/3aLCGF+NsyH78g2RiLL90AfP3wSP7mV//M5X3hbstYlE300O/URUvOu
oNMz3Mta8r59yPYhBRjb6pEXXfNG3aqKqGUSbNmw4nmDc3ogADoiPeIRSCAa3G1SMLOTRfCgUNKP
t3e93f1MeIsw33zQQb+X/4nL0uxJmWv8Dk3qQ46CTdIlXUOo9VuUEq83xudlCJmVKJYUw24RpJ2C
Ot+Q3kTit5X+bCOe6CNCGIPJrc3F2QyywIbAveSwgx6n0qz7ktdDeatfeB4P1GR0Se9wt0quyBzU
LgG/hu5P5mikE453spQUjPRYrMGipwysPQTIOcGpbJvocgZhEfxjFJTCHzKkhKtgFG9Zv9dDLeab
9Uuj1n4tW/DqPEWVPbI1JF1CvxbpGjiQdgK7YT9l2Wqp5W88Xk4HX8mDc65FjkRhpuktC9FU/rsh
txdc98PgZavrPc+lLn8aBK/u6UBGna8ZRzQ0uchuOr8WLu/MHpWJT28t6f0wN0/ukt+4dPP2IhqR
c5bQynyIKXnEo6bl5zOio3Dptq6wRrSrk87WFF+L+NZJ1QJsS3aZPdZ28VSB5LCC/hSlSooTPu4r
1ONNkWpAT4VBLwp4CuIkrXimNZz7C8DvBZmIPozoWM3IfJuFA9v55n92wY/i/O0EfCPWD5/hMQNR
3rc8JBLTTSTIXiECMsP//RdFhFLgWiyDc4ikg589gm5ZxDv+QJbKrLqT93czv8l4tRBoP4uvUhRQ
Wp6fBAucpD8wmwMUQzmTBw6dEGHFxzccqpjnbKz8JRkpGa1LO+orQJ3dJ0hGXRqkRGjTiIwUNTDM
mzcDXhy3WDEj8RTt0zd5aKeMERKa0ZX+GCE3D/QMeZ23L+6ke9CckUUOZe/aphIzBigHIvEfFkHy
jZ8YzxPUMkj+wHFzcUOBl10kjM8c1gEoBIhYNAGyf6Ji8hXbg2+Gt98BObC6KmvyzG7h8w2PjSE3
SlsK2GaVbLzURI4P97bM1cgDGQerkxaWQ/IyYe4T6I+0ngGJVwxjWMgLWj45+AbwZ1L9TuBE1/07
k03BQf7xzBttiKVNIneOvQ7XIO2BoU5aObcfonK1KHe/fOMN8HEnOLCsO+3SS6gdECkkHiwbkTFu
MgOdSLwdIL4fxjdIS3T3VqJi+WBMSmp2DxaMi+ROnO2MF1PRPiEGHw5u3egK6wdGWuKPACXEJiHu
gdzv08nzb/VKbu++do42vu8ZBGGhGRyuwFEgKnX8rXvXHU4cNxynxijX6yhYRA62j28O0ffE+m/X
rJ9AQomUS7OXXvk0PKzUxw1lSmsII8fJ50Lq5npzMnAFJopihRB3EI2EFSmDvecAKtnzsx6z5sV3
sZ0QvFMR/466GPPjqizD9UMte1CIiFnzE0q6y99XL1jQcwujB8b2/AxYLYNn7o/vkIOrt5AEQnM/
lS/HOd+SK8EdtPxCtUFGpXBUW4vtyv7QS1f7z8Ld5wgdWzt5SufOgYJ4NBJm/E86fjUJK6RH0HCs
jz/9shMQ096DPbdzVdxp1IAw/25AEvcH5xgWhByDZdmEY2FKLlGSewMjdaJClMr/hmZIqq5c4gRW
+beDaZ9ktWxwzMsK/RGEL3L/10cLdXCjJ5I2o/LVrQviupq/6dCKBvLXXfK8j35ZNuql11sSkGVs
8nqieqSUBbhL8pmqnWZPWuGeJ5imd+z80u8SuAAFCDCTTDXx/mAvoGaDcTcfI5xpko22/ideEUGp
EiH4Z1Jh5R7wdc9Grdzy9tbzEV8Lg6J6VjNwgv2+x7By7FLW5Nrw8KSdBnSKL0cc3ncBofBH361B
mfblwzNegsoPOIpTH3FJviDqEBTU4P8FUwDHvPB8dm7/bKnHej/E0hXCQatCgFSZQTVI/eYD0mVB
ER5pdNNQjDpz/v/5nwmPP5V2awSf1UpUj903oGxOeb3LOihwoCo2JaIkd8y/cYRJeX14vFWQnrGC
GqtN00eDQqmUFxHE0iy0vFwqvw14AvxoadLCmHjrnU+NvquJcJ17+VXDh8HMqaFzp0RueCDWFR1M
I3r/Q0dlQk9NP69k6IAn2nJ+j7HaqKnLjC6/iKdBGyfUgy3xW6uMk0bJ/7oAClQIsHUeUEQKmK70
kyCLVVM9gQeRMp071bP2wEmhzKtaVIlfVrj7aKOWhjj6MlcOHJ2U6llUfzTrywCZHcGuwz1iKmpu
7blb1wb2lupRMBJeTLbhr/2walidKKFN3AEBPm41BQEUW2ZJVjV2V1PVCitsX4xeNgJaTi8pDfoB
On9ja9c/zv0t/Uk6h6ZsfMz9qeyvV59K0RWcxIcs9yrUcPqmb+mNiouwggb6JjPK2f2sxCnFECq7
ITtldh/zDVMXCHgShT3T8Aprkkrksc0/Hk+q23K431/jlnKcAaKqkc8b8B8wDcbmXSlS3IPQQmt9
PoT/4L2kd5nmgdZisqqUmi1GjLc+XXNuEKgV91StEyR+bNHzFnv+D4QRAJT3tblnx1exVh7Snc41
Qu0jy/xOqUwA+RtW9iY/AvMsp1pbjO839mG13OrYu1zrBA++j9C73jpqBoiBsypEecBzGPxdgdxg
mv0vuc9ZSB5mO8CFckxJIsAi2u/6PiUI+qXFSI4NpqgmpARaZ4Jhln5ArtJ4ppZB+Q8qI1Baaae6
xG1ZJ4ydDzYZ/3f9D/38BQWmA3EaF4K7n/hiY0Affo56a85GenwilQiRxJqoapptp49nzdJFsJMv
aLdBSZTfFAgka/h5XmgDgmmNLhQZ25Yw/7TwF0FOEx697RrRtKmzMJWkBSsMPTdH4LqJmRIO98pe
yttpViMt8za6DqlqChK1tN4mbfXmPXQmBtMldXSagDoBpLiXl5LooFY8PHsDcnT/u5b9wDN1CVVj
Sv5V+Atq3TS77sMSOHJH91EgsjGeGPBvCQEwhVOg7HguQ/aNd6Y11ETzxCuxwKt/4wRnmImNhfoi
POoRdlTf3XbV50PWB+VD9yQ48WLpOhYC/sML9utVWEWWXSgZay4HjIq4IpGDegyOgNofiSIna9eY
TMFXDwNOqbuJAwo+VufJBuxZjzYYVp/Cd0h1M9ROciLsGWD9KD0rWlPRcyLLfWjUTyC8P53PYwkR
KrlgXKQMxodNCG8VojRvHzKL6tjFk4C7DenyIF/y0DvML9etmgUtSstUaCu6oatlY+GoJuHIoa01
2p9aXCx/3M+0QI28c2pL7DfuqmtndJh1hdz3sB5wnDN6RkUCJrEkHPVWX+tFpwa4o0ekU2wAkZRy
VRn9OzSNilz1XPbnFcK4jJL/Fk4I50duvIMmiYT7+TtZ585yqSNP9ZL5Wum20hWC9hMDhl9FF2PV
LiZtWK/BM8t73X8Y4HW2NBxc47tO/T2TXThmOt1gA5Oz7QdUAqJf6Xg7L0/hLTi4pKDgYT1gsO1X
87JyXi9nrFVYRoj15k0nM1jQkjGcGiG+QgURYnkn2G5HFh1JntLAxEHQIzhyWjbDo+Rj+kkbX7dQ
NUxVGmBvxouUnMe5sf8MlbW84MSrJBzePTUSwbIpzWCFRJLQwuMW+LCvOujIFHILY7SKvJzzDaud
IahuIKSBUmr7ex20XtohhCjp4hVL670gAJm6M5OO5GM0naNaFYz2Fi+OD+Z5iftcAoc72h3fDqjA
Yx/bZDpjrSoMzWm+jjtX5sIVOiFdrhSEy0mRTAGnKACU8FX89U6p1pMp20dU8scrp716hx9lZJyD
gECemTRjDxZlDxCg8fnjzLWbZn0mdVZL+LBlN2ITvN1IyJbmkN6ARiIDlgI7xzQFHPS2bKGFOzWo
HWXNZsMbJ7tw4lUnJ3xyrZkIdtDB7J+RB5+YKNAmPtCukILIAq6UPLQt0WRNMNyvsI2sAktylY+e
ymasXKnFzHyhwPG06jWm5HtWzl9Usozw8WFBHCNRa9twzPpwgarpnCN7rwCmwRtp5vS585H/DZLp
G0Gyll4ka1Iuh8Seo4/OWlO4EOcRFBUdYdfbf5UPV1UoQuxs6SRTiGGXvTc7AZf1cF0DOf8BASJ6
2VZ5V77+u3UtUAvWbx627TfE64qY0FdjV88yY8/mzlDRbGbkZOyY+fCAhy2SnBtx3rqNsMZyifH5
ApT34bpAld4bwKhaOHB3oK/09yMTcgZzMeW02yeajOld+oFQqA5MY864uo0wsCbHx5ejCXK1CSzE
TqUBn7g/mcDTpB+5zn0P8dZYdvXLkbibwUk9qnZdDOOgUiS4DUcMu3SiCbXOYBdNQ8HGH4roOTzJ
dsPBu+MgCFqI4YtMz3fT7XmleFfR1yRzc0RjwIigdi0z4CyqvtvsMkmajhAUJPXrIxrYGyMFDqrJ
FMP6RvQECVHL8N+We/KdCgSHwy9yc6I4RpUehO5pp9spoLFu465QJwuQdzpgSGGJGT4+XHvj8/M2
GD7IFQ1J+N5vRTNYo+TC4rIo4VrJeMt8kzYUrFEYqxzTO+wWGWxhNhmvawuQKk2igvgkiLnBJxlw
tbnCi3qjgN42IcGm8oq92sbHZWb2SahSYx3DKEMbt78VjaD4uzxoLJxDgZYUhYcNmTCTnMgzHmob
BoRDmCI/ivj8F33MspjoOIq6at6mUZG+Q5kvRyy9sS2IY6iiw80payc3wCYim9x7ebiMGDYxW4sk
xfja7qV5NQvRw+dypMY/w2KZbwzWj0Vx1HDE9YtZu5Pd+dtGByCMXTuNmm+oG89MZchMrKojQkvi
rSyrHC5Oaz7L9eMaBGQrVR/iYeO7q041SS3f4wF4Qwf4DWFNSMirXsrPO+tzgRiAYCWeiaZvmEaK
Q0gPIVvrtjlp1TgKDFsCoyf8P8kEswelbr550FEW9K0CSSX+k3GAMxAEdkrW6eAtknpAs4sIKxlL
PEefRT+lSUd3kmyhGk+SlXTXW15zv5YTLueUesWDCz8herR1JILDsxcpIRINCzt11rnCEtb6AZQ4
/2gT+qqe2sJSqAINFljVR8eLTmRRanmPaM0DoCEHpjmD4KvZty805uh47lairNu3yE3K9FLsuEKC
sKtwb8okEJxLfijApeMEcOuSHCWUQqOJ21Z0XuDVBVQQAlaHli2Q6JvZjAyaEbeei0QccOo4nBCj
9Xx2ND/Vcp3K6utQl3fnEsWjMfRBtJy5fmB/IJXurdXT1Guf1uA/SpgBW4NQzwl36fo3zyPG2RVT
uPk83d8SmkbqmvmTyv7Ywi/hIlieIVnAz4Q6s7kNnXmPWR+WvhL5dUoX7gy03bDr9aUpSxihyd/h
chJ88sBS3lsjWcEVKMdh5GbdTo0qYSuyM1hKV9PzV2W9WeQiappvkKiOiOvH51LF4NvmfIN2uW+r
HQaUf0ttnverGaHbIn7RyRUe5Drq4A0oR7L3aHryxMWlqh/Gw2hXx6oA0I+STiXCwmT9oXcn0cFp
2uA6h4H8bj5UFRsN7KF27oFsVGEvas0UT0K8xXgzykvgjNYCcYwHEJRuttUCnr8W3lKQ4xdGNxsP
nw8f69sj8o+aGVMI3vf7DFYvUblSDr/0dES4anzzPBJ2OYLOK+nCH3pNARHWA3t3aZ++o/yFvHYP
YpEkj4O0yEGsN0Et7K/PMrgycoMWv4Bi8t8b3rwELmj7bI6ogrwp1sUyRxDHQUDbvLdJJu0zr3P3
bxbfHLZTOmQYrVLfRTyX10wtksZt1Lhm7XKQ7VR1Vi0ZFglN+b58GoU07pYsylFFOSAr6vNHWQTp
0L0seo5MWlwDZfp43mlnQ6HjWkYphbUrdgW/vem9NtcV7P0AOz2dOBrlwnrV7+Bw8eADtQsGuF0j
8TH9+RADK/8uSeIY/o4BzAQgjhGCdjiBK2ty1r9h7uvnScLjTEJN+KNKCQ6/J9utvDh/BgcybWrQ
pJoXGcKRSD/CZuTKD3NeRCqKsKCnCjg+2Vanvof+RCHf4UM2k3VjN9i97yYiNc4JNvluRk6VQtk5
wlD+tOsuLw5xv0UJJLiVY277XdbTHalf83hiI65+xJoaxs+9JeC75JaVd1aj1iF+ZrV1NfE3I83u
AGnsk3ZOPzHSsRTwMgzQA933trbcyx9AD7o8/z/+bqSZ8w+47x5J79aNfay+KSGUoECS2f40FKeG
QEo+kHp+sFXiML7N6j4sD3XT03Gjtvs8l8EodYAgWRYjrPCQSEQWOR9LtS4RxnsHO4nWUfGkuBfu
0wr16PBBiXLmXPkucDp4cj/wH2INauTQXs6/0y/Rszj7kncFkXpDQXEs77IA0XLpfDkvRLVKOy1Z
BI8nHaZcmZrNWKZ5S1MG37UGbHYRsKHsrwfcJnPhdDeoDYZ5QVs6SBxOyHraYGURp8K80+Rymy8W
s5kyspTiRfph1eOkYc3rrQUF0nd9fiH+r5COsNnbjhHoTQsp2xHlmDoEIlu2LYAbRl7WUPHCJBAc
cASzqFAS5cCCOW1OxtwTCkhdw29dZAj2I64ixl/Op0i9nLRTmaW2jb6VlzEbeLLofQ5kjp2w6kAX
5eO2nMsQfZMWZ8hRo40CZ+n9aJ0/DyS5jN0R2Xstts2rrrsx+NB5jzTMlbOZNxgtomU1GfbVtiRB
r/msCuD7bUNt0EVGXPCmai04i2nq0dZwMve9QBzS5IcK+DKk7LvxrlPpKr0x0VxGgBfGED8t+oEN
ArmquH9NnoQP+XJDPt0ztUz82k7Ri9gzCz9/IhCDWbJ4iu7xGneXaRC1RBRWiZkp1AF88uGq9kUM
se706Z+ISQAXii9VYQm4m6xheL1m7eystPiLEOJOgHzhW61L5MGj61lBchb114jfpetk1wCEqiWf
/UJyttgdB12a+wiye9qK83w/dMRGRXFFajfqQpdmUPgp9JT/beHwg5PENQDkZ1U9n56wDdu4tn/c
XYP5WlVMsry/eP/+eEg+eesz+vfc76pDPHox3kiZpcQzS8Z/xmI+yfZIU7y1z+RCMY/en80QKMxV
zUsseXDcg4vB51ciY1UniYfdyWCYB6Wy6xV1MOF71ynALz6DXayvMyjeRjcK0GfBIMT5+FgvxQ/a
u0QAT7A2JbubS1XVzZK/jZ6F6FuGMDQcHcFqjr3aU72//WlQQgKvMy7+ojCQSJW+7peODBxIpGuW
Z7JmaBsxyvUI4hy1fJncKW8MKBqvW0fNWKkQVR0JeL2ALvLPyXElYU+YVpFcTQvAN/6yKtWlIpEn
HM1yNYqb+Dy7X8LdbxoU3C738LvWrmGVO9jxwlC3aGhB9giLg1g56ooxgZqtEKAtypm25jxWkNGY
eYk/47yxYLcG5gnY4pS3oWxNoKYOdqt8RWs55e9cVoRO5KRIkyT5zXzkUxHeapV/Lil/lF2L9KDs
hyC0VT0Hyc2M230uTC329Fq1+2hDhjelwD+hL6eBRcodDqn4aQQQ74k+L+UlgxUI1cZMySD1wIya
OS5KstOtPig6S80FE4V+NfbRKdmH1uoT12jXuB0vDQ3plG4Ij3ekH2c+xKN5JbN9IBgA8f0xnsJk
VEbjqnClRNeILUKJ+VJbVCeKFmK7g/Rn0mnHdlk9EI1cepm0IXYXbHAxcgu1Okf9TWHMaa5HyVGT
Egjp8FXZxRqM1ayamSWdlfW49lTxc/h2NM+idkTjVKWAtn3fmYxrFpuJmrp8/ZZzBo6nuQCkMiFw
fESKYCeEzqD0+iWFTkWhnbl+hbhNaJbpGNJvruzsgl//RbMIyhlXx++Vq9GLjnIRSpKaCzO52GeE
sVMQlMP3W0pFalLYjR/uV8Zr3RUW0wLwOvlK417NBfped7MRVrrgq20pv/YJI8BrAaY3lvG0prL3
8ItcITE3jFdGyxF5dA4w1WfYULo0Uc/+EfMBwLLrYYGk9hH9yR8ZedZcphlXaqnCYkBi1pnAnhM9
GtKQGiimrKBUHGJcFYE0iUE/R8uBhell1H1hF0z7iB0swrI+Lf8rOsDHY8YhsGThCZeSSzwQxsWg
KG8yTe9NSuRtvE6gULrVnuDi5mwEJoykepTy89b8lDvqq8a3UikHuXECjY6FaOEjSbYuq9cjWEjM
3c16UG8FfE4EX36aOVZWX2bwMAjsuUqLYo0ipzc2acTPlFp4vZiOZV+WsBHxwvFqdecDTVn1TSa2
fPDcwyVgMKe6D6gTX2J4k8wxEu+qaV9vBojzprWnju60qEJUGBEgGdK77+ZY6yHXNyK4G2nEJCLL
KzyT4qu4tnVtPOpAqcz/6JlzQsq8kYlw8TWgPwS9HyHZQMHiE0FY7arWF3Tf48jyws8Ku8DoHtQk
WWoi/6hjPyh34y9dnzB+WOgtnfmY1Exb7CIesDG3zRWd33lmO4yPnoG4fNPhTe+xEVwdLMoNpYMe
6MKdsUwNYjscws9OMXUzJtOyChlE1GHDP+HM43OgBRjS5M6fkk+g4ZgqLk8pKsUaV6LRDBHh02oU
WoD0S/55IHzS+mlF7nk6YFJbdN34HHBFh88eR4um/Chj1rpU/SkcHNcw8/M6fzgjj5PiPQTo1cUQ
/Dfjnzruar+4vjlnayyWeDHZTLQxwLMAoiA437bnsNaqwVMMBMD/WycYELeMJCtq/+3ibuyNwSjD
jEa3famTUm8Ue5y01ayhZ0vfV4JM2e9yYxciYOwwfYWI4W5hfp/xzu5WKkIKrd9NrrRltfapJjwr
pMj9+coUvoOPg8oXg/xeUHRC6Y79lmyFTafYOJWCuq0YLBB/HQorhagdLTLUzrHLhiVzBKJH+sCd
N6qzJH7NKBlXVaxYghe/ttq2ZsYKJ94vmTRKOA5QPGT6TOY5t6Mcg8ah1mH3tvpdS701GwCrs58K
GM05lco6pd4EGLPniw0NDPh4GLuatd0ywxqpIMbUhtzEbQY/bChueGbSHOHk/30Sd8yVVz+Q11BJ
BTRiEL4OUx007dD8UrcgijkSzKvlfu03dK0+N8km8mTxXt+LxXQfsn5KS0NvsQjXomH7iWdFp4nH
qW0aUr6SDAIay3P++xHd4K1mvaHTquDPZRuya1fHgQ/cvq7kYxW+M4feJN5/qCtMh+fDS/J+EAD4
pqSX9BIJw/sjUsbsEXWFFktCkNHlweHkNpOVjU8DH9ughOrN+WgJKvHlMVaMNaq0Vm5F3a0Sq8dp
jJFaNvVv6ktzY7ieV0a5zII20PO2fRBrX+9Cb9nM15P2relMzeaasmcJBsFxjYqnT5ksGDqHQ+j5
B3NHswbBK3uAoBjZMDqXfWnKNdqVeomeslhavqEjSxOqycSYDHk4sNjyxmi4dCVp9/TXdmjtmd76
PVErrgsZoubLNJYu5oCQnnnU1tiOq4fYZnr8Qu9tyntx2nzzUyU1kUJM+iJCMvrA436UsZrSkR9v
w5O4L32oA0B3QRok0Zdwtmdn4PIMQq0ZYvFPCZmCuUFBBqawwDis/KHhd52ILNYJnbGgq/75A2u6
itMw82kYHmuZtKvbjjORFGgxp4XCDOuY+uhM9XtampOFQjCisDbsNLrWpISNJySCjgQs0si9//Cw
uwK7s2C/CXLK50Whn/eWMRRycmXMPVdIjJUvtjVmtVpyHm6hfg6a5Pam+caRgiZuwoPrvVexKTen
z1NNMXswWGhS1PtDjizrIAc9kjXLalQiaPMSJJ79SFJrQO58YDMDHM5HrqK3WfvTDI0u4ZZrefTG
57C/HORmLq3PoBQv+PsVMdV9Mq1PQWZ0PksvbGZtASsOEvyqCW/goA60yx4bujJBqDX2PyyNXEya
/05PlZ/lXmBxS7hMMLqT5RKcDs5qggVwn7YFjByCYMbB0DJ03mtI5PC1pga8TQXq8bEUDR7DlcI7
JuwGFTA/X8l9zHqp3ga2NuimA4zPDpmIboM2FIIDrKLVHr/UiJesrCVLJfwo5Nfopecx1B+LP0QF
mj35KQd0uwAyN7OczT2VTTi1nXFMUFQ7j6dQsbk91tO64XVbjRfWvYv92H0ZcqQt2EQxHGa7VOEP
sqvRRJLNW4KuXdI2uUGsuiZemO4e7/adBB+2zEratCiPOQUwZNfDLCkHTNERmI2cVC479EZP9gET
RTj5HvlXfTv3vb6Ov+32g/Y6Bvhdh0PLT/HwIHKknPdDO7/DpK2WNJjoUuVk6PFcqUnsrvHrSqPv
4pvNeOX1OqEAwRTT7LOFqCMR89ui0H8NEilm8Ax8ACt2oBC5Ypt1jryt3/OspoIa2N/ws0AGtVxb
Q5AjnPrbCABwL/LLxyNsluscUByy3S87lMWgs8jg4oSbxogMRHzZ2Gwgd4tEpe8xbsNhy3AIAOhz
6IgR/IVYeLJ7PGGQ7GueAVseZBA4JUt252g9rEI0YMdzNSO+SK0pjUJmXB4vKQIFXIUYZ6ii7csI
cdc/Ixqc56Bio+5CATvHwHJeHOp9jqz4mVmChitAI05IrDlUfVblxSbg4TqvrRnBxwEvQ+BrxQYI
x+tjct/zL312/G035LGw8bhFUiJZgUIZ6+2RZuZyfKDUo93h0Rqr9I3dwalN0z41kUJTxXZ5v5TZ
03Yaw/ozg7zBbox3qOIj+YQlknmQko8TnyJYb4lG1cXIFqro2y1N7IxbPfuvbdjxIKUHp93ZspPb
ALhYOguAIsy+wHXiIU6cLWCPKFNWE263ZsGufR4Jg4RMuwxrGrMwUDjqRFcaYe6uQ0sWd9VOJDHj
DVqP5R6AQXnkK6XFIzQEeO8Lkf3zd32rZ80NKKAQPR11MWaF08z1QiNFtD2g1CMDMXlLdXwHBGGd
UYeA83T8ZYD3c7ZcKdlapwjT1TyBMxk0V/2etxJQ6nTZcCQB3lucYQPjs9H5tlX9o1YAkNxwMVHe
rOLxVk6OiHfrSRtKe0iyUHp6o5l43JfC14RJH3twQMYGx4WSZHnKEpXJ8p2+xvGAcT95MP0plh/w
BhVUoebMdSUOoAr62x68g+fEHV3kEtTgCIIbr+49SMZirbjhWzQTp3qlYLZRMXwg8PQnGPQyXbsr
61Ona8L8fGmL6ayEfNp6MlfV6eIFHuJ8r//UOHHYl9aJiZpElu/dKHdUobp3DqGGP4ODKkPDRjc2
jYIYfWNaVR8z9/E6BO+8h9QM2tJIZMOfzWwDTcyJTLrOPazhxvGbr7KUQKL66w+Tj279guHw0r+V
kZLMNfDYAicKuJeeAuJ9cYLIahUPgsPV84HjSFt1WnWg8iKiTWeKrI57I3qwYl4n40FvJ83UgR/c
qaHJFg1F9TR1/quv/ej1cT1Q/T5a/wYOgZ6ly2rGZSjIhsVdQ3nU8JM9nDAj+FLm/608rFf+mUq9
bEvFDysHZ1URP37XdJ6o3R4T3i+XBRIyrStoFiaccNw7Epi/cZG0aQLUwhsWBVyfHlvRftwi+1yT
5qAsMu/J+ciygf1HwElweZJnVf5uatDEIVp0v1l0QdwZQLJhFNWl/RGgQOqGsPQEYQJX8ImVrkh3
EilYCqpygvu0kC/WbQGp/66IfA3oP1SF2gxWxa0yCcVfYdNFA98808bqbyBmcS1uw8L3kS7HCUtw
3CYNeD0Jh8Hm70cB9RWwtskgdKbhXbpNHAo3YOjioNwRl3thLZG7Smj6QApE/71L+srfDWdnZAVM
dZkW2aoB6Rp0sxAUwamS934CXotIsbYiiElkXVMcWVixL6FZHqW3CJo/QJuSiu1ZfzAEfSSBt5sw
5HmlkAK60ur1xExSdC/IR0Djq8raykrau4ATNvYRTYSDrLMyYfavbrRf6beMUczzZtkNGWtI/c6Z
PxlP/BVwjKZZTaDB3Bd4bw/7OZaW20gHCVmcu/GLCik7YybqOvGAketa2QjxG8eYqU0iiPN9NvHt
/jcQN37FSsptlPQEo2NeNH8fqvasZlKMKui7np4ge3zy9tKjcLQqPOlLxhdEYhAC1oFsTYIaZibE
hOvQhEesOQDJdi2PFaULqi4e5EiUPT1zuf+SwSv4QwwKe1X3uJoPD4LrUB5TSXyL01TKUbvl4bhD
FbeL74kCDnXDbB4qbzmC/2YJI2ptQUd/GpTOQK2z3Vv1SAEogOr8nyDQ59+ENXF9EzaysTpNZrY7
2bboqIsFDXA8UT0SKLaZGXUaSs1KbUdzxn+xYxY7SaIatU7fdT6jlSe2uOUY90f4VvZKZzJqNPaH
0YP/eRpt7/JhWaxoPvYlOuDj8lABMKspzlJeY4v2MRaf4ovJbH0xvOAD5PAgu8OVlPdkxwsqZQbZ
Lp3lyT6IxzUamv2EfianaAmPyEsb2gSASrGdsnyoZBzvh5lE4BQU9iG4onJNZGNH8uDUQvLJIcNh
BKHfdJAXlNslCH1reswBcGP2wHFr9TSUHBfA6MZJ6YC8pXaeTCC/6tiZ/r9qfM+5zE6+ATS6ri/1
KsTCWUy1nmPiBVbeFe1d3Jv7K/09vpovGqJZWovd/pdONxjEx9i/6BxO/oor4pjUUY3dA7Ue+l7f
9Zsh8z/+T6qMrschv2FAq9j7s4byJxvZAaJDdNpHBYONMbrc1IaAuQzTq9m/LYkxOGPHl47WQttq
hmqR/4Ac3ix6Dg1vClehAe2GoMwq2L5jl2KSIXme7R8cHTTHSvv0GCZzRt3EF619CUHnI9OWAEjj
QhnrRrPMdY3DfIyHV8vn3rCnaC11iCuCuRnIm2/vV9odM65gnQaBAE3i4blUSbkSnUBgaUBnBYm9
yDrpZUGEjPAvmXv6fm4Kv8TM8vg50LSRQHf9EuwR60pb3aFY/vhfvAW8JJDJpufUsUDenu+1vSs+
ZeZzb9MU2m/uwH15QbKIGdcBf4bw3mF7nFcbUAs5+EVDVbFS86qpsLkU+A72FKvCrZZNShTE2hoK
/l5Haeujs7P+lqsDictaQKnyOzLa2SLRYMFZ2ch/csjV6/GUoshi7EBDy5RQU891YtK3BAgVan7n
NFS7wN1bXgxoogBqiyZ+6OhBiWG3HqiR3Pp7i/DFSPDq4bqLzzgem+t2RNFyWxjVNZoS0Ou43KD4
oB414AdAeTTRgqfAMfPpAyJKK9qCSGBs/K0J8yjyLcuVAv558SfmWK/8q6Pb/+W+UVIVwOi+0kE3
Lh6cOZFMD9YiTvlMS3eYeo7qeiqQqtnJLw1ti4KfalPGH2BZ1Mfm8O3sqGX7ZRG86xRbnGI7hgKw
vx3rbZcTyBnQq7XZZMxjdbpS3C0xMUHO+uFduO4OI4snJMXFQEvWjTSe14kPAs6TJmlK3fjR3IQj
HWipvdhvHEwTEWttpklNk2N4059uS479qDhY7pZxQ9GdN/vG+BIpC5Vau567MyLq3QNfDqXFqAAB
ivWZqssYWQTdjEa54FczWBzD48IMqhahQ46t2monHyKo16A4wFSLn4qsCvdYOcKBSzEIrpy2ulTm
xn/gduf62ZnTRTt3wh8TW/Xutlsgy3WGwTWQM+WQOhAtnl1CDaqTrSAldK0PUbWPzSxdntmg7XIz
mu76csi0ypa6DSF6PV7Nza1iQFm6y/rqZYUo2Es1kVRU/k2HCdddN5IUioUx62m1tGUxivTIcPel
XYSnGmr9fE1e3K9u6cO3UQyWb0FQtgxiiN4vDL7kBtr7H+SAJGDgZMrT0QQER7mtSHVr9l04wQG+
FwLtxXJgj3GFdu2NgwIhrrMTmECvi28vzHc3RyRv+Uy1utp6C9QV645L0TSnm3eRvDHX7WUD+8D1
Wg0Xww7XP7QkOxtYSbVpNKXfTBdddYQWkSao2CzFC08KSI7V8bM24BGsv+MPIJtfhcXtUNP+VN5C
quUQcxHalhJqJU2oOCjIq+PtbJ5k2hN9USVBdbqmsN0+tniZlAa5Vj4ZdgvZyCf25qR0nb2tZDOR
UA8lMX9JKZIcmOiihHxKK/EaEzFPYjyKJDqEij8NF881uUKmk+T8Frcf0jOjP8JHsIPz2Ls7GxZf
T3ReiGkHduyrWJk1mV6EqHlUTHu5jtXKTx27gxur6zVuY3XBQsUYpgpGsYaLxRz8wYhDjpE4rjop
6Z3knjJHW5FUwZrE33M5Grs8e/pWapSn7UwJdUJum2K8bv7+iXxE3b1Csy8uw772Mwi81oi3WQz/
oH9wQ34AO3kclvL2u7mZsGGOt96r3vy3u/XLQvLlyS1pQdJ0uoykw5N9jQRFhQEA1T4LxNgywFZl
tIqRrQtbChS80RU+/uaJ3wQffFIrwdf/cYRaHGshLOerZgKbTQkVo5ggsGe8+KXpkpPKXd+IIwa3
pFEdmGoAUdyYMGbfRPSiQ2zMkUvpMmqK3giuooGyu9DgemEuqO5XJsxsjK6i9GAbaDjDzcY9ADnz
VXCtswjNDkr55IRpvWMf9S1ECxWss4m+aPeBVfnZqKA6JdGMRHyw9lV28GmMdZaRDzkEfZXlaqv2
Ctl/xn+AMqjMdEh5G3rb4sS14rIzdHf0Am8e0/SZrYZ9A+P5ZBOwPRxt5ipNfhRRScGQG+oCz8bC
KAOWwBoGvDqcbumTM/z0ktTMwoRiZl0SQtFRbIGb/RqbMHzah2TQ1fWOP74xWQ+VULIDa6Fmu+b6
rstK/7sNNjZYhyF6paVcHA6ZSlj8L9OoSzm0f/UKQ4C+DKajU1tEDDcLeG4lciWzmSZ7HUWwxwMJ
GFY/jyFxUAvLCTY1w/IdhB0LHsVmgw41V/wca9Fnhy/IS1/4YNZw74ZjKw1YQYcEecesyhtJBVSN
5f39pcAQ3qx2ZZBBMYREhx5ZaJ5OvyNg9eYxFAeCmUNLZXsY9oyvmQnwaiYgojPTfHW5uX8uq3aG
V7KjCnG1BhZNeJJxR+kc4Wibar2VI+1hVapkXgAfmYHVFwKN6eOXB4PZmzTiZEepZ0pS13JDynFj
RIn8OjWpE89rEhNeruzSXY4Q7xnwRyznuU4CZoQf27YASpvlTWUYRScQ+JOJe4uCn+J8K+byhLiu
62du0iSePTMqWmJzwTo86Kkea7dDj3JH5M4FrZG0PxdHNUuHh9m3kLdWiVg3E5lPIsnrejGBiaRg
ctP0++HeocdkGsAEnSf5Og25xQQms4ogt5CvHU2qH0plmPkt1iXN5MJDA7M6TfTSS+0MpSenzcWR
8JJQSo0wF+6cBGws4hmsC29Jf6JSbqUws3aOAjcmO9e+agOyuXQ/MB2dmd9RACy4FcmYubuPmuzA
En8tzp0jrHFwZN0pwSxC6QiWG6/S/Y4yiyuILYmLKysbBPKUoBiVzswR408m9ofodX6GM/aip94B
gaStPKcXsSAMFPLamm1bToP7vRX2noKLR0WuX7X/YSOlN0Q0TGxnF4A45iZo+VHl61hhk1CxIK54
umFzdD+61i0up8hjwRemx1Mc/KmkHA04ery3TnMUQdVr/0xKk01ciwrbp7wF4Ck6+8riiC5Eu2V4
trSODKi2eTtl44ED+nzImsMGfoWyM57+FaUl9OPLm3I6DSjoIjSrb92nRJy4t8jnRv8WzXo3OZPt
OiqRg9hF8G/jlx6hHkSqWYLJkoyTxELqMawgEwCR7+pG52t9rPPyvrkjGMpEZKbMSWZe2B2VzgkG
lqRLiPFkdzi8n0STZ1CwOKYw4uz5jDJsmkZSuFhT0YMwdOiK7PvTgZ9zgMlnPcfC3gpAGRing0cS
JHC1DI3fadNxqPIJIGkkV6xYEu15ynmMbcayr6F6XWu1hfQtscEENtFsaUTQcqqZwjV4gl5aV5bR
kWKI74L4QPX3V8v/V7SQcOoVO0RKfGGN4+C8Pv0JbaxasNmLIxXmrYYGArVzuHhDTI7Nf6WLM2BU
+vO+AXPbnzqSAZMCljqLrCYGZloXDd1L+5aHDu7lHpvMgkVmnMvIQMFGq3shnJ8IarOFzvB73x7p
WYZ+Z4Mnd/UIQxsA8dGr8/1/hdGMy1fUWvx/A21Vun3KkiHQSvQiwumwfoT7O222qQI5faYg9gd4
DL2c+jwvVrqExyucp/aITo6DkbSTQi8gA1xzsiuJ66GO271CyKmJUZKwGVnFCaIGbTyZ0RxCIfkW
ijIbZBlTpXgpuW5rW0vzvkKnUX/mfLUDFILBhcq54rCiS+KG+JXOUmSn98emnvbv3ou3vpkTe6ud
bXmlk9euHmyMEV5mux0kdQeEA2j3TjDGlCiJ+JdsiAdDKbO09lgqkUwcuqkT7gI69hJjdAaj6i4g
TxfytD5d/C8wC06L2+Poxmb5O8Is84zgtDrTdLXh/tgG7hqCb1vPc0ljTNSmsU44YgnkoYLOprDA
ZIbhCYDi2cN9XpGZiaz5XZJ97Bmn5cZ70nZtvlEqDk/cU1ILy3iZ6yV+G7KtUB2V/hQ/LNuGGSfd
rrLHzFswdI/tkE22YHEmsrPQHUl02Mz8pYMxlUtdr8LurUrOjHe9RCX8P6c4k/uiAhg1QLpeVAI2
iJlaHD8ih+qySFmNASoKtCHzVeohD9Y1+KRbEWz/I8uiMSWFeB3/yR4NoL/HNCFAzH/TGljAZR/c
zepeXczwNMVnoDnVeLbYtWWh72ElI7u8avWOf+NJ9f/QAuvcKddhBlCCsFpnYlF0bpcNryeskI1w
1KBnpJgDwFqnXlebGnrEz5Y9JLFXf6WphsHg7XHlmbDwqjZQQR3VL3Cq50m28WYl2A5skOWEkSVp
v5QLbtIK76kY1dRqRB3Hbv+DtO7w7WiEtTs8bQubZopxpmPfDCF+STc0DP0YtskxRrih2goURMBu
xnX6+FUMvB57KdtRp7QpQpc5h76slfPLRiFIknV318zzQQElw8dtur1FH64E0zJYULm6k0tnFQ/Q
eIacnHDtfwJDaxgp+14XCqHDzWHa0qGD9HAFqL7VfusHud0l0akEHu1G9Zoikldqn/1vwG8+xwW5
Kqf97YccJZK1gPlfnIYDz186ZNT4oR1DrhSSeROgRxD+tHuu47XSrGzQQCd55FCCvutoYlF7ReS3
n9pu8NHIWhIU4f9bD9ABzBSrPdfPyhdMbGFT725bYFG2Xc76msNaUhWY7pCFQkUbtvKa3mD5+ml9
6ps6R30E4QTKdjFkhaJQHjQlaxm0gPwXw0Ke31p1taMwoaC6wIBw2hajQZq7X10yiGpoUZ1YiUyk
sucBgpkpfLGttubEXdaj0Qc0fno9ViuifO65HTff63oYR0ngCn7cO9Bg95GzK1Ny9x80XoIykrG+
S/ZihWt3SNUgeU7m27oqs0K5ltTW7iag+TCfiCRvkdS0jOa1DITtGuNlBnl8i8ElT85TOc2x7xJI
QgvssgFRPyHA7S/3VDC5KKUWJjktQ/UiXJO7gQ+/gQbiAeeSTSw+GXfYaNN0nYCkSM+XSTnX8uvt
Z3MUPQZKZ3ufKGKx+LdcaZJkmhxp4l3wPmuXU0rt1fMkAHfV2PlykNTD7ZlsEGfxt/vIeIlmIjZ2
nMG7tTG3R2xloqZLXMRSqPvZiKoywVA+rzK9CMl4axz9px7VvTaz2xhq8CD/6XuPMTbL9w++jbLx
npQjsrQfvqodZLQMa1htUfMNNT1rcFPXsMLM47P6WVXxQZvHP3m5Luy+aL1UeMItXAU8MyoL+EZ6
ULjJaEkfE5za/v8Yjif4z15m/1dRHEV1KrKvdUC/VV8EdPdA0LvA2EwDANK6bNi1xrVLTz9oOPaH
+lbg9BaSCX2HlpkkzyrQYmNPHIyQcDmkqhAXrMBd/yvqDx0P3UALLQCPeAFyw9jfFiq9qlPEbgs8
h1Wbw5eOIPcgVaOfNlHrH9FLHEJA3xWzamApLDXajWEYBen9NgBHLtCNEWCb8z+O5lR8Z58Wr4N/
4mxC12b3jZVWWtXg6feNINY8EhjCcXTxp6k2uyYKXZe0VsDnWoXNdICQPgO608bMSkllkARB4RDz
WXB1JEM/3NQfFzcwGD6WrZkVU2iz8mDgHMu1NGI2iNrVC47qifMViS+QG5IAwsIZCymtmMZN3b6L
9m1Y/bgIjzisKJjUm6zcJkbkUHzbjoiTHJ/XwKnvpJJoZRVt+LX3eHbTZukHnH8fbPzrB8WrkaBG
PZzB36NlxGUkMssjhBajmzeCkQZQBvA8hCh9GBFMzVnYtK1/jmcbbx9PofcTLq1zQD8JxGpW2zbm
gluWwAtD6ZtyS3hDz57fj59CuaaawIRIKvs4vC4+sP2QnwlFCghhU4nmGSTMvi+zpeHXkK8/eo8f
hkNftN36awnS6lq4Esrc9XiJx5G1lq06dCkoKcwejKryFJvGgViZa6aK2VJvMpwL2c6IU3Es6l+B
NioPrhlvf0E0Ai+gkMhBOsnYjwbxcz1/87ZUb75nhyiP6HFpJTsJchdrJpqZNvgJzUY8XLds+Mxs
chUlOBmH12f5orJyEKPburqP1PoObay9AI6OUMP5r4P3aPTeav17sdZpH4itdPF/nuPcByAayNZX
SaZTfzHepMLIbUQLFAQB7aFksslqT21+M+ghnlQGd02FAH8SUuh6OdfolAfnKuQlZ9tOr2KJ6BR+
gIg52h69zWuQkc6no/EgZYU+AJ5lPaj2zhhWOIobIX0Z0Tv5mvog3aV5AVMOOCkyrIfLQ6T/uZpC
GMvOeKTQRgqE8dJ267LLVtTHqu+8ZSRLprk3NwDp0ia3Y81hGbTA2vT5qGGJGKWxrxx+n4FrfZy8
RYw5Zn7WlB7GoZ1fgOwk+XkNaS+qQ3BHEka20DuUH/jMGuN+0RAi8hZ7Otedz5nvPkfFDyz2XlHd
IvgCa47Z059Y4Okw6GTsTJYIpymJCsVmP53drhr2oYUUBxYfdzNWt16cEGutM+X8le4uq58aIk0z
vht1oghj2b1V4wNcPEaICsLtj+kTc8QetkdTrFN8sL4Rz0MLpk/Ihz8kn/EkjCwuc2rj7hXucjdz
o5EDSPOJYX3ij80dfZXyFCQt9wqsVVBVMWQYUpuY1A7nAIH7gTYw7tnINJB0PjDZxR0NXeyzpFKb
5b6L5VUoYb4GXvsri4ndPOgfyi1ChR15Wa30dGWy5X+hmAAGtPQfhXgk7ZeENItzOUHN7dQHl+4D
0vRCjjUrnKZRB2Bcs4wayzNhd+/ukAN0z+wwWFILOo1fbuvpI+jv0W4gu49kKQPEfIGRAe/HYUNA
8oQYNpgmYAVjvu3RBR0axwfaCtZmwoNRLI9D0EzrG+eIYPvVF/bBbxRHodmLFR4T+AgLBW99m2La
tIG+7WuqLjZktSMBEB8xwpvCFU0TK0uHSm1MlE+YB6aDKZL9EavAfJQLLDaDfNBRJjsq1iYRE0Lo
2fHIxeKhYLVjYBn93xhPS31Qct2ptCsqpILe0pDrFBk8/i9WdYtjyDr7gmUpXkRdKhFWGP0Tpnrf
YKXA8REfY2G+u1XT03NPutB+OEIS1qFBdWRSh3JBqSlvzMRKgLEi0r+NrQUwQOXWhrjO9dY1gHi1
t+U2xVzL7pOVwnvjfevwzJb1iW+cb/q5ZjW7QuLj24Hu3cntpHhegT5CefMgeRQqYR/Ulu1D+BIl
N3OS0Ay/7C+fTK7h35m/fJpdsuqev+FztckWBU7vqnymCQsMIa2G3kqUOYA1qDBGIo0IC8S2txJ1
o+pIJdKCsgRvWeFpkr0GDmbs4HZYE0g/qOCwHjad5F5wq3iAM3ba1eDGLFXXRrjWcDvDCdwcuvrZ
sO9gd5cRRbu2+lBcfDODFihpqlzKnNeoqZKAOgeuI25TrkpWTtFT4PPYE3kUBfvdWdG0YDpdW5+e
4PLtI1kZST6N4GZ0L5/J8TgCgia1Z/oD+mkzchF8obi7jq40fVUzYHnkrvk7qjSEY/1gJSC5JTyn
TdC+5vmXAA4c2lUlmES5DQnZPEk8XmYEI0Wzwm3MfqBtlLPgvL50/KV1AOS5H8V1/3t3mmmiICSO
YztUV2ZrQk68KrGKQ+ii6bogzk+uBsf2gO/8Squ1Nz9Ely1YRN8zVHVYygZW/Fx28xXzR2Ws3Sh9
LjeLxygQsTWYwLRV5gy+JclCuYyJfUE4WoP7PY4lznG3sy7+zJruLzirTW3Q+ZgVEdU92Knza5G6
E7lQ5272YvdSFmt6TzW0JNT0uTbN0WdnRPAMZDye7QZYaEZI8dvtwoS4BxVvt5BQ5DWKZ4cK4kb1
TPI6WneMIPI9vyo/tHEVsRdLImIWRuvJHYyy+OBw+jMuEJptjz2+GAPgNlZzKY9bqh+Xgq9Nw9pK
1RwVK3V8xBVSChVtfpsJH7VU2bpXlXQniR7YiImtYY3HjNRIBw/LTug4l99yRTDhI4YIRzyKQUf2
0/GkshYUONNovh6KhO8sDK7VS10uFmlW+dzhz4pvRlQa1JMPhstQOgLlVrlEPi+hGFdXK1K5FINU
WlL6+34O7JjOMJ1Mtox1JQxxulPHQeAz+cG7Ysg04X8GY9K7co3QOLiIlgcLrrAg3hMo7R3fObi9
fm4Yjqww3ymy2OqHWorlsxRxMX+b0nVqSKVMqwCuRLLzUlAbAf8G0lW/FmXRy83z9Ullg0H5hfGl
Igcq74XUwq5scFiogDC/KD6HJNIOEvPNtqIxnDGt4mfDb1cNky87Ch7rIsi3dGHtXTR2eup2x+nY
1N3oxvYvQK7cLIhSeUu9vKJb7wYt9Uq+B8BVJkIVY9vAgW14lxTIYqRC3WJ2ljQQ39Gb2q6UrbEd
PCoqqhawzBL73KXN0Um+2gvP1VXDxGPRx1Po6vT1z/W6Ih9p9DmbTIUOtVSeYkVvDwGPUE3WOUmw
mhprmmMqej5bhLn+48GKZC+DtH8nr0C6tu8yvDxS9Xan3MRSeoeagA8n934VjE+0O87KaXEHqHfI
DPzHKmbOQ353RJv+eJLM9QVqOjRju8VJ3z3gyxUOw7HpYGLV995mw1+KWmOGmQFgv2nb7q0EKr5F
QYgd13pjIEnwh7JvaZEd7YPWa+gAcmgM8MCO3JfxDq4oiXiCu+7aSAzpTv0vnLCqjJ7FhbZufAsv
xVELhRhgNElXrLaWB2Pe1pDlPP3xE6MtopYsGGT2kIeQ5Ebj3+kKOzzgsNa+e8x9qP7o7JBlpaia
IqsBxXFKA0iUVBgkf3tBxx7OsRyTQktdEjtkagYTIqNDbKcur3zScJtU1CtI6xgTtt1Ea+/brc5K
iij56eCqa3pFBY3bC1CfeGRH46Lo/H3fqJAuMZkAIwmSW0LXDmCtiD/OpV/nvGbzZkY1V41AUgq+
K4xOiGcVXeSmp9nKEZyhNIM6nce3hvn/FyJdPKLhbbrLXLWaHiOMnozUT4FlQ3M6sQG1NYR76HPG
oqx3Z8Fi4wE0GGzCZenSNq90ma0VMiCXZBdNKDGpBfY+y1FSANP4EquYfijiwMt2ly01qxI0nnS4
JPFmaEAB6hPfDvruETkNQIgddOREgf+HFxVlbE60jlWze46wYnafarUO9ICbwLyJxgW0HZqw17EC
Waq2P9PVZYjFNNCbVowBSqnsYv4mxZXoHhT66wxvRaijnvpHi+zxNFwwST53xt2sfp+O9pG3yQM3
6iP2uGJwWaxzOo5jiFXlCov+pT1Ruj7PHchpHb5KDSq/qHgdMIFa0nC5Od5Og8Ysc+9wcvAXuvSa
QS9lCPkqp3hfFWzTXdfukA37AjoduB+yEwb0FgybLZzqoES8j9ruQsQ2y8Qa7pTCA9CMOOK8jFjZ
m8avFM0WolR97RO9h6M6pUrS/RbCPLGNrii8a3ClFSY3DWMZF3zF+qBKCah71La8fK8LNwF3Aj87
gVEC+SC4akfO54h1T7LcEbB9CaWt/p/wJxwqvMYwKr/rX8zST5zbmCdMW89Q4/uR6p++I18+nmid
jgAEfYrKmQitemnY4ryYRRpdLhuZQbMhIGMv0ST1fI17vfidp/HksGzMaU8M9TChYMRruGOjSYaB
Emqi48P4rKmxsFRH2anHrwzO6SfC4wLSUQ7nK+8WlqbP6OPXXoGg0p7ZnASRJhGGca4lmrnt4D4A
pZEo1B53hAIAHk1vlK9RryONjoNjSHTDE5zmNI1Uw2VxkuU+Lih8yqpmVxfhaftFi/sB3r89zMo9
4xumrN3vBD+p8Ixqw+NwRxZ/A4VF/BMINsUyidoc5XJWxomLN0QdcNWbl27ZmvU5QlGKcrH8DE9p
YDEegUNBnKYayHlhpctcIeszaxdEXJIMcOq1AtCrRhMbOd7eAWipV3G7CfpO8+1n5bgAK+7L2mPi
VfqTI6xvYPFYS++FXoUhJEgomIHSqjxH0V0xtJeUn7Cf3Gkxy/VEbwfvAwIjG1nJrjt/XBDH4Q2Q
+pTa/Y/+eexvg7hepjv6dUB3cn8SUBaOd07cyV/4aTkDNA5ePlYOJWpa6tw4UoM2NrVm25xqKNNr
xiw6fg3gshslTjvw3kOO9k4m1MdPer+NUj5w2J5P+EW+HJ9jzHD9rflreeGJUQH82pvJ5Ju3FqQJ
faLRzPVWjlKTSJ0U/OlPfkDWYVjZu3t+AXLQq3qfT/RdSfWqU54xxIOZDZUMUPrxCQbvHqvZvKht
U61WOm29HsLsTbWQQSJY5KITvELHJ3E+Keu1sR4n7lmufmI6R1xYpqHDzfJJeEEwn+20VEb2qaCk
MuwLFxMuosCsWBueZtmst2y1F80VBV2JJi7cHBG7tDMbaeIqn4IaJhDgIMQbpAOqBoSMC8d4GhyH
QrdbpbnBPU51odLqIKNd1gPWfO4CYAtoMUTG9EZXe+OSDGb3UUMkC0/TLbxiDbgpxo5NyonmGyQP
ZByt/mUxqJhXWeI5XPBwXbLj62M9dbv13cQEw98qqsxsMxyCc3YOWOPAC0wnwZ4CjQdamqyXPS1x
J8X+suvx55wy/y0KTT2Ox9jM0J99SoefgyPLbilghOHDaWYTVCNA4vr98FpZPvGmChwR37CKVKJ/
Ea/z503XRotO44BoZrzj4sv9Pa9a/Cu/WGHvts04zgv7XhH3x4amju5eEUseyK18lpvJ6yFX4x/J
gaxB///GzU56SRqu51cqnVfyJR0aBsxYxYsYl05o5wMi94D1C51g5p/pTdi2ehPJzxP3N9ONMXAO
uyQz+Q0pEw0lTj4bLEHNJXlAYTLLaCU61Yt+/CNZr0X8SFOXTWeCeOxxwVoSh4ZrikVVO5iyVKkJ
tr5MZbZo++WpuaX4IctT3f/BlgmvwWG3ETgPBtW7n5FXAIZ2eAgxPhjmTUva2Jvw//RlOoZ5qtwT
4lqkHGRmBRC5Wd9VLsYehC+pGKYT6LTpN6Wcr/+Lg5tSZkarVaL+B2z6+BMZVCISbAXtp4hGhpT3
XTMBlhUK3X6e7vVGC0ewwbfau5AhRDu02deo742ovZjD7OwL8+meWy+2a91rvg0MhcG6NNCXF65f
Y1BgPHCWQdAlINkv0vwiSDFSKL5L8Ziq1qRHBcqEjd9/vrFN1/geQpK4yuboRN0tgF4/LRDH9toD
WA7W81yNMQRdHvDfW6xg1hkgV/SBkvfxi0wD3+w7o6gQbpjqAq1D0aVCkkMnBMjQXpXluiv3Bzis
ZhFdTPt1hZU3t6i0b1xwW5KUrXfpe5p13nakuOrYc+mcFA8lo8t/X5+iCT+WFjP2X0XvlEjlPal7
3/GDWU3yMST6FpgN9nn4NxGhEVpcGi8Yt7daz4MhCcbaBAFkRfzNGCbw1pch9JC4B+Q67GqbIEg0
5b6GBUy1nlMrLYrGpIcVmCrFaDiwCJRs9Wk6jJ1ESAyx/uYvY5FfDYVMn72oMFmHzARuHnoxKPG5
6rw+VjW3d0YwDSTYIKVb3l/LUmuCaPALjLo3BYj3iIyhW/u8gAYAI1uAt9T6j5kWKG5zK2ki73jj
HxIMfwPXR7ROrim1tpWtjyw8vMNhfmW19fRpvLmpRKn3KTwLFCZR19yIuqXYD28hEp3ROlLOsgHF
tX2G98VBA9qsfAeddqI7qVlONKkLBGc6qI3rbjk6FXAfEKq2KLmRfW8vEBdTnEAVPlalUk2gpblm
TgV0bUPh1T9wFCfjFCKeZh+fFsN8O1X7V0QCfLH/iZeC7iRzaYiZqa5AWi6rV9zIc8FvWlFflCAJ
hKJFzu6EcQkeO4O4pyLPRFEzhGpRcrFXrwTsogD2t1PLfVMJEyM9CUGfoLqe7hnfJNvJo5v7osxq
2vmLpe9Z3QGCabsohN88sllB98vAKDqkrWoDVYB156FGwQRT81NxYZkseqfb+bk1ZhR4JoKn74Jz
jq0en5SNFjSkIfAfY31lbhHLP9KeuWXa9zKSg9o5Qrar6HdzEOTpkma4RI12gFjbte3cnzeFuGVD
IrNRmrVuUfFZqe24X6EOSGDJY7SchCYsCkS0REf85wLSAa70rBwD2sRLsUVenhtDgVPlkaGn+IA+
QhiK699exMVQSBWwxN/o0Dewt/LthEG1uluLj6QoQ23LtnMgbSY61WLQy8PY07uhraJ/0biSgPfN
3kHh0BIVeu3w5zFpb10h5UYSWdyUzn4ELO9VRY9XBk0QirFYTP70XXzPhC2aRLzzR32UvCA8eOGN
4fhNiWMEgTdMZioJ1TWGZ1b6jiyDXwxW51MrDJLOZnEySJFOzV1Ourvriz9VRERMQjOt03rPfEeB
3Esp8CcRjgUmypLB5qFwQVRNndduXFDCs3gytjhGPiUKiM0LmU8m6lluY5wgt4s802KNndtc+yYy
zTZSbOQZVMhalmk3GcOXIUPzeryhtRt6cFpspZjOcTZcENAuKhV77ApXYupvGz3XK1xunWKXVL1J
g1N2df/1Rcc1iRANyxQCGKayMCr7AAYuU6W04oQqgvatgkHXs/txFXd90jAKJvAJcBcgbN4uqriL
OwuI6GLUpRG8b2WwkiZB3Dx+5P+slN0PIh7A3tNijRb4gfUstbe1YmiV04uNI3H5qPep/RwbLyQR
XUDmLDhCAx46NGLJzWFgsDp2AOnNlYwDYUA25iQZfyxjG5CpYWs9bsQNAM7fbAS3+y5+8EEMP4bG
P9M5lgLn40X2Bj1TA7eAMGKVpnxnKDhqeNYFfo4isFB+qIRtHprkUazXJ8WhyjSQMmBWz0c1k1SO
+Uo6B6V3HW2MLpKeR1E4qbYdOEcm9vlPkUm6TFWTW1GoSWN6YE0M6V9qE8DTmgGNEY9zOn9ePXbA
+VJVYDyQNfTNptncjUn7bwn5qVWZTN1IALpDWRhkNlEXnKDo7HdyUH6qrCB9KR7zM2X6/nX2HahM
/4rAzk0LQ34ALuQBClly11tAh/VeiEbm+rsm7GroBNPcCo41PtjR/6wKfRdz9bkrgM9K4GZxdGTZ
W/JAK52NKSIp+r6vaUY7FdYyfsepyxdWblS9j4zyhL7pnj/saPxHRkCsSvTHMRhn2Up5fP+bT0pX
gglKTU5q+meHZm4KSUjAykRc3QPe5gptKwPE2q5ll6uqI04JW+Ka11O3vq1gnRss2yx+i+aDTlfH
DjQPNVJm2drT/qmbON91ld8heaqs5LBmOkM06YqBglti/AnUsDWnB2iW8kijFeac/6fTj6VEy1he
9krjR+SFhtInZrD7vSzXMR+BeZXOhbZBCAOee9x3XSwr3jYDHhzyG6kO59LONeD+g68y4t0fFfXu
DGApbu0iLgGvGM4g3DHv+0Ua7S3zPigrlEAft8Kcv+QnUTsCoaGMfLpy5SgqcrGszRfSpvUfXvR/
pELQ8uF76fGPSqZaW2Jhuya1+Qa8hKOQO7rcgSuPJt80J7JnGF/PNplCGKYqNbJmnibkakYeeJDI
P2VxtE8gfppVNKrn5G3ey7e1xo84qxoMSTFi+GoBGRwFbgbLBxXWwIuuzn1+x8SxEcoV3tEkt8i3
OdVDWBPW7CCjT+i3ii0i8bUW2lm6i7JphcAq0dYJYqCb4Wra0ZPTvCGd036OgGrN2lFxjD2FjdxE
pnx8JBDxiYSRH7rUiZH5qEgXlUWWBl6z631DQ0GwWQGxu6XncIgeWG8zOdiNpddqSonb8Ow9jSPD
Ge+DOmgK0QVCUyfGb1w1+b1F/u12FZ1TPTvTemoPjt6TvYcvOa9DZo+U/BY4BPSTKi/xwhPlN3zJ
j2bAXfqqey/N2HXTz7PqBpI5hlR2Djax25jh72i/YFeH/Rp/JD/bPX4pA5XLKpZ3rzXVvDeby/xK
NmpQLiUdwxazW2xyZknt6KvxoZLGhBM4Curq2NdqgnFIlX2pCkYBN/NANspd63wImMy1P0ubgY07
BF56+pbOzB1ZC9WZ0MLsPuALF7qyfcjtW46MxDoL78Hz8tF/VtW4gKPqXREBfshJ+W83EjBX9HDR
DHQp/zI2ZOEnf93jfCq3KEFKuMj5CFPZr7TUqVBQdOaSDrA1uRM/Qc2ajwLCKeASpZr0z82y7a71
bQ85LgoVi88cGMdUn/bzorhnUHOilsvtH1g6T6JZwsljMJfHmqYDU8ZtCym0BCwjgvLJwtkmsxXy
dMo/ZJOvXgKfrQelanWcTk9sAVtvmau/Yp3cbMAAR2Z41aSBhc7bGws4OuVW4F/1NdrQ4n4GfnxX
8AtfUyCan+KJLcT4eFbvQevqEYNAcVbvRdjN0xvvRTHJpL+LIlNeRp7hPvbE6g3Iz8n+wQmdBPep
mFYT5oDodyXR8NWs62U5IMyVpavIEoEFg2cP/NRbHrNryJ3mtCfmCgYxYpvduMBvPSGifc5KF/St
xs7Yi0z/n0gCh1tH+spJIZqeo3a6FWNIAe9DTCXuB9p7zCLJWNGOnYMCeq2G+AX1TA42M5oHv2WB
0d/ZiXgVPOddxyGtfFcmlCnoJSsZ22XNRFhZc7Z8HIwa4q2JO7bjsoY1A7MXYWrVw+plwVFwMbO2
Vc5wRecuCbu55MPc8gwHXO3ipMrKi6UXMNWyJ8DEooWzIr+C9QWLjIOwO2Plj+O8ApKXkMuZSfQ2
QZRT+j3Vmpq/AVFyBzkv2aUwfotgSu8WlVUpurXLvgLHKtrt6XI8V2sYQn+NW+ls7F0b6Z8yq0zv
6sgrl6Zj0Ex0dkUs0rEdiYRVRbSZmouaVLLKR5+c8sCnV+LUoOXxNHn7evCY3qoBhjPS7aIkqdMB
rs4LgXB29Okyz16R4A1R8EqJuDcQoSF9tQVipvEFWihcIligesvfKZxPNGImZQD7tJezjVPw9082
S1Dke8KmNTyyBf3wp4SCj0PwUxr+XhNQUEW15txybo++zD0PqSU8nVdRjB2NTEwXC8JzUsJrGqHB
jNca8KXfR2JufGAl9Er9S/XRPAsFc8eiZLLtnxtbjtE+DGPX21aKScYaNhjoKhMavC1IRrQxlG2l
/6sIvODrxHInbwcOam08XWB90yZR/fIz4F1hS+P1psfOdzaEUdsvK558236IyH+Dj473lQLQS8vV
fPndi1dkGyL9QreMEVdvRU9BeuOkzXjAcH0zN7yU07E+JYPkIcJwyx4caP5IUtX41PMPxoyLz2hc
6Hj+miaVLaRSRuoXdXWSZCgN0qo2SJ4m19i8BsR8Csh2UEnHLnKDDuuUllv9RunBTjfJLCuuKWku
9qIR6IhpIcnVVYK0kGUJHS12PTqoM0vP3wIkfI9EWI8vkNCLJdE+Qi6+6yQhLS1joaeaYoZk978R
okREzR89E4CeYGSCJvOIcwJoXcGvXs+daWDX8mp6pBNW1z7b6KKKZ5JyKNxc9lAtDODZey8/jFSS
WpoEn6B7xhnxRe2pfOvNhxQjFtZT1tO8X3AcDymc3DeF30p9brPjqZQTgRUbomJPadvQrcCBjVS+
rp9Iy5sAFz+o9dGvF2oDyn0FnRzn3M8ohptZrq3tz8XsgigJ1pE2fONSOTYhEQjWqXeT8g0LN6OR
sPcfh1izWODtmqyOM786Ogkm5i1GgleIHMriFS6ZZ0lq6ym7vltsvBjW/m5UXy4NBwS0e6+Y768C
UVk5yIOk08kU3qEo4AlkV11CLGoawCTLbOjs9doqx4CLOK8u2duH0ZlP+z7rdFcA6xtFJpdGyGI9
9cBQWTzwGOi8LePwXkMZKi+/HdsIkvao+mpGe0gnMHxMB041eJsLzZFeUSY7CFfryFSScmT3f+Ey
sBDbZXJ+Sgf3/PISuTJ25w8bBkyDy2DHQxdkDPkxND5z1+qL4TsOFCMrn+br43TC9D3wOJ2CziKX
ip6Nkec7GH7iWD2Fg4HM7T+QJiHHvocsjG/zbuqV4r1tucaQtMrfW+//DgsBLrl9qK+YLmtZ0Ae/
jrhry9GjhmKDvUipejY5FPO/YQ60vpuCvn7xSs7oEl+6Ar8I9xvRQ/ySxIwxzye5BeiQIncWJ7SG
vkA2I/GroTfieDJMYCcC7O3nF29apEZYPGeJ024c4GLLVYce72iauKgUAh0bbMj8kG1BE9aP7lzv
DYzeOXxfgu7+Glw/mL2XU+CxQus/Ppvfw0z1xhv2y6KGjQ3FuxWiFPSZdVZ2T2NcZVzgXP6MfCe8
9r6KNSeJIgIkOJlPWWUkjkKkFrmD+sWjNXroMquRGOMODwZCWOuqBUhdCbGuy0dYJmms3KfO60h4
6iS/zExoXTd71sMmegpKKPZCEzktj2GN28B2ltnlZLm6AiWz0AhCrvashlVDymombKoHkqn3oOxP
ahoQoWdRlEwYHF8be9RPGYLh0q/Vcn8OFv3dgGRpY+ad2V8qt6J1YvYSwW4nesTBt2pHCKhvN9fE
X55IO+3+1a+EWpBHCpmgPOdoBRjb46KE3Y+CgYlIdRhBrF5u/XXdygxDPq6G4UjAfYvsTgzeDeAx
7Fj0Gidd3CcdGVWz3CqJHm0UfDGnzRpaXkMBW4usR2jD/uU9fnfcHjlZZRe6eX0bPSxhXtuBk4Py
hkQdLPFjEARzpUMYKg/vqbPMtStAQwY294KajJD3T82k+c3dlzjCAVj17hpKsEfEFDOAEhrsRWE1
qSXQV/UV6rXvczopOoil8q6kTq3NqJF77+cQrFhR6SeormEREWO18OdQdX4jKUwtnSC+DQdn1rs5
7DJIYaAPmYsagH/J8pxF33L99fQBCl4m7kTDFU01SrGtKnLCc2zVkKAno3V/Pgp2RNnObPneTiEK
w5F5DEJVj3CqmspbrDq9PtAStLlPfdAsE6N29qwoF50uIzAdHw9CDV9tsso2dBb9zYjKpLy1HRZZ
jFfiTQG4yK3BHR7H4U1JcrfqCKEKEzYhNyrbSzpfyvyl5eo16JuEse2AeuGocSzVm7KYgETka+4g
Ro4LvfkcjORSNq9eqS6h1f89rESEBFMJ8R/JkMD0fnZu3H55PQGpd5nHnhymr0UGgKk1yU2DQaGw
PhgmnqmhkDDbI+zi6kHD/OtZEAROm+kUm75DYaKMd573ygMkaETvG2MUyXn/TabZdq473RJlxmOe
GE+Oyj6KYpmZri+hi2pwnughbQzPohCHuTW5EpeqJIDMPOuLFZ6dQVK5wc0930bTjfCGjhxyFeKT
/e52kOxnCDH8C3Uw6OvzajVpfE1Gt/8iVLzMd1yD3SVoJMT26QFM/NYL6QdoCR4GcrfJ2biPSJaf
8TgpYYsf+zP/8EaEzvRyjna4o7cWZ4U3yWn7Ckgw7r8z0P7QgFrNMNGnvqdCKNi0oYfU1Y/0ukB3
vKcQv4o45e5Jk7yGhwH+udiIbyZY1sWQPr4tCRUxA000nPQPw/WSgjLATDWCUzFJwAh2kxGBEtYs
daGhByVjuP53vHvIPf3naqmM6GprvhY1M7zuC4xS0XOQcYkoci9TerjWYd+rXPjsvSU6lg11tu7d
NCli2GQ9F4XWsI1indn3ZK3rKQ4an4PG2Md1Df4Bbqw48es6BvGR2U3/QdeF4nbIexhX5Xu0MLfP
4XyN8BLBJBMJA7D6ZvgLrZtiCS1vOculMIP+taxsFFDx+AWptHlgS6YB9E5wgikM1dODGhIi+VHl
G0PuPYSnvLq5VvIT5y1eg849Q/MO3N2pfwsDfTWWzvW9f1TXiMZ4wLeLzII51BI2ghIWIU2Fvcly
rUl0XghTW2EhiWD8xrBIWet1A4f9eacTJgQGRvCcdlkua3oIkfs90MwYuDLjRzlcE0X57PawrU1K
8oPiNxhjDtRZkp4gI8SvGcbXPxcrhZNFTkePdiaIYW3MMJoXcvCbJc+dl7eBh8+J2xwNExnMd259
eX76DDUEiVLhIfP+4XuwLHzz6OoPDMeBY+7LoR9fiJ2Ss8C8P/61XWa51+RHKEPJ1j23M3FIaKyn
/qp6CfUDI1atfFyZClordmViIre2s7ZqbhbdwKZbWHhwmClfMKHbmrSAwhTcANEnfGNoBdvscfMb
h5yIKgdSsIX0owJVln6f04pouGTuU7gpxWoTY5nXzolz2EbVD9N+fa2FngGPKOvNxRKFObmzeTps
CBJ88SAiWUni5IFVvT+QFaTlObMTL7Ffzh2yNmvhVwpXRbJNaNiEfo7JQxc8OOsYXMKfZiXagX/d
JEGVH34Z6MZOhD1rAx7aLomduK6Nb8Yr7AzCyjAY8mUCfEhXkD+GRCEt/pN9XDUc/SipaRnSX40y
F1l8PnYjMpMwE66rnABOx4EIJ92/7w9YWrzEIr/P02GXJakflYA7DO67OgnZYCf84dxrIhnNZYFi
5lEJTgDvSMw6K7j2ymI8DuvVh8T9zOC/tehl+Ro1K970xD3HD5EiLvMJ1pDfHzmKOpywa2F+HJyX
hebHvz3XlLz3eput4sEmpA2hhVCO/ajkzC5lVMWhvxM9MznyGG4mz8Mvwht61CP0y/4pXPVKigP6
LzbeVfII+VeDmCpDfgsQx066feQcjGnZtbCvurN2Kmjo4MR/5xQDq/RHKffIETFv9SCwG0th24rX
gO0H8uBhyp5ag124JeBeBT2NL0Xd3V6F/f7d91kg9DocBP86SWmpP30elQn3OVpzdatGg1QWkjuU
nROf9VYpLhHM1D6uX+MYj6riPFw4VaCNl2OtrrQQoFbl/01ZQLHCOIjyliwfEqUmL89plUcXiQak
h2lm1iVSdc95NOAYRT9rP1vU2+BkIXj/uz2Hlz06L0IV+NU5RN1Kxlbs6Njntfm5mchwyjhJbMzG
FCUBqg4rLRYa5+Hlw8UgIUA9cHd9pU/V9EiAOp0xbeI6ICkKtQ1cnpLL3q5YpiMJDUj1g6DVRAt2
qgAaSzc8CCMJBXSxlvfwrZvegHGC7PwLL675Ieg34pcbXnUQif4eAmQCaM4vdXsPFJg455+kTw9K
wyIc+dvdQC47Q2TPKYOJ9jqjph8QPBd1Jv8V9lNeF8YK+mHEIAqhFAxT40d/492/j/WDxvKYA6Mj
Nk8LwhVU7P8QyBPDJhu9ugDKI3TJmTd4Ak0lguUCisZE/MfJqxGDyZ8M/phf/dYCl6Sv+FNqoDsG
UIL1+PBlul1YePRrcoFMEptkAbfAqJh3SB+57B3nA4l3cGNFlPNMFJIgzredzZWvk4dvV885CTKO
AJK9zkLDHiv9N1kcFMjCCoUiKz8V2sZ+Grz7sfvj6aEDz2ZF3ZNVKOrXehtQhIiwUagrRbt7Qxjt
Ltv9reLz852UmriKN5c5Y+q6Bh4WYbhims7M8kNTEYO63yq4FGqfXnLOMF5mj+5wFF2aFUZ8kfe/
F8TkzUpwvmqW+bXmIFsbNHrB+HdpS+wye50SQA+aH2yJF4WEcpmaE1DLeEEf8juZK4vmM8adNVu3
wNnVclsweozVe0zmjR0WpbdDASotNpKwbB6ZXadgvONsBsSScFXvKsBuE/Pzhhpc680fIN0L4svr
q9LFb3I/vNu8okz6m1I0qvS6cfXIH324yfYSrT2QixBTMovloJ1KkqKBnQYlLYsYF/StmkiMdNAr
TYLbWufNlB1+axCblcLoTMOREB4lUA8r8rl3W7bBJteRCPVbfheX7QkBuq8cv4NC0GGRuU+5cg5w
7hXd+5ory6e3QfHTAqig/2crl0ONMy+7FnKFAbnkxHz7QTgxh+JHjw+Ztls76sMXV/xz1ThcYcSv
N+O3QDUzDmAIIKsCYpaRWQegzEfnSgqxqZX1CZnLWLSDTGFR5FXiJ9JhOoWKDQJ7oINWaDOuaanG
kAinxZwfXLHXK9g/54QtzyObEfe2UWJ0FjzrKfY2ZM9qLH+K0sUj9dtXbT77y2kLy4l1Hx0EjPHm
zqG9npLq71xuYIUxR0Xe1+POLUtMeod4wZBsM7AJuBqq08/lJf3tmHw3yWRVgB3mK+zcp2kHmXZ+
FH8exPiiRzMGZOejFF7Nw39KaeBm8WONPxJc+j4azZpkjYDZQLpdT/t2+kzI/Psdm4BD+sqiFJ7Z
TpR0uVtqp9LoxUhTEr0tGn/eBomdP5FkOq4pm+MXwJq/g5yMpKNpHnABta4An7lpk57UmPJUVmbl
9Jo9PhAwx0isrPskmt6kVT1Z1iVinJWmcYIc9tKwKEmr0WqvzFOmL+U5zkuksJdPSiE5sVlXAHm7
cZiLmWfadXTWzx9Rwcj82UYFvfObICvD62sY7ZnKqQGWrEy29+F37LAUiTiIBbHU/9q/OZCds1Sj
fvzlpQahDmXk6j7pQ45mIonUUp+9I8QTrVtL3n2ytzgRUNvBTVKQvLii4+FkvM2UJuN6qN1mQCIN
cNALMNo8yP2v7M1k71zfRNYLjSIh7Oqx6Jc/3jJ/H6Z1vln4xkTpPJ0IMAHlQRN3lHaYf5vCn2YK
LmhHZFlysPQTT7Z9omWvTA2YENDBEx71TPAi0W0+VhOx1Pg8+/jyrjSNvVRUcti9ODUOBh6NN97H
lO1PGAdWRGkuM/0N+Bclq7NZ+2vu5f0mnRTfpdCNjF8fYI23ccdvF1UcWlA4PIL31kUxh2SgQWsJ
t8XW78wlhTYoowCu9nW+de8ad5rTW7am/pedZUu3tXq8IMjniK6BWM8w8908wjEJFaRUeKCnv6i0
BhTgMYprQRMJxSjveTtyyvM+jCDd7rG8bjHbwj+/6hnkBSR6nIPZKn9kwlNCF4vRrD02ux7HBrvL
mi6k4UZXoNvP4tSc5e4IQNANgXHvIhk+zRPlZf0h8MnhoGuKn1HVtLKG6kBmodXrF5pW+aVgiEyk
stjDpEZE7SFtcU6EmxxDOALoF5HBS/GtzCboOGTcdCQdlOkKPbwvC8+glYY0JW/scUl/fMjEgqAK
DAN3M7nkg6URCc/buE6sAfj5cylN0k4edAQHTPLuFiX6gdfcqWRbzSIdJcy2Cx7WNCHJIeXwMcxw
x8tXYieGRLtVAFfNeuwvh8W4CCT3LeVLWpDrXBBiy7YcwwtmGNJHSyv9k2arC6F2Ph2BYIswoNfn
CcUKHNrhLTUnrxKtKDvDGaIF4KFP0gsxgAOtBL3/WDyMYqAgLqCZS24ltsvqwT0GiXvRf3IoiTWm
m4KnAUrms0c+KG+3TIW8MGINzjxtUvN8BzTB1pGXOWBa3uTzwDzDkeO2E6sanS4exwUqQTZRNIQ+
+YrdzAqbr38t9lYo7Pp9uVO+DGqNUc+ZjdNxD9n60FSFr2o5D6oTxBCuCBkAGDswFWXZpm4doUF+
mRawW8evj8KX42RGCVsvp6hRL//d+rJGz5cNXtkGCTevAs0TGcSOI84CKD+Wd6D90VEKT5p7IJBl
YFMQStJ46yRz34W28PPh/gyhlVsrZCc/K8Nsc2rOfPdLy4Wxi8cwXwkRmMxZMSOY2n7m9jS0XFXz
ONu7HmdTFOylxSiSI+6p+PJSPRtVxtUH0SdU/TJT8FUSC25cJLWlIm/DmnY3fOGsvR4VCFLFrZ1h
ansHKxF3auOwZKQQE4vP5p3CVLv1MIWBXhucMu8nqbHvyYCSGaM2MqYJCZcwN8KShxtyq+Kry3Wh
ESvPiOGPGc0lSR8gazkO1Qwvm9PSsiLsCcZpClhVBTOCR72r5g42bv6R1aw0TYwGRPB5okf/Om42
gSD9TQuHmY5mv42QfU6aGb5iIAh8UCOtgHq/fqca+eBSni3g4bKBZoG8LSPNyA5YzZZd0JsyW8uN
PD2mFXYdNuSa3Unj9+4pAkoFd2bq0+t29shFndvLCG33T/wBb97w2rezZBaeeOGQY8oKjIKEZLrl
A4aumL7EDvFqikwt9v7/RP4552SSVRkn9Ih9okFvFnj04jCiKzTkGBpj1T2JFoC/Fba69vqkOGpb
3fJY0uzyt/+fzmZjgYNJTCi/DPof6Q40x8Tpbt5GAlLAoT1UeZObDknkwDHnTNtQg296c6Kc0bOy
sokwnjNcXnPxdG0WrL8ctZGst+d15sNKri5Hp5ZZNOLueY/22Cy1G8e07qn7PgzqSqwGdkc0w8Iv
XeZj2U06y1qDfJrs2lYt/kfdQanknr/OT+ZbnNqLwdROu8ZXO5ThGwEAiNaKONJQ3KdAB4fL19h/
DqK3ondOIafHEDb3CYJpnWhtE3P0rMId5HPjl7xHAP7NN6ZjjuI1hHWl7CwxC1P+CrpAuSuRJ+TJ
3SLq2eV3HXryCj7lHg6rxA0oHVjJrFnq6hqlUWy0yL5e6KN76Xg8KxnJPvwnSFFpMLRYvSJrXAHr
mDw+xoWARGKyACvt8TlCw47C9acxKpdwQlKCSurtyYAtnyzfA46/v9wm+B8fjWInSUYiw2sXEvuN
wH1DXOUPZLl04qC3vWtzIRR6QZYiCCsS8Itsd8+9UI1kjBVk6YitNRsNsaQvvTzGaB8oHQkk0OSc
Z3/BpZ/Zw4mQ+EuUC8mgKXWHLcIApTsaxEa4Sv5LiRYdz7f11790tE/Oy62OOk+t2ouAt1c55k+s
T75v2ir0nUMbhs5UJ2nRbHVCxlzLyDpHUDRSi9ILYaY6Jm2oNKzT7WeHYSjuVgkOYv44h3PeLjKf
zlPJGSscRS9L1AScuL7P3w4whwl/eUAzSfflBfByLY03vCIYf2ZqFFFuxk10GG0Ph9dHJMiQuG6i
a3heaQJFCRgxX1kNHXrxnzUB7JS3vacXSuQfoxmnF64IfIDFk6XFGlfuVV1XpBw3YxqGbRolrEQ/
4e6DRJZcLAK0ZMVkG/gNdNT/9afhVWMg+eYT7DWr7gjBxi/qVTenH8aDNr11hNqLIFYwpNvefCsA
R/Vt/XeZ6yR5crNz7nbu7cWWHKG2MIlnnaBgqPnGjuADpbacHwGu8yg2efjB+X5FoP4Gfy575BR9
P9q27ZfU6x2u8cPFsFCKPpnyE9paOcgR1fHS8gavcNfvuTL1XHNTtgsbmX35aAMxJ5OUC+SRZQV8
qQtkNZ5z9zqF8boa7lbpLx8XwpN0n0lasqg7B2qmCACM7uN+xfDmJ69hziVPULehkx9YJh2ztLSR
bRZGn60vwGRWmC+w15pnRj6noKei/BNi2SWc9BzOYa28pQiww/fcixAmJdBrsVK+XH1J+73tesRR
Cfd1DHYiVqYU5LcCR5SQjlikWGk91wVrxaNAsQWKv5cyknEFLcUj8NRd4Z7hoy3UFTPg989/Xb2J
9K6Je9owHQHRzpAbpevX8ROL4pROM845Y2ZDNC1i4/HIOP0RBIOWT7teQwfj8gjX69kabUIReedJ
w58uYNNT3GG2/3RnnJpj0XI3Q+lFi7Tv1b7/9YusuKxliXZTRXpB9LRg2zHw+Iur1wFKFCJNm0MK
HUJ/kVHQPgQzktCjNoBC4hZoYVZVsHA79KB02hM1lgfWz43HgIR6lEQu6idZw3r1xBzUVEzdDz/Q
7+nD2QxQLS4dAbq64nkNc2+Da7Poucg2+54HYunk3D4+OcSBrW7JRKGEOLlTzrUJUcE3dxL0iWJk
ipNTIwWJzBJ8DOta9NPYXEhV6uWjpeqA3jfrtc358coO3XFZ/1hkbSGeNJzU2y5j9lJ2b96ISv07
nzpiiVugT8u4nhACP0NsG5nbcVGqd4jNsa095Xr/3KcFbfhn0dHLFLppVl1CGmj/9xi8l+nxCtEV
S6VaEn9hWb+IiS+t9sBOhwtiJPKW/nIS7dJGyXpC/gf3Si1oxa8YOaFdCbsRhafv3rQQiZkPoWU0
evDf8gsU0Vb+UFzrd/UJ8iFgMFy8sow/emNPAlAqd+EZu7EPjB2DxdLOCodjbAfRM0HoKUkAPuEO
p4CFJBwFxnpGWpQB0AqWEXejsPqsF/jsAdi2msdKzuFD2UjSz3BFGdESdT+nCuaS/JKM23koHSQj
z0ETC29j2yF/hFxeR/ktdTR2vBXaZhSKlZe3/32W7R+mobE+m1OBcGvSjPRzELGsbCFwgiiIW0//
83C1bFrzlCvZi7v9SKDb4C3E8r4XHwutsCgbVToGcZmwwE3Aok9uGEHXnGssZQ0PwPWQK0xTxU0W
3Q8YM7EiCSbmggjZrCaUrortjwsQKdOQPAHrcCKkVdsUhv4Evg2stcgfJxQ609CDrWO0xucToSQ+
fr8Q3vadgdt8NYtoyJ6SUhD1MvX4YwpfXjkE/1gHWRRkijKdWpj/UGF9uzVgN7+7c+cpUd8tZV4R
/QSNCgFzFYqqXIbKyk92Kq6z53MaYmbqCQcFiGvr454wE7WTgZyTuk3RZ1MpjVIVpeRGpIgry9Ng
je2a9toymBnwLcdE1TeOfyDP96Mg334P2cd1ANlENl9IL6Bu060EWTWl2+tHh4Dloz0CGaH8Eaeo
JYdFsf9Fkw7PqCRcfatdSMlMKW+VQYSjWP4LJF5pIFlDXkiOW6C2eD9F2NJ9KjUaZ5DU7l6SZqNv
v2aDwHbv+srYHLaMdI3Hc/DElimKGUM0ZNFQLx+g0lOCFsq4prts8c4lp/p0y7hY0wepErJWy81W
KTQGM5R9DBO1AvyVZeWCnCpO4zpzNlOmTPbLa0/QE5uFrOXTHGxqcoyOc38ErpgBTEGIWuXL2xGs
4vrwunhaU4Xnlr1jTmvyRcD8LL87mOxkkkQj3BUhjW8nxQpRI3JkeWt1ZoqUlHXOTBzww5zrTxSM
yha8ptbF9EnYewPrC02xlZALmVV1kPYZwzj2Oyj0Jv/3/sKBQHvs2nlKQBgz+c4yGp3dsCaqg98+
Pl6+SM6NmNp0Wx6/Hko0Qnu4u47uv9o5mk1Q9JFrB1Ywi+L/1eTTx8sAEz02/4JcEzZxBPqB3ETK
q4ZDL5d2ZHZ8LBa+mIk66nMywBWhn48V0gmiz1AS0g3z7sz4It2WS5YJ7WHMofB9etzRC5C1gEei
ax5zezBHsvHBrxXio5lsAcvpGoGeVHQs8VNJWO1p8PiiC0Hjn95pvoA2KSuE5GJV44ipmJy8yxUV
ZJukLOmXgAs2UJGO6A4qM8U58JS/RoGTNDmdwQjrIxKRfnOYuubc9j8f6ZI/BGtZioOieKo/zArq
iIvvU+2aKbEoA4gSTPyddXzvMfGrCw52Hm6vjmSqU9NXXUs8ZHq1QS+a3BQNF9zSALxomXeaGknm
FdYzabs/i8VdkWypSF60xuY1PVngkvH5MU6F0vm0n55tnd18nqur7ttsM7AFku0tPR5RxZQpx87Q
1n4MK53tQ9hhPUnjCxdwDhf29hK+xnZ3ERl9+c0DUPCQAeUQ0472oCnbXD+A0NlzAFgqel+f0CEX
XCmx1TsQTgYq8Ps6LhU/F+a5EtXy+82LcIA3xlJ3xGY20rXnPdmC+qFwE1i9lUajV4JDiO2vxCWd
1yEi/76Vj+/WMF3Q727bOXNNfof7lRpZb72JOV7IYwDrpqFvvQdNm539jTcTOR9kCDwHIwOaEN1u
hra3gNf1Cmo6CudSuHlCyX42HemELGuKQFGtG9zpBRBTP9PC44RHVRKhAkmsTTQuIycE24hA332e
2Uwt6XLjDmz72qBWZAk3CfF2AmeDDU5V4nrKfogNy8FvcT77WlSdkqFQc0yHsPI7nKwjXuRyrFBy
suTBSokbMFSySGXdsUWvJwRyWlqBOktN2XbY20t3N8BSdiji9IqjSHoFHT+dLrwn3xcGaTvnSQP0
nGpw/kP/hJvvALNFlJEUTg1mCDGXR0NBk5jTBruRNT9M8VUWt7pzWoKFpmBIoAkGhLeS7RDGEQaL
Ic1a9HyZMNQ+7e5IaTQJFLHPhvxJTMHmLHNARND52V0rG/1X6tGR/mqkhuqDV+hMpex0IptVt1NY
Fd1JwXrZO9EVTF1g7cQEWDvMqgjUx2qx0tB9vC0S0y67WCbsyNQYdi0uQtD81QrdwRgCzS1E9ZnM
3KuqiLbp+BmNDWaKTLVgIJ5BbdiD/ojuDKiEpSk+G4um99PJPkJT8c7U4j+k+VdRzywJFo/SbkA0
r+GtmOffTK33yfxGeo7xOE3aEw5dbi2R7tnuJl6SK9p3Msqq2QuhFBGNlCC6zFaPKtgzUsZ/h8NH
pRttPSWf4xnIVTzpVSiENs3teUcuPlY2r1siUi7wSoTnHkF8aQ18snPzylhCiayVxObabY7Y/fvm
y50bViQxRFgPuo+dhwqFrwEvrrVm9+XE9WgUrK0pCck/rDHy2HEODX5GBKrdTnHIqzvMoEqFCJjS
k2Yg1vUI+M5j5ako/A6jdVOGvlDKZWapV18+GV0UUDFjgPtXTvHSSE+OzKj2268up6w173piswoO
kN3Isd9JVw8Exml4c0v3QzgrflY14aqQY+x86hqoLyGtQh2lizG+bjg3NTFN8WthvH0Op9gw4MJC
HrrOjqNrGGwDTnYxJWPU5q331elELWymRyu7CjvwNHgIn17i16gv/veA7MVb+16VGbtN1TqDnyid
4IZp9vkSE0VpfEdx3i68eB5TAvwp656HYoAibZE9B4raAvoHTcrlPi9CpV/+VpZhhjwZ8upwPEL7
JGCa/W1pYDefymcGf0I+YWcWPUuh3y7Ov/iF/4wbWMrY6vpGB2ZUv7bpv2WOi+hbjM2GijmSkvqQ
WtOZOFm9el5XQg40hhsMRiTDUyEMkQvGQVNMKaDYPo4qd4c+s7RBYaDfMoj/Pfk7bB2L/O7hPejJ
4nrtyMbzwfJAQD36sUz4fiYdIDg2OW+pMMjbfaUFLKOnycLfHt9y+2WA1okSmDy1qRuJIi51se3D
n+p9xIAxmI5C2J9xlCLYUDZfpICJZzkwDgA4kFjUWqJ7KW03EE6uGOjPBB/eooUrxlKHMc9BKEiJ
SLK0rtZduaKQhBXsEJBM4Ir7FkBnYFxQKaomzM3qrHFMn6LYyltJ1kYgHtkSNd0khLOIZP8fhOkR
f72b+GrQsPpOGOuujOIe0iDJ80vbpB0yF7ZL6KlPU5J6dVKL+LT05EBZpRcOEtt1eapmVv4H4q3r
I7q8a8/C2e54/1PYU/rlTY9y9C8sugxmVEps/oHHTjJ1XbNp42lEU6ij4UpavAuf7f8EVqxK15IN
+YNt+5uh3M6k837s8ZFsmyueCrArMHjYIa4X4Poqv6JhbndmoG7K0oqiqxS0/F4fm1K2uYfdev5j
8ThLiB82112d+Di1yACOuh35Z3kUGNXfo3x4mR3tsC7jpZ/FFE2rNbPBHSp4XEcYX0Af2RT02Dob
FtXMWXGf3g9OMAoXX9iR9p+UNjd99pKoswT+N8GPKWzrOkKViBJ0Ex6ws2gN3d+VBuM0WnYob1Eh
+saFEXWsqsU9s29xaDSCHzFIZKuT23EcadF4MCvPYiJDkCKEREn0JhmEdhcmWauXZr1YVgvw2Gyj
c/u+9CoVe5ghtp/iezEOsch4xWhDnkq8tJRWbv/oWuinv7IuFdefbvCQ9klYf4Lm0P4GlAYmslAD
IlFrSxnxNvO0B+FGc+ZKyLIH0aQYhlIqhkD1WopvXdmgd0/6RIgganNHds+RZxRVIHIR8S/SIEbC
m/EgVCu0lArymA5L5Cc+OS57Z9AbAzagVykC4D7wWGsYI/hzs3jbUOqxI7paV/QOGOPEt2YWdEFU
CmmVg/d62O6nUBi/Az/YPhwTF9cW6TVuVE90UdpzfGaDnt58AfFTBJ7/IGuHsPzkopTnnPx1NB7f
lFJxE4umc3lftm5tVAUruJWG/lQ/YC4EqrJWoy9vgxRugDai4+J5I+Bya8Bq8HtTm/mXNXRyA/4H
iI5455sqDv6JlY5PgXy5dw4hblO2cmdCGx7BVB+ROoFyRJqe4To+mqJJWihogWDRnJdNkSOjf+xK
ynv+jzRtwt+I7QWxibkuVNxXSBcs8DrlDGYZRhSQlKVbiCpRPeCgqYmOf9XRj1BnkldF2CZLVTo3
hWZFH5cpJAnwd2QQm+Pik8EVofVxH0OehVcaGWv5JIChm8e8JT868xl05pJwN19vB9z92yvniUJD
lPW7wJ0zerpA2GEthFHDclzupg13fvMXI+FED8yThvA9+lebND9vKwDkQfVz1UhT5jgbRHzpf4Z/
eACHc+11stGFUOqJVoHh0tHRgI0hhfyp0AKsHxPIhTbYH85WunCU8ddMGfAHhTa4lfRn1bd+GxxK
461DkW/GH5j6+j5Ig00IbQKD7Jywo8E0UanA2z5fR76sWjjLptgzpg//LUn954XbAEmr68Q+cF6H
ro3+XuuDUuYvUvkkSvQBvcLGNpT2WN0aBlbLoDVasDyq6Cu0TfcnKrSwv7SRiGO3uQN25K6rf78J
VgYcKJO37iqk0w6hWYbaETqZzJraZ4bCBSCFumXiUcAB2q05SdVpPasleHb8gIf1xCbSzKippY6T
WVmv9V4/TuDPv+UIRYgta3e++LTRc1t24L9liXiaILHVye17IWY9dIGBaVyVws7qrzuFGdGwCJks
CE+Rf7XbOiEbEOJTU4/zASZqGW4ytwhv82mwWtwyjFaB7CMopiVe6Mh0bp8dYGKVPOVcKjm5XKKb
C5gh8YWYboZJn7LTItkagWRfCt4gityKd40ewhOk3c33Wrg/nnMpo8hHkx8yZ8WRMusOVnpagiYJ
6J96eqGya+U/rQj6XB5x7g+ylvoWTVloo8Av8MlwI20AaXejf4V4JPW48RlbHHMRlD+ViREwSnUC
HsdGRbpV8KFYXI49AnJl2w8v1qXZ6lytbCQbxmpbauUj6Nu2GWTc7mAfQZrWMF8GVJMnOP87Brff
XXftsaUX4LVF+f1MFwohYMo9DcBzxFdL3ouq3cFwM6kSZHCNDmorcU4/Ds3bYhFpKSWJH2RgrYBz
p9d55gPpUNJJI+hQDvgGAEaNWKnp6VlSpTCobyVnjmrapMbKxoV/JtyC8cCXMOIj8dZgPhDcNO/E
WOfrERKdu4m5jkg7c7KbGma0n64RV/mrqtCUV9c9LGz9ztAy0W4LLy1P41srkcw1UokzFaltYHz0
bGUFtOg+8xrLBqZFooEEcEB1uUSS23DTxMHxd7iBprQa+oGejxVPBnnMLcrDPU4T1686RDB2WKMG
4OJxWufolWYpM+hcPA3o7vch/tc9W/dxY7bHcHxyr23bxl7SpV+gtK7IhK3McSX8dsq3bL46hiMP
eJU+5iM1jEy/77U200v5SoF2eZSsxxeCk2ybywp3Q275PLFIgLQwDdFDJDwyqB+tazt/4RI3yhPF
lADseDLbk5rKXzmoTLq9//GDxbCN6SiBuEvN0E9l8Bp/fEto0S38WSvHoU+cSCdq2Jv54HFSMwIS
XaQX1B5KDV5vBtJWnRbPNflBI2Fd45MqbzeMx4HJ5tkYt4HZhDfIPtumLInpY6nEKZ3naR5+ahlO
TiaEVrS3XbdRnbmODekWouiWftJVEYR9X1i/QvDsusIlEMJh80BwG9qyheNPlBxBe/J6w/+xKjy8
NAJVNQ7hfZF4FgDEVgrE20biH7t/gXYU4o1TgJzswdIutsPQ2yM79DlxLHnomLVKg5LFx64L/TfJ
N4axSH2/Rl3Mfwug22ZNliG7eKo80D9eEDsUOxIUBd8OtsEpEtGi8rUHfKEUNdxueCbWvkVP4jtl
p1BpcMxvkAuPhjltDw5rEHYdGUVDzbuVPu4XOSA1YFRvAiUCXm0FjzWjeKEtVfFKOllIkFmhAjdh
hjoBv5gADLSZRfk2bfgLDWLZ+X6X1nmDanQNI0qGwabNBqUQlCmfKpIDNOKSITt5AtWv2HnPBV5F
TzAKGbkrdhpk1qn5IjgfMc+7D8P0tSM+hPcOssZEqlTr1USVDKv48ALB8jWpA5SB3q8b2sUibeoM
U+UuInA5G6pGGNtuP36/7NQgdDMkPontulsBg9Y81jCEQ4axQHmJTzQjPc2oGVTpqjV7uRIAjQ2B
1M74l+7eyC7HFCsPRWzEtB+yMsNH2Ob0acbPWc/UrVYc0IAXNoRV02zLv78Zv5Kj/vUKCq3PjmEp
dpQPj8nkqRYhxuPJqhafuSd7vSDqGQlFbLITpXwAtcalb/u15vdx0qxOeL6ZKwlHVdwL6ws9t/yR
AxeExEV973BliRS/vGv0Hgfgz9wzTl7FLlbyXniGZXwhGuolBGWvwJB10lzsTun8/evI/MR9kZaw
nGW/O6AWWYkcsNT2R4wWtiTsTXpTngDmQ+YkLFLyuP14cINGh32m0tEO2jyIe3WT1+1c4aiFaJ7B
UZWHlhyaorZoaITgtiucXELoc0WxgCgtmmw3ENxybQF+O9PDPkA7DwN77oFuD4BJliJt8WGp5zQd
jNM4+0UjMa0y50ZYQbeAu6ga4E0vJuNF3WL2d9xuNJpSG9Pp4mXaNFldrT8CzJA0rXEmP1puBX9G
3nN/wDQNzHYwBx1AH5inn+Ham20RZb8lSBUgUPs09YdM+pMvJTSOgCjzcErLwU94sz5NQ063HMfr
yt1POOABz1fYsLk/VAoc2OnVExT+MVnFqVZHUFsbe32jfLj7eWP/uISBi8SItwcO9SJ/ESs4NRnB
AhOmeDJWhEjXXXpcaoeZ5ezGD+eJL1e27zz0uskEHknMpf5pJ4nq1RL/2rcNZ0Y7/GnzmZ176xLu
iWmuxwx7CBw3exWyYKKJ5P45JvNU3dSmJtrEFW9plugK2dUATEvEDd6B8s1AIUn2YInSajiFSE6T
bX98xJpMjNHN86joJRaNYxYtslirjsxSTOedRNvRwPV2XUIr/mgpZPa9+nSxUeVcYtwZN3MQ25V2
b72z6krQ/SW/qGT6Mth5XDRyDRp7h5/BDsN912diNgpCdMdigzqeXZxj0jOzQ9Cd/Zg8Kujw06Gn
m4St1H4lhNsFrGI+PDli7C/Y0SHspkJqBx/yV1T7oSlZIW5yho02uUSlbCZ036Beon8y/5ronXjQ
Y8TJP3wYLaVTJXAO9tZ3Bpf9gc8As7Fo/hzfoH+xW7VDb5lxfkapw2IkgRTzdm47R4IzMjEoaS9b
5SoOicR7ufGlCAzqskBZKoPcYeQelBM78kmIn4ax7uQv/epbGjShOfiZHT5NItI/l1BXLMPeptGh
ohxd70n1bdK2eqfMULj5OvB37VnM/Loyy0CFWNHmzcgHgVgUsdsd3cvuQbIt39SgWOMazhcMFskH
YGzqm6DHtFxmOHGE3h4Bt1aTFraVUZmpr/4VJOmShMETsIQbSG3RJiupqnijr2MFKK+T+0pgd17C
d/L/vLpSWvDPAP0CnHYH+AGubxzdh2TMZkn8o2lLqrk02Xe0g82U7MyMb1cgBhXnBszSlHepZo13
R1wb7GMzZmfyjsdN+4mF4zYrqOZBOqeaF1TcDf2Dh/qFthxK5SXdw82Nx5mxYbUK0fCK3x1vSeHp
BGLzeNnD6siK3jq/fCibZOpqNJ30UBPf+spx3OAQn4RqLgNToN3JVu+nGhqVtWl8ZxdrgR95VFmM
8hqRyPfl8mjrPnY9YHPwmyLlieyGGetXtsLQO+l1SmfthIEW+9uc20BvTAtXhP1lD5IkDKL3eCxR
dXixpUW5t4coCLatKnTACA8J7YCXd/N0j2vLxeFzilYv7/ohYDmk8kKigAPPZutESW7ncELmb9SF
zrLThCHCeS3eVhfuNsNgbw//5I+AOE2A1MCdtbWIjElHoEvsKHVEIWpiJlnDaknpuCxvNmegU+aZ
iDg0QGrS6RBryk6FYJ2t+biVNXhc0oQO299H4xGG1Ob+Yizsb9x7Nv/mP+27+RNsOYQbq6mMRpmm
95nD7Kc/DKEsG3L+WSFjrZHeoNPVkliK7s7C9O4P1XjnyL4ws4Tjk36yMH0nEijMsv5yIeFzL/cl
JW1N0t34Mb+opzE7oyKdpDgabdvcLyB1Q/ljb9L6kmgHh/jwVsgDYtf7Ne29BrFLr/omIh0ynjxz
PRcQ87XDTGfY+A0s2mB3QDbwBx0u5VWK2UkqkXx2rMeNphvHPiJOLxCqfO8Xx5zL2YTEURDhDcib
0cRBOdMPovRLlDYS82IhY031vdHkjkipQc/8WLowppoUomxjPLN7ePPKFP5y74GWub1xseXlmQV5
LhO6YbSGjVlPaWvhAZe8rCWFtQEYbM6EHLUeAOqzuUR9Uffn2izBRnqsoEC5cMtuDnPc7uHQ7lnn
jZ99iBkDr5R+EhEEnY3RMKpxpOU5ta7dmijyn44i0u6A46J4EBN0/2u1kiQeqSe3x4vUSnoiNoiJ
o66TmD+SWRXTsmG6fALNA0IaQe4uw6UNj7fhXjzkPffDAPzitMVNm5GyhRnJGjZGEkvv/0OAEOQl
N6c3tWiJb7peyPgFXn5xEHsj0sNeo7SlNgbgd5z1yzsrajD0O32SlzQ/ClfdeqK1RaJWWxYAp1q2
XvDubXbyHLyvYqot/huU1G4vcMayTvuU9y7ZqmBQJvC3+p/gzDHE9q1wPF+vfIWF80FaQZeGU1CJ
EFpQdPaCiuJXJWdrvLMr19vDZkACpL3UjwfshEgA8/I9+FSmXLb/eIMP9NYaMcGoMiwVXjg5okHq
FG+bn/lrU90FnENDx6ZaglToqzkUuQWBxj/9j877Cb1qgGxqLPaAXBUNRkXh40TvpZlMlzwzStUt
oJ3sIPI9rPrQAB++WkpGGUA39kUviTqW+cmGiI6rqRNNLuOqAQBMl3k6CgQK5R8kEGVNG86sy2G0
lr1pHF8WPGF8bzTfDjs6tZFfdeqeepA6yBYKY3GHKsMY4uEK1/cG+EFamCjEQDguzB/j+RFgn827
haav8YdyKNRmZmobXNavJz79s7rP2ePpegG64qui5syn0P6C5EqVeolTDzFZISS6GNf3T6NSt1fo
yUwdh3X/7Xa0ZHuFnFHhoJ+qOGxFZKyZnmdkTktraYrXnxWGcG0gbmV+a6pjK4XV64Fc5ssxEAra
puwsqmz2oeDSbVal4u0xk19zSzPIC8BTVbLbTvyCHpGR/myeA2nBEQqerMYojHapyVKuZ/CizxcW
5lgNtDcLAkI9chcjFZPN17DJ/tZuvUpdSBCbtC1Rf/nVurnELvUee0L6QRtf504xozRIlAyPlzN3
ZoKWZAVaMc0SN9ZtiMCtl64AcMKIyaY+OfCKt10wgNVwX88OTsrj0PtLxRi1IPIyP0/nynf+qftb
LTk3EU5q/YgkzhWMqSp6IRXv3lnyv1Frj3R/kHPKyfX8UZj1ONZV60o9HA0lgaCNa0ja8gLzzbk7
D/kcNK8GBe+nPyat3W7MFWqLwbMw0k+/wpqdz//1E7UxmGJFBuZSIgjTOVMI4+dF/ke4+hJ+/bvT
rfY6nVXbdrFROjVF9m4gSge1cPiPPS6FiaXnk/Aw7AnWgGOQOd9gpevHcoZ8r9GwjCVy4W/150s3
5OhPqpX9BpKeP4T6tL2O09FTZxND5bbd8VIb+Y0KcTn63Kwl4RaYFPF9j/t7+nDIDirCzsQNyKHo
aQjs+NfCon/UNj1SvDo7tb1rXFL6rrjhXT/S7SDRVSJ64jv6DHsEiYY5+QRoWLCYIXH8GqE8Nhz1
N8eDTehlOtQqiE7+AM5JthrfpfRqQvSHlZ7SgjF2hdlZvLx/Mhz3Ls1hy1Fm3sKjCXzpgYwurY+H
ryG6SbV7+tFuQV3794RMkyWZ4YMRjYjv/69A3FTTNIwEqOXrkYZq02W6q0tyhIouoYaA/ui3PUya
9L1E9e1sk4Rl1swQQvdvi0gdiQr9Vml1Fi9HkzTtRDg198YugtpaRYi9rw9v2r5uREH3KjEYpqWo
GOrAfQZIXshuxpqsF4euTopmApD08HwloLOYeZN0rHgxRvEDcEkTphhW061zTGUK2gDIS3fNIPxN
oUbGv+xuP473K7iBpDfmECeCk1yxPY0B6wSDIjcYAaTJwW7Up3adntLnePL1blGkTDCKQwBnzpuW
8aVI3uED8GOoLF5WxuLVXVMBN56GaeF4fhmpjiI31cFB8fLu+LMwkJzQU0lyczBM5unrKcufAovS
7vQyAN/W6my7a910roQJ2PvaVw3OYfN5SEUIIhMQ2zVTUbLQv742DT+SFEU5b6z1ZNPkUx2W6aXW
vWytpdC0LRHT7n7yWDt4HuRlcTgjhYnSd4xdRnAoCWK5bpckxMLjzueBlDKSbQOnInHq7mOuTPbl
5tGnVAKY/Y64xwlGBpU7zEfVYpH9YvB/WbpQYAytpJI2Ikjt0ETiirkORSXaXGz5TT4TKgzycC2m
mDj9dIrz/LR5OPuHJCEP/xBwFeLt2FpLN+k/TWBWOvw/ZIwApvdltC5jIMFAfM6YQRporDBnu9YB
i4Tjvx/NsdU7OLt3ZlrKJv0bNiCKACyUT3XZxPTsKEadtWAm0ALuwa52jrs8Sizk47ioEmQ4HZgy
9K3TBhVmbXnB2o91dyvjsnHtsEACetcVNuqyTJ28y2gKfqYVCnrJchHNVPIzgwQcBie/nZ1AcU9m
6mUyu1eKD0yapj9axqAce3xMLUC9FmwkysvH9KPeYZ7zZBmG14d+sFMN+G0pema96w2iZlBis016
63INJ0PUNkb0x/4lP+WSm0etHdjH8b4AjmdcJDqImyS3VRg4mHccE/qMpM4nsJ3Zzy7VrvRw2ZaD
iHuWI/3WhvVHWKYWOA99Y2fMy7wp6XaJlLtpDvSgRmwaicplNAgkAheCbH8l1q6EX0BLhIQo9SA0
Ln8aJXfY77JB6W558pAwjKg/X1wU9gWE+9Rnho4PcSLGLG1O+eWPupP23iwWFWSdhpKecKQsKWA3
uvWEhTidY3zYlL+gGv7PugwIbndb34A3IWGRO0KASfkf+goMvwEaQ0RyQar8sNQ/MSck7qMJTwvf
wLh+wRmG6EnkpnH6/gn1q9Gh4gsoJQSA3nEqIwWFNMBP3SrYtO+fjxlyV/jvt0OtXpKxX5MQKDpV
6rarkNAGHMXXIzlOzuGAIpbbNsLcjkosGvRtznntZ0C7U1nKyQmbAXT9soEtHMn5UznhHh3LeBv9
xV30suy232PM8T/vLq93+ZQnB1VXzu1yBoWAST8SlLX4CNdwWjmKltawWPQWsoUAFoIgTRi2xdzB
I+rSydzKnVZZSZp5gnK8pCAZLkE1ejqClqkg8KGLPJZC3uGWZIlzB2R93C5aUrekYaFXg5K3SDgB
9C1zzAqSZsDo34KWefkI+i8GYtGgMrD7xFFfK59836qVHvMmTHki1ZkLGjgosavMHgi+UZAG/N7a
bDxYxOm1ZerlaZyJnMHxyuL33AH19bzJMnAWbkuYSfkfm3AbsPoRp6pv6PZrYlUCNJL7L5r4LK69
HvVCoJwOHKbLH8QLJXlOyWqyJOXKWB8PUbBXWuo+8Q2yAdwCUHJHGZ+jJbUEAk+4pVbG/xJzipvH
R/QuquXxtQqjmyQKabzOPhdpiyH+dZMSviRl1cV4lFL3lkjaTrujK+nD2Ofd6VpQp7hXzaM9ifv0
C6QP6pCr33RJhIZ1zYoWutxQOwx/bXjqTmkA+FEUzXB8S9uymRy0Bc0O1lkiSYiAGEGgCI7cHl1C
ezthw2+FfhwImpk5GfbmVnRCzYYW9ja4X1gbdQ09tu+au5PHbh/4ATslIwqzofT3jl8bWz3D2uL2
TuivklRG3FA/QlM5bvSWsaUjw2RWURt+kbLZ9aIkBcIDXj3cb7F5ZvWEM9Eyzu1G5UAosoVsAslU
si0vDNPzQvH3YQACkAJeBogAVuxJFx7QA2tDw2PEgf82nmO+VFCnhtyskfE4iFNpwS8BwPvmRhHV
SZcw9S1GO4qp/4j5vhrNst6I5kwCoYGHzn642JqUj4fNeB2Q+mzItntORec5GmRjw7Ci/loBadpA
p8Tj/e/zsk/vnThppmX7FH4scSCp+7riIXDtrOP380Xkusset99PbcCp23amOEXF2dYVA4pQltgx
3Eo85Hr1I9hTBKKYHLyefjogb96ogfClgU1g1GtGv1Bq82RCA2Cunp1WJrefd33wkVcXjZbmpJX0
dQqoObwXlCOfS9lx5QjCn15W7NZ3XmO2X8GeTfenJhWkjslVplWivMRNAa6Ipc2Xe+BP+s5ZMxVn
TFdYtSf3bX91ztQ0fKD9d1wOc0eM9ouojBy/nUhXtvggTEQN9iHuNJasolWMZFRN+aBP6DV08iKH
qNxMz+dSuUpQrLsrXHR2B3A78TcVBwkpHsS6Ivx4/7qe/ZmEXDvYhfTUIgeIPztGyuMxOVnNfFPT
e99TXv2sdn+Q5XHpwLBeQXSj3OpHwbhbW2pjJzF0H4Lz8iqXOvuIBcsZcoeFcYrqCGB1lZ2l2w/4
CBxnFH5XEhRFRLnFS0JBALNT1kPSgkHh0eBTEiTdxwriOL6i2aKEWera2J4jVSY0o+K5gbcSA3LJ
pdegu5pW6m589UHJm7J1ZU14OtXmprf6WV2RtwafST4jE5Pq+/z3xGeX4ZsGgKiJpCEoKQH75icx
qXJoP51fCx2ssYNJU+9QzB1CfJThlojw1XL54QWwOySaGOdqgyq00tS5UXINovU+eo0OLc0xpSVx
Cl+JEBfBHwvRGhkrfK5UKwDoCYT0CZdgsIewIUylTFayIlt7/THJJ3xqU4sRRhXShuu3uIFIr2my
B8Sbui0aHiZt+3JsMKV/CqeA7gC5gBpz3h/mka15gSM5vdSV4qPEA7K+5fQsCZB2WTF0hJkbYLx+
WCOmNKlx/K3ybUgU2xajNY9nlq0jXXsb7Dv19kux7ZxP48oueeRygDP5vDihExeKOrnuVNjnSC16
+hD99117q+clouykpqyQdFJRNVN11cczKFCGYWT2gQ8EWHhQtxVIf9a983hMEXek2L2TIXKGzA7n
y1Tq/iIXu+WxA+dG0HiBCJrf8RCcKpbyT3s4Mi59jl5XX3enIYQCqIWnWb6IdmTcopE+ZZXADfq2
ZpZapwQPa5g9yb5/5t2ZZzDtViZ4IDWExFMHPsh/rWvXPI9HDpFyzB10RLFZINVsdLyxx8TOxwqR
pzo1mblpCcBdMPPdzHiSrxqTT6TYDlKAR1tOAGZpwPlVDpMMdKTiE0rlzX5T44ACQB5Vew/O4NKQ
1yhtvaQ4PtbfiNrRt0hEEfboTrLqXsJiNKkfhzaZrb4wwLwhO9wyCsNUYdimR5jZHQLuhqjg9ded
DA7rQhNW789rvHBUUyRaRCrgIub5YS/or1lbx6769YfsJmKB7DDq6NJni3akkpe7bwj0V9ewZx9a
VwylnwgmpoIT+rPaFc/WzAFrc5iHxyU33kXT53gtA7DrLl3VjrbWmtD9TXwxt/ToYLTunehNsnEf
10RJbJZDqGy2qZYjCqYyEU/CFb5qVpTeFZWrNZzs0mP/xzlK0hxcxHNLmY5Hgm0D92svHaEbAeqA
rlLc5N5ZMv3ZLOoxp+OlN1fLNoxpJzTYxUnQT8zou3eQ6OSP915NOfL0//XfcEdMy1Z2GYB/Dmsn
MOVTYipcqfY82177OgcxJTeo1woZOCaaVahNJnBfyWCBdW5P+Oqy0L5A9UmRdMmJlpkLDc/fpmMq
iRvVXOAo05811M6zpyklcCPHyerj5XkhfwPLABGAGxs3PHFMaEZwDP1YACSYXTggDKuhw2gBRCs7
QgtJscwzYLPe8f5fFwNrgRzmB49CHE5qgeUckSvI1GoBBU2RvLiN9hWYJIzN3iYkwBfqCmy9j8/e
WocLNvGmv9LiHQB48Jxpcia5LXAxf9eSnV5nj15DMISAcxv4joUBGdPGCdlxTJ2NXBaQVGld/TwS
KPa9P9LzTyrHUMyKPO7ftTfM6AuK5VABR/loDq4LRjxzcqy3Dp6myTJTR6EB4wFpZV/wMe8IKQ+P
8UEUmS0PdnqIsr+W8zjYPTZ45jxgInriRt5AKmn8SHxyRrKz9zApV0juqrjAPoprJrqtx4QAN29z
cjmVn7roTpbWNLwIMTbJiEKarBUxlea2hHCXut1sgjxy6TtVdXv8fdF+YnoBB9ts5dsgFzdjls6U
oA6Km+XYsG3A89ajEECk1gqzXl+VMhfR5w1vzWd9lGFmsVi3uIv6llu2i78Nr5TZqY/I0ILx15cq
ZbiU1mNYKwdkLnPcwaHUQjdYJHDSrWqPMR63nnYCbg3THAxKaozizLgTK+QjgnzJ242ZVXfvWS/K
CgMlDnQcxIo6oUo2WmYiWLTCW7stwG3UfPbtHi+oCsk9mKqXDuwZziGbA2gPNX5NIOLNvIor+ghW
vWp0xaaehZCNVsNY9I7iuQJOOcW0Ey4JBi15zfKtkkLHJJSIyAslWekUraGlPD8icx5GuLq2eQfO
SgLeXdUXPjII58cJaSkkdTgcQX6OzszgL/yguVrj6ymQITyXjsEnp9+F487q7mvlEkfaVwsNABRp
CiQXD38WVzxyuX9DafLkq7PArYBRUwIL/230bdxuKz00WfjNVTFHMLy8SCWUNhQ8811Hw7Bx3ID1
BLGAVTUZWg5tvA40m9UF4PWGIM+cQSOz7uc/Q/CT9H8TnKXBJczfgWvWHI/5PpKJh+fzm2mMlsvp
5JdMJ45EOHwtWMYIgdLwDnMuz0Sryxf7XbwyHQG/20xROS1R5ubV3xm/qCat7WRerrTQnJavt9BY
Rp6KwrvoIEco4154xQYL2Idj04mNQYMxdBW2hSXwtLJbp9gBiP7AQF/a7+hUGi0Px7Vl5SWJ+dE3
r/V7abJSD72mInoRQBsxxc8ItaqAO0Xdq2JZRjlq7Wf3DdQJkTcenMoeaWQxtqjvxWn3TnyXrYnU
xgoek7MgleZiddr1AKbuYLhz71OicZ6QP8HQyBRBZJ7idkBfL0Xlcg+fLBU/Pp0UFA6twUEaEi+t
dB0OAK9zU1Ik2/TfHbWk1R2mI/2jcNpPC1iWtXA9L6pt9mFFLywZIINbSSlpVmnh7hPeTuJ9eR9p
FOPMHMWrX8Ua1ZxYUVB4wGOoYV1wawfQKUwydVmyZ3W4QXXbzeUpUg+knE8RtIRmETeiP7jiSb0O
Ypa6hWv7GeyJBMhmV7d03pK4coMeUpSmUE6q7rQeCf+V3JHjcX388ngQNZ1NbQAlQzD1r318FPmB
krGQlsmNo10Oszj+drkpJr/OMb4OKjSJas1lfaaQ+dp34GwO8+sWnY6fUeRyHM08ESPqVmPI+hnd
JO9ddXCE0C96cdsfOJwKLM8YG9y3pMMvY9jfMcYKhM/obghycBiaZtRn+t7cLEQuHcjwJo95zOY+
YVarCI3GmpqhRS9yKsY15fYjcIOKhiZeMwEwyMOqUOdGItgmwngFwAS1mtrXq6HoH1bqVwG/uotQ
iTRKh8Yj9l862tnJ2T8hLi4GHqJ85cgOuVxWqiX7uAi5rJF3jZh73Cv2ngLH3XQGRz8lhQWtx3+O
aiKu2Ag/7eHUHDsmcqXMY2ZG1LLbaRfrOsqeciEUqmGjXdr25EyN3bcFPDjj1sP+Cm4Lx+6SOKCo
R3Mwcyb8vypfys1TaGQe1dBExhFx/iDfFw/jjHIMKzBCseKWj/6G+abrzV8w3cTZPRm5pi8cCB2n
0EwvWvXaqf/xbAvC0SiHg8dkHRwDDCrsVJioELhBOxwQD4+f4kVUMcc4a/7OKGw52v8gRzLKSlUu
jrDSj9JN2xLJGQUkkL5yguh/5j2yBuKmkipRSeqLg1lzEFuG8ut2CkUASKw9YzFT0yy6dEr4tkVK
i2SrmWd7H8A1dzA9Vc/2BnOhhf4jVxuP95tigE3pmXx4y7+eh5EgVMOxj/QIxBBkyTBDpRV4nRka
HVdLdRuSVFiPFues35rSuve/jP1BFhqHx+HsTb1F4l0Vue/K1BFyThYjce2KINSzazhGP0Xm/2e4
0B3K6DnNbTdMVgmYFd2chlc1/jp/Gn5YDtqs4L2gks1fQmgsFlRwdoNmPrvvbKyg/8Zb/5wSh9Ix
YkVCGuVqbkJn9Nw3uohOl7hnxrP1ZMT7o4UqzNnueIvx9LgVLo2pVsvd+MGTK6wJGMMF0bslH5j1
lpMhrSE2wO2uarkYUQ/HoaIQzq0s70zgKshFwDS/rnBWGXkDe09KYeewXKMYGmBC2lzzEd0x9qo2
kMePYCJAqhjXcjZEeGliMNTC2jRyj7BiaKg7VMAY0eKdPqQqH7ACbQWf4NyQHd3YVnmxoVZW0hEV
b4jnOSvh3+bMx+VbaeBLlx12AvBjo9Ff6FRcLk356HaXU0A6UxCgYnmlhBei2hRYak7CQOTFOVKW
xYEDtYMY6y9KrdNJ/WXF+JJsuYl03uHsiU+7fEa82S+ZWvfrt0j9I5Bj5OeX7EioaJs7NbKqedY7
d4NZ89xmcHBy7lCX/xJHI/yCaaCH0M05u+qK6UcBNJjWv6NBmiiAtYHFi32fJuXUj/pfr5+1Cngp
zyynMhNkU/UCzFCSxiJdVVScc0MKseCYXbHcsewuHhQtpaV1FJ5zp09gCHxWc4copTguY5S9XFP7
6846iImf+UCsXyob7alkEuZ1Zd3xYl+gCqBNAjcdsZ3s78TfgsoX1NEwu0Wcb+kWMuJjioxl9YEY
bt5NurJMRYyxMZcbZzsWqoYJn17MRSV8XijfKc1ICGVRlWNILNqzXdBoaBN9nnVkd7/mmOmB1nXA
MbiKGLTQQ1RXVy311/xyk3LQ6LOr5uq4yn+gXw8MmMamdlCPWRKE8R7e0C2OTB4X2B7XQkXJFOgO
zpvFldKvAHFmp0Oe7G7QRwwp6wdcEvaWydY7Mqs6dWHeJVn5B2mM6/8fdEAfc0OQHVxmixJzhUG1
ygPSzRM51mvqMLY6z+ugRCKGtuzkZonB5E7XLCEUrgXfJXVssAbuqxdOSqazAA+uDsL22CFoQMoS
z6g/mfVEpByYNp+pKqhOuRq1h4IBZX20oRYA+6y1UX1lLtIPMoxqqreXj9ffvvM9dhsHVcXFdpDY
VInxn7I7TyyopVlq+hUNkPPIqaAgr4Cu2HdPslyazzAB2Qb80Dk33As8cELiGHwAhnDWsAvjxzO0
G2fdfOGKcx0Qkex8uPIcsow/ouxISZZ/Qyi9HURGA36s65J2dbdLC5P2pY5irZ/zg1f+zwqYJ03H
ZLSQDJchyWqwcbYoSTV2EkWCoYfWL0f5IHKUbmKsVtwi18nUSsepvu4BfNHbNWm5xnxzBNUQ9BAq
HrEnOjQsMlJmciDXDUc5bRYZQB+UC9eaWvIUH0WeBDd5j9kjThHJmGDJ/bUyUQ+eKthR5GU1Mpqe
VRMzHQcMf1tsOtKjSPIVghZn8iOoLZE+5X8ztydV4Ybiy/8hIMUI8TsFgJnkT/z8eFV20eDT0u6B
hHPid+66xzurWrTB7wUxELPBrPm5XvhM7upDk3T9cZp5cox6W+wF/pcMIVmzFx7JEGYcYQZbvI2b
6YBzZS73kcZAQfS2jzDPRcdJmTm7oX5jO39unDJ4ZtVt7AJjTETsco9kNgl5w5TtNWfIjFRqSIs9
MLtxXWzhOApDS/Bti3F35l53atKQYUo5WtE9tF34z0pVCvqbpGaira24Qg1IK8izcvb2cM2kIsVI
An5fBnCXz8EY/KJKeMkt90KhOlfSh71nxPEFabiub+kiZfOFxBPl3/7ewZEZI58sRMikgnWukY+W
/bl8MYy3Pn408gAp5X1LlCc71A9OjKZrRGE1c2g1PzCKiV1UdFVpa5pIovFMOmRcpSqdf/BMutyE
PexBmaRxMy9/u1zO5GLh9dxlU1tNzexUajtQlXMjWoKXoOsIMciKpMdzGJHhn39L3+Ih4owc1Q1q
E1aCgGidhrNvLqlzXb+0mx6/W29J9hYTw0Id2bSH5GgILO9WKHydZSuGZPiIhmy/u9gu0MEDeFzZ
XDn/fhnuxVI+b9noBT9RrvDcMN70pPq96sxV81egTmvZLlAQi3pn+bfsjmzg7g9uqjqTCT3xg9Km
yssRJUkbekUIzDwib5NPmyNjBxgTBirn7yTn8LTxYm0wo77CNJMOLD906xYziyKX/fK90TsFj4iR
/xEUfB1fCv0QBLOtmSN45GYLMDbovROHEETkH8dOaBsrhJX+SBW4J2k7EsLR4znjF0blAWxE0J2Z
L88VPZlfclCultnMkn7WYaH0RMg6RIdDLjfDeWT78VNHZMAL0J+LKsHecB9J4lEpaqxOKv0glGIs
NNHq+18qaGpnBmHj/p9o5cOXK16aCyStHHCG8xIlqFcLduKyT5XrWrEOMU8J60R5aZbv/xeXDhT3
xjqzgFTgZ7/dDwXQYHA7HG80BdGWCa3oLLBVyTKFxaHSWqFRv3qoQ5pASiGBRlKN1DU+g0QFqz4K
xZa54kCX0/HSc6gue60S4QenoLltK//h5f/bGiav8VUSpgelzgY5Of9VAk23IEYKZwWKK3rTqjkq
5JeSiSTzPCdWNEG58b8v9/uZiamorE8u9oKegZc3LTt54LJvLIBPVs4iCiNRluoqVheIy4djjK0M
OWxJEfISf0/ekmj1oIwkRaDYSOYYH/uHytje9r6iEOsWDRtcRfm0Bw8DrMgO+O1kIqYPAyI1g/a2
hg3o0zeJL3+5iHXL02SNpFwQWT/zpgTSLK6YuDp5g3dQTE2IHxlqaoqpa3ML8hC7TRz4XeOeOkwW
mw7y3YdC3HHVrz6vN9sHPNZOQRRCUyU+GFfFimqJuxtAqWuf9BjIeoJqVvoetk1GUScuiPQUDy1c
xiYVG+wRiPL9NPqJWpbPvkZuyTu2WxWOCvoXyl3nT4L4WCRfbGGMxlzb2XfiTzJgcxPLEZwky2c7
hZHn3ul/4P+b1g54hP+7751NWuiJv9Bi7hCFpfR5B8Jn0qvAjsUhlCHpWryOWUnK/Dlz92IVxiKH
jJKbI69/zmlZ27tcygisemNbsLGqZM25lwc0/CjM/szvM1vjER2Jsxdi+ZdvFfaXitW8A3hdAd3p
NjlJH+Fmq6bp+UjiKRfK02icA1hl1O1bA6PEuSBKg46YTtSnTPiFZNDdwQQBFe2Ovx+QBsTxZt0C
fPSUZlt4ch9Jd80p8dnQpdlZhM1pZ+CjHSKrRBwkucv0OCkz2scOplPGHC04PpYV59FdYZ6Wj3vr
lPclQzxHB1icTbdfe8xI96nSXdeqT2wQbMO7ESKUCpWjYa3ZHMl3cHiIAlbaInST4nYbDLkwQM1Y
OqBYSRTBTm5UFqy/19VrZrtLd/Yk5zA1g+UsRJHTegSrv+k13jUdQLxQYJXMTy9ANyrRwDjOoE8n
audrupznkmmCK6tD/YtyEakWTNs3ro+Shxk8BCy657zNQV8ksfMfScrLosrzNSL0th8YRqR+0YtS
icmh9woyPvdX3hBRfvbVy6SydGh298jOTMNIs7JcUiGlCg5RxhVRCwVEQCdlImtHlCJQErLcBxm2
A538gpP3/Jp/M4OGP32724Msqu1pOnr1dFzJa9RmUYymFxxfMjgnvQHKII9M9jVCbBYOQE+qAaYP
MaweA+vGD37QKRspXw2OzOPrN8zL0vGRKnz2YqIEsSdrkV06KzQDIZng1VjNFTZpWJ11q6pOscp5
N84fx2L9rEnSWPVdz6G6poEnCnioyoTk7Xtt8+hel0OSnTeYDPAVjB2zn/yOK5sXwtGFiA6batH9
P8+nCNvmaRy3KP6jw7JKhPd8U0MO20dE2tfLY78uDW7bpi7rwMKYtTBuw2C43ssNsNzAeKHmINIZ
u93dmKTKc40V/Ea8lu2jEy7WN1s684LLqn9UUw8HsO71lvzvda0AlPZrkoYZtxpE9lWejgOUvGFC
2eo8TP6Q36RFS3Fms57XX2d3b3zm8cqXIfK8X40+YjzH+g6VX0zA60oy/OHzJIx6/a0Oc/sx/OTv
DKI0khNldUP8pRNl8jKkNdlhY5voS+tIK8fNiKPx5EMPGtAnDTc3dMVEe6PNelJZi21l/UosM4jW
CBfX57o1FqjJ5EOP0kXZiqPVA2fo40Zk5d+kuhWgIvMN3kNkUFIsx5h5xC7sMnuol5anCSjmamQW
73/7Tj+toh97AxS7QQ8wdFwQ87QMzyMP7uNBEynPpieJ1BzW0v4OjyNzrEJ/LYJ3bJb5tqaC2ZI3
Vvdxot9UMxVcL8jTu7TG15oI3OBlLTbQgo3PYdarve3eWfXbd52XZKlCcakVx1K0R2Us7fgqfGaG
/TTOPAJoMW+NGeMEZp+G/ci69jEhS5zAA4JeDJjaLEu6WHR2GaFliOr8weZJ3m0z4XOxTlSbmOI+
1tCZDdnqDUkf/YXZsNgBTAJ6263jAQs7BvL5mGL+92uA/zPAGNENOyzsHmT54a9s+yVumkGOcAjJ
KVw/nxbXhXn9kVjPX9l0db+stgC17T9wfxPjitACTFLLvlmhjpQ+gR58QjPD9LsBv7D3aj7WCfZZ
8rgviYyNrTwuP2shK5/RxXUb6Oxpo2exTEZmk6YLEkm3wXSJZolTDbubcWI/Z72DZEZJUmIsiHg7
wQaf8w2Zr2hUUUreOHckL98/OsW+a5OZS51xF8zCzKckQJpdNyxJXk8AcFvkvn6tDcamTcs6T43m
JY4Cli/iq1MyhqCGwFKzpxtK3VKVIkPa8oDPWnxBLfETXDYqJuf6v2jJ8h+z/4sPBZWCQqNCwfd3
rlZmBBhVEZeVyIbgSmRxZ28vV/n3TfEFUudmoNosi6BPNDRd/iaWVqBnfzymlAejOgYaXUO/NLrm
XK9UZzt5JF6Jf5LxK9XZx7MqGckSZ22+TG13tFM2CpWp8vwTVU1sR9E2mzfz9K4oFHbffaXXzUyw
ZUyPOojfTQqObVkc5WNoxycgeSZdRp4/ZTaaQ4q7CQyB1jwIU1BWNDYEiPoBfoJvySVpejPjgkzA
1R5/tcjnH2ahJOstFUWZDm9DYCWA1hQugo5D+lA5PyRHos8wShXjmr/VuqmbCl19HYFpEAWjdksu
JTGnUJ9LXVmikaSYmtElTjbw0/zgc081mat/WOUe+IfL0tlJPc7D79Vc7zFcOp/11LzLL6nHiEUP
Jihh9pZcq5QVP1HrFD8GTP4wMVaaBDwK3+syUjeI/2Lk1qsQnXGogn1orsSLY8Add7kwooEYjdwB
QEkFV7toamhMuQJ5bgPCwGzKQFYJP4jmtx3j5ExvLISWNLPdkyEk0W2gGo+uRAfePm3cyj6g55LB
6Uq9YaUFvtVB5UwRgunc9ezbSTdRl1M14HqOzr7JwL7b2wlAotTwNLIObkfLTNUDK0w178IP8E9G
011lVBI4kELA8eQpceEpPayMQoLYkLd2d4h0vbl07XU/vDFQrWXzxcp8CL9/sBFDEMizt4L7HVHE
nXzfwkF5q5SKQl7lNSx3fUrrpQ8kOj4yDpHi6PMDDnYgdgsbafWRdEeayVd410ze9dVd8dllPSdd
xog0HTDgy+keOArrxWfjTqfcbHAKuvcOa7qCzqa5zjfiWjXugXg4Q1Qtl6QJFx3QRpK9Kjac4vPd
OT5Q68c4wSOO1j9Pc1hD81MRfludHEoKzlY4/SsXTmNLhJsu3jQ3ewCOXd5JiBUURJfer76Agwfx
GL2KyWocyEqYB4KgIN5/76Yefgy5GDOCmsEQDWuqJLMwUCu2s7hUdkzU8PS0PhKh5kqvUABkhv2Q
IJOy+TcedtBcdDuAWepF2UkPm6HXv7B07eenCy3ZD4Zsb6ZAp1st1RTmRcaFxrwHPla3BKVGOsK9
WqGT5r7tdYiPlibHVxUC/HEHJyOK5W1QgFIQuIwdM9CS+iwEMf4IoFrSAYVwvtGvxLqLZ+c0N4ZO
WdXjWxorx7MByGipFgaAIAoR9tNfFRot0NyC+P+U8tUaPyoC+qgERXkBX60QbeOoObemkIjRz2jg
Bz9/PdEn0YCxgxyJ4pSUTrL5a26j+t9wAqFuCS4mrjGNFCULlx+UbAuu9SMhXe9yhLHwszjxbCXn
HrPHKM5GWGYVWcSmi2FktzKO/mNfZnWfjv93SA4mxTgH7RAdizLnVrfuo/UwYwaxcWEM6DRcrwCK
kq/4E0ztSEG7E0yLKQUAbSOQhXXDgMU59ybElXF3kPlkYa7EonkJDtShX82LjM21JEVkidKMVk8L
FSnWuCxzHn6OmljWVf4JLNw+hraQt9zAYKHMgaGWQ1lW5F5/mRUE61o7S+YJRPxV0EnR0CLMO71k
xrZSI9nRTvhJS9m37ZSzhWFATZcshAfsIviVNpstFjr9dbpWoSCdITWVqVNp3FM/mZRpmyHxyjWF
mXgf/c7HRNTGE03VktNr5vVTy6jbu2UyA5uT0z+EsLgTgU2+/oSigfuDjlfBR/QwNE9p8x4zzl/A
mxybLgFqcmtXVdP74a5x1kAAa35mGZB1TNPCTtuHLhoNg3iAwqdxGd4ltIu80TTqTThbRVR9LywW
9WbONNN5Ri3lDMBFw1+679jJshND1FUmZUFVdoav2A6j2/xHagJmgSRx8PNpijgrWegLqiR6B8LO
ZFULRztULa5wDf0UFYi7APckzUT3cIS+tvE5WjP6w0j180D+knnkXDfhVIZtCQ30QMXAlZFz/uZ1
AtRNvkEof72lIDM0oILmfdx3hncw++x3c3FUg92nK2BCr4PyMsLvE3guly29x1zibEMN5i+sqL17
joQKJWWCNccMzoItxZA6Z5LrkU57Na7Wcqy2n9md7h0gEYxtOW8ZCnujxzUHD8hl/ShNY0e7W5CI
WcWhfLVR7zjXJkDGGrMB+izD0v/9WiX/iE3rJy9bzHYP3UVyqRCADXms0C4sU6fyOlBScJPSV7lC
psC169RdiltfgqRSU7RBOuLK5CBAiajdYGElF8P18Xj+6Z9e8T9srs+LfnxlZ4ctDIhwc/a+0rbU
EoCnGu6F6PaMcmu7Eh0cte3DrywXxtQFF6FikvkiyWuPKZDAehombcUl2FNeKAlaT2lIN9uaXDUO
gIwnql/OhnJx+nGwPyOZpoPDasuPoAilL1I2qD44aPWjWEfpBj1iFvl+iZlTC2fQzOVCkU759gri
5VlykWUtz+vwFDMof5vKDYGKxs3LGJFWNHUQgiuIAsLtDR0aQ1bIBr2JEo/DJL/dBkQMVYz35Wcq
C1zKJlL3boKp3EsdoF7m7XzC6qNQvfFXHXVduljRngp9qEeh3Ye8OzXewHcf1r2w2HYtEaRxCz9p
Rikp2TKCw8bUPEEgSQf+mUkxp189tfAPXXilTdhdh0n+WF0Pi71owMTUPvFXN8BSvP79Xfob/eAX
YCXnCOplY1RC1K1gkID9O6aKEp0kbjxZFuikCBjldWD9jDfuCwfHsEz93DQATRka5wgkk73yUuQd
rfg1iNXo5NlbqAzXxEkPqs2Gnh9O/OGFj0D3OEHwPPamfFXjpa3ZVknDqc4WQsIPcmhTiIwHamb5
yN/DyJs2jiHE3Eu6MqyWyvHM960hZuBnMiJ0YvF0eejY9LhTWLypOiyiVHceq8iVrh+BhHi/UReT
4oziYJbf+K0aelGH8Qc3B3QPdnO5ZpqIQ6aUlGg1IRwnoFLhT45CGWkEb1R4/r+jY6RR3FwQZKyQ
2sfNKx+mfy5cq8fr1trnhJUSBZfNRi99WvWSCdHgtOdc/aXERzNI8o0reeM5vtxKrQm0Usr6VVjz
qmGmup7F2k2hiPc2SD/z1fl02pO6TF/aujELTpWQkDl+tKq6CJbc8T/8VzwnEb/HZlb2A3midlUI
tP/yc2T+xODqqSMfiJGtA8hvDWExACcRysSzY+jC5ph0VVq9yTyfQ4ws+TvWeI/mCXcBdmu+k6WT
a8ZSQ187YejsyQlu+9vRY3r1FAXpq2Wb2DtG/vEFi5HpmPgJloTODdoxYSoj5HWeeNYj0wJlJXIy
huZt7owL0ydxUBXECwVfSARdFjqXE/mujCWH6EraAVnYZFRLKG6/kjQIpE9a1+H2M8/GucK8jGXs
z9qxC3PttpAH4BwyMrhaV62n4MVGQUFBH6GuH0uAWFpTUyd2xv81pa7j8KJx1Fcp9uZSiBdduJlp
kcU8yO3nTNtNzqOsvaTjIugzLJojOParix6SCmPYkqwP8mz+YjNcIRcBHCpNOcMAq0RLfxJyZ7K1
+cq3Ycd6noDaTu2k3e5t0Csp0+vNBl0428uSvwvq/Fj921OM1HOOp5qEx378fgxRzWlFYiU9GBct
fLxlXkGvyhASwgEo3mPhYE+jmOzxHJtWifIlZVCyfd0vm9wGj/cKpW22cq5YUZ9ANxmkRyp1+Jhu
bZo9SXV8sYUwMdm3bSbhNz69ERDtMJ3fIrfU0Re1MpYi4+gUn02Czb6pKtm2P66UbDwZQkQRzoGY
Cm9L7qeYWReU8ON0Pxc/BC2MV6yeD93scEqRb+UzunhdSJbQNlFfYn+koktUobs4iWhr9tzC0RlZ
sJEqES1kmd43roTHksyZxE2a4hpw+DjmzI5bRhWUqwPd0fd7i2rZtm6Q5YfdW4sPdM75oI7HuVT+
wLaHskPEqYLVIH+iBQQ7osW3Ah8FZfhFRGUMyCSEyys6nAmIRljRbupk2uTax4sFKX49HwWzwGZZ
h2ANwB1V992X5XO+auPGkXIcQNEqBBJ6rPs7SF0LhELb1GLelIbx8k/9CSl6SEOdC0fnTZyvAwX5
ynCRhzmqSlhJVD2M+rjt43AibIzzxW284vhLiI9NgJTW4XQYW9yMJQwawxd3Y91whnqcAngYw9lE
Af64bCt4QqqGbIPyqkQwUFO27C2xFT6mHk/8uImvt1/DyOHlCSQW30rHulQ1IUvyaEgDr9wBKDkB
/g0B06tWOJb6SFGrSP2tjL5OvXLRhtOpKt6y5mf1OG4Opdi/V6up7scpJOz4d9GJQxXjmGCpkHZa
EapZL/6t3GDhhTYnftJfphSRLEI81cAezQ68lbdHbVIyFIhUssUWSHe/+Ao749zxaWUhD9oEYvPn
37temKLj6VTNPgldOpR3u2WMBalNYT3aAV+82BKE2NZnWYRkb6QtZwNLpF9VcU9/sw0XUyVAhJYD
0e80ykhU2XCFw4V5zkIlgls7gDHl/+hopoiRpBznXD5CCyoMAre5Dz2gz6J+lUC4rj3JA8g8KAPB
ghT08m6M/Mc8nCjRxLySo7syHZy1PQizB4WXefkQ3J7mUJWknLOzRCjDroaryMgItNI2k+94BvXQ
EVimNfyvXnQUfNom166ifJPnsxhl+MfB3G7PfLkJPNhV8+KqzfDh19tWWnhGKrSXDx957UYDyV05
8OT1tSyseCcWR/hLTIyo6soD7x5DyihBcytnkR2Cda0jb7gZiaVOmY8G3ksc2prob5tlvie8ZZHv
j3kvCg6Xj1OkdygjQEw4pOyJbKh7bIphTJ0esEiw6sjouDuYRHSXTTecWYZDar4ADEaS3eJW9DMw
JZRgl9yAvAGzg3g5UrtDVoazt6q5vh9DQ8Jb51X/xJTO9fEx4C9X1sJrA02dpfVIizz9AjVgWPvJ
aryc16XV7ZCiMA0pIGTOI8C7ZQDVPdb/hIkLRj/JU0deBEhdJCkIcS3XvFqA3h4nA3a7b5nMOh1a
Kro049g3b/nxb1TpBXHHG8lf1/5eFvNtuJ3sJT9aWfDwBYuXKX33i047NqKq4mo49hkeUSB3ZEbS
Pe7o1NSpnRlAy/XnOGR/xj51lsgMHzDqlmF50wQtxF92oVwZB2E6ctIKEJVIuOxDiSBurnVKgC1X
2u+KZIWY63040E3Gff/wDTLA051Td1h0IsypH8dZNCF9lN8Sg+HfIMjuRfJR63Q4dNak22nOrcI1
XPl2R6F2jzscDGfXIBkskNUUJTPtKYAoEnuBG8Hfm57AWX+16SE87VEw57M8aL5+EzNS4DZd/rOy
Q37+LbYF34sM7INmViybC9tsn9IPkUCBTzK+L1c+SQ7SiEA3nWPAUYTsEOWFADkf78/zjMmQBlFR
AT3mlLIShK7ZbsfrNmq1RV7vwvlj848JmjoMNDhee9sI9y+mZb+iBmmBRTMnDbYoKDyu/bSO+gMS
aKc/pa7y+StgKmn2FKaX1uuEY1PyNjq7G7Yv4cOqnzge3TeOUawnS8RNunMGCR8ZPlKi8CnVljK8
gvikDnWqwwq9cPHNUt29gS7c2aio/TuridqJMZONrPGPrp1ADgABj4ekGgnEKckETSKCcrKgimUQ
taN+UH0y2hQV8l6undCGpYqUjsm5DydLpoWWcnfHt8PIJliYgnSghZ2WLWUdj2mLdpqo/DUp8xIs
ZTdx6NGOhUXNAyGRBrOXIoXzMwwnlz3Z2Ho+EMmMSOOgxSzMenolI6QbXsaIJWqOyQzgOWDVRoAs
GnmKTrMUKoxVs06fs2v9kEkihUurxIfi036NMp2b3Gz6rOBORwlqoMwvibTnThr1vqStS++DMwTd
wioCXb2u3tx/zefApxG4Fi8FVJOFiZ14NYB1ok6WATMJD8mbbpG9wSYjEO5Ookbi94+VrhNP+VsK
tufJHlspkKpOnJdEAyjfxviyLGvV27AYQcPXRFaLzWvYYrUOMDGuPHGR9AAtM8v3YKxgyAmLlgU2
R87lTVjvpIjuJd25Jz4C8JTAgYrgDpH7gAsWxspmp+nhH2yFv2KPWU7AxW/090YAn+NZhrth5QfF
mc47PpenzE79gHzFbmkLwuuitCYL0vz6l+edX1DOgL/wQxQQkOErWGFfm5s6CVosdImajF9eUkYR
+LIXZvUu2DBPIdiI46Ft3/MiPZK0De6RuoOBZQo6lCMaPsx8Akv/MluJOS+RAdpWBg6dtpIwpMpg
Ms0oUKh85q9/MW8rOT66qSRbtMIMmOjGA0lllXwixxJGWRPacfALuMjU1Sc73zajm4n6MUZigRCI
ct+HA1TpBbETgL7TVFTBsSj8w5ZKqyHvKLh9vGexYUeuo9N3YywCj2JFJmThE5qieMQolbuhVJIc
WzfMAnkm5UOLBx8UT7CnMXvnbacyZTKJLhszuKHlzcgGqe7JRPQVxTpcxOU0JeFqkwYBGM13PLhL
r2neCsx9xFZ59KuXxcwiMumc03vyrI0IYIXGyIGt/PaDTFw4v84Bayf+0FhC0YKD2PlCHRW+mIwY
NrLqxIjBxpmDq3ZMZoIIPI5xc+9oyxMeXt5SCkqQsqrGAON5Zi1CJOeTYiqfmA9ATwbSCBKccqU0
E0fcpYwm9bEZwxVCNjIGncEOfAUWrryQbsI0aOpyftNyP3RyzCCTlqHLin3c/ZNu4EqZ7dASgwTG
UfXdGu4EnKgeTOooGohJxWdutw6vgIo12v6MmRSCOBv/hxg7rHYl4dRFWqdYMOkfvxotwY1Ri95s
L2WBbBwCa+hC2cT0RvTuEFkv5G0iSiWhMl2YI1rJvBJWJKqwBMcDtp2vPK3fBfVCGmX++tkD9av+
N8MxCd2q/oMkph/LlNt0l2jT7Iwk1uRmtDn8+HmSdQeFuka6G5DGMba5W/B4t4D0lq0quJgindNm
IUnKvwN9t5AAAn+NrspiLK9DpKk/z18jlLiLMZIsxXKxsiagpqIzMCRWTLqj4JA4sKpSrRF/gPyI
cnhGNrvkam8jyjhe6g707LAxyozkB2FRCtPoW2G5bdzcFn+pmkCYXtudo4C4UFggKscCSEl9W8wi
S51QZKU3Vs+1m7LCIeM8fS5jmslK6bsSf6XqHGwSkkza4xkKPLkGJotP6kN2Tylz0iwsagUv+Cfy
y7QthSIjljF8BCulkyGySnYWdOIJvh11m0CTSG1hS6HTIhSsesj0HjyM/y+RD5fqqlzqkE2DgXGz
oWrMrhkfBZ+DXkHNyfZ92NTAooI+Wj0bn1w40y1RIdUNFe5dwRnM6PCa5TfHSLqxGZcR08aEn6U6
anfhDS0i9XIDjLLjMHWqBC6XQmcIdbMAxH19Soo6AA/QwUhVQ9p6I/o6ygiArhDANqCRzzQHscN4
mx63PZldoLM6PkG0vaC3VwqBGNZ3zhKY1KjKCJ7lEizI7XF67oqhvTT3PwuttgBlOcsmuFAlEKbU
7NRBarwiP5czSWQiAX2NPgXaVrNLLBIvw9L2qTHarN64UjO92y4HpZKk2+dLA27mQ170IWYeMEVI
E79f0AyXvVI68pfPHLGO3IBNoO0VJESQr5tbsfrODkCRe93W0Zkr9VjDceMfJsb94Ze3BHz0ghMS
5eTQD3TAwRsJ1aLYoQOcXpkjIMN7JaORRc67Mx1lg2isON57dP9W/O5EDLymmuE5ZZO1kcZ44Ql9
0tMe9ng6wEr4LTzqDnY0DeT7KdsD6i1cQOApgGzGEmW0aBQOVSuYRDnrvCsxkhZhWMCFfZ1nZfEr
MRujrh4rggVivzjDwGs8lTIRtynYWKoJ/4g/Zz+56cJYZiF02piOvIWcPv7y7wRrJdV8WpoIpE+S
rYDPVROYfbFPwUmSh97LSaYYtuYI4wvIRy51xveM3zhJK8vzi5KSQYlfgXUydntsi0Q0UIXoyk0Y
vYx5ZfBMnKlWVXEmlXS6aa0pgFa+UvaBfAaXF2T5W7eUy2V/kTSfKFcFy7ERldtk28Qd30JJhi52
vyRVntdvfI1CevHA3YE7liHoblY9D8OzrwoX9sbsU7NCP8Hi4a6h6fehS6mlLCwGKj2lBW/7+K8B
yZFU914S1AE78a5hchXijfN4h6D5T5vePJu+v45YMI/iBigjzprD8wcqciI596xqiBHyOw2jNp8C
JdunLjnx+VdV3CkBZLYpsjErnT29EOMaYmJWUsbupDe2pgtRPwzij4SjuyqBgr0fMxv/4fcKKcZu
Q1kPs6EpXogtJrTN1rFb+6XYn2AOFb0rld7YSBTO4sd7UPcMU/Ot2jD3zMUJ8hQ/nMjdnTzpVihJ
IMdjvEztzSC2T75WdClJPM1bgtrwYpDiDhmoEs8LxyyXrKUae8RacOncybZAKyKe1BqW8i//xBNg
As7KjwgrAmw4/f76FLZuXZ34I/1/PDnbjonoj5gukwbXcUVIWR/B27ky59O0TvgCZkAZUeO2hd3B
UKsWYcrZHYr8ebOHeRzh8ggdKbBcpXvl+UggRVlIpAuWbpgTrmFf5tvYRYZCDI7n+5wVWIMCveHt
Sk+dn9X47z/LkOjImnBhkR83MkJRANfd0MqSCei8aqDvv7GON5h9Y6734L3Tzv74Aab2ufmBOjGE
AZMS2d6zXdvxxzDv5hX02pVfPNUgVSa0b4qe8gzj6OZxa6ubnH5yty+XVA1UuVyCHddMTT6EWnBk
TNhinuX3j7MrnUDOLCW02gpCtCugUI79oUJrZ6p60UryEpCKpSxplUHVmojLW9blviJmNtniL/fh
ZeBprB28GnKASYWXVYg5CWjgiTYBmY/cEZ37gwgEGcDJNZPTISp1YxE8O/DBnnbS1yGHH3RBrJbS
7vWANUEchuKyI5OyGCAhIDrzAB3EOSHqmXxXGiy9QZ1m644ZnIoZdTxjfk54TEYLxktE0WgnS7gy
uXbpwgboRfVZDEaON0iEFJ9z47Af3uzjw8a19+SeMk0l8XN60wti0EJ1CeVp5pZgNW7ODMYKe9Ek
eCUe12SOYaVAVXZRlamJQJc2SzY2V9QHR6c+/ktnCg01djndruGgMC3b+H/gw5pPlZVJGJ4C4eTT
eHde93v7GQsV0NKu3jM6zpyYYQdfpsWy8vaPUdMBM3xmLbfKgT3JyqJPrtBM9U5Hnv424aQjq2B6
goYJZCSauaUo58ysAOzflUxpzXpGM4HqyiJDFomruweWOyseyWHQomRFDfsiVashTM7kjarFbKHa
nh6s+qvp+ZacwOxnMkwqpLB+Gmf0VOKSmtpvH0rIhn4AAYkuYt6p3mSDrMwVCB5jQIdT8D+eJpNb
xSuYHiuTwXI1lRDKIIs0yPUwqLwAOE0ikvNcryjlm3bQz8NQ5c/cLkij/2Rpu62rb4ViPXTu+wfn
AMSQymCibLa/jwu44/FREYyK30NL/coKb5qrFfhjorytomWY3/3i8iUHSh+NGh1N/BjxBbmb1AEJ
WwTTjWvyD391B87OKh+qFsoZs4Snvy3IqLIg+gKHWfdCC/43n/U33MxgR31ECUjSOMNqCbgTe5fg
lqCPew+DFGzVgGpq96hRGOOtXnNLD79Rm76UuLalYuBDkTTKE0nNedYWHjLCKl4a8R4hmGKZL19M
nsWPWUh7Z2irzQ1vTPE3X7B7E0JOyZychEjORhYJW2LiNzWuIveO46YbuKwm3euENk7i+sCgu6kj
2HsosuGpYzhFHAyEC+6n/9jRSo6kZMMVIBj23tvd1k8SMCCizhT60NVYvd5raML6+g5CEMsdU2IN
ae4fhvX7SemRSYLmp1N6oidLVWSIuy83IJ+rJAea58grCACpyeBCnSCSVaA1/VbkR27H1Nads7PW
Er7pdC5jlKA45ZEDmWm6M7nDoWwaOHZ3dgFm1XhgdoL8xONV30BH8cek2x75n99oeHdf1Xo9isFg
Mv5RSsE7tdsF62+Befz8vrcooGdWVssbeXuaubO3CAivaIjCSrzkecDerRZYjWr1bTOP6j20fbDh
gobPPgPEomeDyhnYqOOsYx9kNsnA1vt0+65taVC6lyqtSzCTPlsQsNmFJBKTJwPO+S+Zs+KlQfrH
9FY7gwN71lONy3Ya/51Fb9eMcUMqM5hlwhqvEVPv3WROYyuh/kfXDNfrsTuP8bLgaLilfxjnsooX
14HvaIjk3F98GjBQgU+nv66MT5yxbs9Z7boUAJND75R2AJCzsKPpxCEKKOhQxXEl7PNMKQDskyKw
XKGelhI1gG0KBBxL/5SAyH+ojLZj3QLsmsdeUusbu9FcNxOxkrwyQ9bYS7A/+u5sUZc8dZqUz/hf
XtIYwNnFrd4gYzk6j3eLCSLNATbn4kOmyHpYosA3rq+jr1DGXXuNRoMctSCcgB3rgV07LiZojaVI
kO5IBcVsK1Y7D0Wo92xTijn7xYyDscnu3BT5jhEOs1uyJkjHbpWyl2a8BaBPaEsOyN2Gbw72S4DJ
0B8egc4RmH13YhANSw4RKa0F74YMpYs1Dhdp4Etlo0qwWPGmatdsVjGj3WzpHeebyM2X11j/iwLM
IHU5/2+LK24XZuqlwT+4l2MnHOgq2QYxb/ZoeTNnhVMTJlzgoqglnWJaA6VzNjMcw9hvomkIzB0X
HFv4jYS0UlpXxpCPna1aI4HI5GboE3pETbU4xO5u1tro6y2ozShsaIEEnT/ofK+ZRphY+YEfd83I
8jfCVcs9JYWoOr9ukyTVrPv87ZWr/ix5lW1B+8Z3ZU8iB+OqAgQ4YLDvNpRW8QJo+hCjLfqpXGCx
2xKycW4Fj84NNPDHzF/6LgiR+pgGxB5qiedQ3tsbc7MHt9N5SZaM6+Ez1RY3+Drf3sKqEVjDGHuX
EvdKnQoG/BM0tQB1Iy/XLu4Ur7Hd73+3INSXD4xZ9aUX61dLgHSyDM35YzgvvS203nw8kaxRgtKQ
H49qdAqi3YRNV6jcU+iZOz0O/g+vuyGz8AmHruyoCR8xjCO39R5g8J3r5kUd9d4YgtKhXCyr07yI
fLaHjoOuZVbvhGqMpXUDFcjAhC3LLiS54nXm0/9YgGnhWZH54UVx+sJ0O2MoCXgPDpAlwwNwtart
9dJKGz0JRp1nNEz8uQO2gl9L2ld3zZlQQdOfTZS+KbuFLgD7vl7rCqPB/NSthMdgfBeUXu/Zm5Nq
ZfDRU6dmJNDoMaQTo4vHl2PvFhX9OUXDoxZygHqFM8mOyaW7g7qTYbguCq7toInjwN36tN0UQ/3p
t9XR0xrowA1d2E3kBpUG2dsfKQurrqEZRNhHRN8ANlbury6y7NdVxvTFU/0OJ3eqWUqWBZWfLG7S
4p7QY6wePmQcUHY5beDzxZPk9o4uwlm2VhLFnKgz8WfufyKPX5gFu10aSsZSVtDsHV70GGDikjrk
hHrF5BUXwDs5Kk/PeSensu+aB6tPR+zGYWtY7wHbB/KWVdSv/w2NFeiLizwZzekeohRkj9JXpvT6
ITdsO/AMFYUxIi2cR4/5iM9oP/suJFCS0r7KyVbhq7ojKP4Ln9/YEy1xN7tKSACBeR1JQJ7KgAyA
HOBGv51G4wINhHWY7AuViNw/aCFX3sJ3EgGUhXgxu2Bfd3yTbYsp2hf4hszeBYPEFAWIBzaOU0SW
9ZPHIHexsSVUO0Sd0mMCoY6GE2ZZ2tMT7o8HYR1y15MRGtXivP3LgYcD/kpJunNyVHMCNZhBa3Zv
q/HVwU08iwqVEqR2RnZOq6pTW6RdmYWFTuICTJWZLYg83/3TUkHmjDznpjAVviic4MzmVhgd7BHh
Rtmom/NWDEIQXu//ElnuIyBPqkX8pSmlsG0UC5uWo2dyJvtzxao7kVbpntiI/g8T4zUeeY5zaJkX
x+b9mZ3ARtEwz/ADT17aGM0dLs6Dvx8sC8nfHn9QqQp0s1f/UrMsDxf5i31E1/LtpxW+WwjiEC9y
r0mOfwpiMMbzynV/zH0CwhkNnj4TDkZ0w7gyFbVj5B7JfoCA+sjHvQlDeet2c0zp6MZSy5ZiyTh2
QDUAXDHSHoqQpAhN+fApKVRiIoy1u6v9IXvbKyEwstWkuTEU0WbSViVUe2X4KzJgA1NxWOCpOLB3
v2kZLNPCtLgYdQ5b34v2gPy3EO7TTSFcLMyl/JoBbiy4bMozfMRc+R3ZD7s9DdWf2WERZZQik/iJ
SJaWVR9DrfM410ZECbGsH2WBurRPCRMn5BdttVETQmF9wFr6k+qOm0UZVIE8x1+wqbQpK71DOIM8
oF8ibu9Mk62xyolfrwc/WaMQxxjHU9vUNVVQXGsO360vwRSbtDvodEi3yrMfhLhIIVosvc/OCiGR
yvu5ga1enOgEEGlaV1g/l7wo8lsLoToKb9iCkpsVGVHca0DW5NJM4eWVJxnCCMvYtjJU2tpAe69+
kWegUFhFe0D/7XflvKZCzcbgORQFDeX6NyeWqZaZcA3f2SDyN1yyR+bjDmGgba0Znyr9zvSZedSP
9xvIexb2bIzk9R7Jq0WWMMevFR/wJGw/usdet1aH56Oqx8ZBvxEG/Pf2JKs4x460wiz0Lkc7OWEM
1ObUS+HS6ocNMfBPPUGj16CvPeT0/O+bkK8Cf98lRnDecPdOsYyqeNbouaqgJ4bEp0NyoDHUVF9d
yf6vQuS8oU3D0zJUFeL6Cn4VTvuaquUSioaB6F/1utt3wMiHJhwdjS/FkQGtXbFLIJDAc8MMKPp9
izvNtRPKkyXm0fmSErMJdzw8xNdrd8lx0BopYifyeOdXWiW2i5pRL+FISEs+UsVatZD9akl/fDWn
esb2SQmyicnIUYsFwZrJmbLUY8JLBZC5mdLU5J80+Wd25yqEjv2RVplojwPJmdYoSfeeh0sNRmZV
ffAaeM7clIRI6O3ZfLxPG45cZiFtrQgVwEMttfI5wxvak9KF50f6WlvZd1PYxyBCT//xnzP9bCwK
vO9oI1OM7wZI6or9QXlC9Ts+wrAVNw85l4VeQnl4/w3cXN13uMyDqf1IgLnWeZm7LO7hsWSIJclV
reL8ZSowLVWGqT7/lmhDjCouYrWcEc96pRO6UQMvMNHLxG0XYCUymnmnYR+N2epRwYzvAIcdUBVs
mLQWQZ+aUnO+s8zFlv88FJR3BlUARk/Ke/m+7Z/du2RAwWDQnISJLAXibJcwNp9AyslUlvoWcU/9
jkNe+uv4S8tdM2vrG9euTECUWzKt4biYQptuJr3KD2Ahwr5TzbIv0rq96e29JFN4/bbEqKAI8HlH
qgFkMxvIa+OOs3koqVbthuBsjVQqgZnAouK7ZWHGui9TP+q0tvtMtGfsjoIeOlbjEKSPbCsgwSMW
/yuWuRYZciePvxmQCtMgGGYLVnP6JGfYlTTcdRTOMIg3vgMQSZGhBYM/zG3Kmy6H6U+jiiscHpZ4
1NQ2Ynjvu8mheRvQSptMq3JgKRu+IBuerILGIaVMsLrfCTgLa0i4W1jFzZQ5I9lkMh8X0o6isK4n
lm8xKo1TbQ6GSBZYJ2+F4IeDtQ0ak+ccgfHXNAqkLl36OEctDLca2TXk00wLHZiZ27SXFBDHNmP/
UNiJJp5DcEsRN6oiMo61PDhWecOsxSAiQZ0KZn8HRe6iWM030QXBgNJ4PuPtBqDQhuOLPZLSkBLC
M81FrxklaoyKfpRlEyhtPvUFAjRMxvKEkywIG55cQ31D9WGOObakSueFA0XYwzngOrXfZQNoQslZ
1QlXOD+dZMmjB08qzY9Lv9rmmF0ypP/7zECVnOKZJYy6y9IQ9HIqHXN35JBJ8NeP/Rf/PYM/WfjA
5X9aok2QjlLk4U5RN8+qyID3CC9i/fL4o4oqyy3zK25hTgEbFR7slBIBMMDN1C56MJNGVchK7XkT
bQTYNqkL0xTruBx0ALykDOXZxepL0Vb0aklrBsb/jTnndchDvl77fwneDd6eSPMpOITdsPTbpxIE
29NxwaNHIHN7sHbyzc4eY8aNzkHwTQUBJpiwU6R5iyzpddONyM11mzw+7SyPAHdrbMTsMLAOI1SY
qRwYYALTnIFh/Z/83K8mHt21pmvVHuO8hP/wLssFYzBeLlu7WRKiY7cllThD7apOCWQ06scxUfY5
/Obv+gFZveLnzHfG+BCXmU0ZUHr+i5wsHbnjPrX4VUQy44fowLV+c1CDZ6dmGP69dEjYjDG2MRQZ
Qf7GDnU695P0I1XqOmEvMcqU/ncXnXSSmRAFslXUmhl/8WcspMK5Nig1CvQHrEQODsWZWM7fqVX0
fn0PGAbq1g8cVJhzIQqwDNPSPcFuFjtz+3f0cp2YPM3jUK0zABG9sZGsy2wR4nVw+q3OKqC2Zlim
iCJXoatk7PTE4e1jMqWZosVpSLiASUmXN70qbXbCQwRI5sBoXFlPJrok0BOxC15bUH55D4nJYxH0
4ZcG658b6kqvwUccnvETp0T4mMNaZHATNGYXZRFdeAqqTIW0xOSvI7wNqYaJuvNBESkjG6wS6VE3
Nvg7qAEIlcr8m4LmPuolaK741vmwGTE5em7QU2WZIRUTY9IzRF4f93YWKfRuSSbhQbS6en3UOeKO
875P+w/LDH6IUgjFRvuTX/pvTLi3GtVewgIV0TCoV7xizwSkr393ISQznisbmtg8Cgw+L7Lz67O+
uViyuk7pExUJ0Dg+WCbdtoiXxnuw6k1qC3d+9daWTio9SlwyTcgxxZu0WffAx9M5hKv3QMAlY3+I
aQDwe+k21LR+2X/TkmMDXbqGXVQMaGBq3i8aTa5G8wA1p35ZkE566Iu2qTa3rT9eE6mbiYClmprL
7KULV0S+vhu4osXyIk/+lZNOJ+QTuQrgWk6pUqqJrHWbZKuG/NQq21Zw//JYFP8/sXI2aDWD75Rw
3+wAW6osXnrIIV9B4cnUCMBE8RJTM3wDmRoZppqe01fZmc8jNR+qQ5z6jm7Ed0Xvw5uW7ClZDDqc
l2r7dmXS/NVGJrtLp3IZP+HfD24GXpx+JUfGDq2YHsPMsxzvFxk8XXkp2/jLCFbpp5yBCElhG/9J
EjycbR7Yrd5zZgET2I4RV9Qp20HZKsgbCH7HQRLzocuv3x5RkdngbsSus0w3HFJ8dPYI1BWaGJxX
LgiwnudCNeNLMtSbpgcl6Qu15RYPGZgYmaZ5YF9kdxzqQBY5AjcTaJHz083V9NgXWEbWlHmmGcIF
V+TTtPgCQfquae42gtAmfm3kq0N9TNQB8Bd/9IrDnfHgvOTVMios4revis15kSUOExb1y2+6KstB
5Pahi41Ij1hJntfFhDt5aPuYEQlXo741oEbRpbAEyTk1pAsBZzw9sAz22+caEpM3corXTr66dZ9D
IHr6Pfvk9jdFTl5Y8bwTfWrfgvvTgAWpud3Kct5mKnA3UJ99QApBEVRL9HWv2/uaNGh234PY+/Si
jJUvTjAl7wxuZCnDbanrdsHGLCiKKVtO7PYb0CjR3KYByIKGy3hxuQFzAhI5yKTiW4uatyzqihmx
dINNUDcTnSgBu+CBQiYYJHrxA09slElBU+rREnAnPWNHgun72/CwPp6W6dKqArRSivtyeudwgRxp
lgP26K83P4bwrDsF6BHKv5CSGJAE3gXViIQ8cr9C9lU+chJn/a2+ahk0sh/J7UetC2cIjEbOp6t3
1JbgohZDv+ZfrHGzQbzbytCPeyHK6d+KM1Fyr6b3JuVTsSX5PkJdGR3a3NKnZk2m0RNqnSbLW4UP
OgylX5gabftUPoDenzCFNS4mIrQgcD9bviVPkW9DNmHKvD3j+o1ODLAXmYUX6KwirVwdmc/YEAen
dpSEQLK7tkkMxFniRvNy00DW/3oQa0kEUnYMsNnWIu5pS3tCfIg/EOQSyiw5dfJ5ioS12SUJHFkX
MXpcjX4VN4AhE6102hHKu2IOr1wWxBZw/NhrSlUKgQwVN1+ryO8LOqZJ74YAZosuBuXd0qoNGeks
ojfKC/YPCFvokmoaaUKEvUFly2B3DlXwtMLmQFD2PZnKD8FizoAIK5uAk4RU9Ny1VaIqKdWZHdDT
rLrzDfXdPFqqaPfa5C87fl/tIavDKlA5TX3y+IX9WdTTJCVIaU+jJR7pHEe012565wI3oVLqL4Gw
ivZibmjVgURILbr76Z8H/THi7gYisz/nohob/TgxtiwzD2gJ2gE0aTKm6Zud2ciPj51O1Ks+4s5a
Hsp2pE+pzg5v+IDKK0/Z8v5XDs+32wn1fnxfd1WD4ue0x3odcQIGZCk6YH1jGhj/zgIpbz2yCEWd
D2rCFOyX7wX09DAk3qD/XBLjaIJ4EykCFxS1Pr4tHJiTWDdN+ZlIl6oepYkw6UWkHsxwy+VVC717
kpHL2fUTNQi8L91nu0WLZSsfyBpwSpVd4ckB2XJtgmpq8ZjI1dvaV6ADfluteqyHkGnhXSAQeynU
5K5V3p9CmiInVfIAUQnGP8Y1snq82K41OeQewX1ZZH0ZxB4kEgTLVlmzLylYjmc9BCN0ql1yzQnw
GOb20QP0SOfi/E8K8fVANuNP5n865GzY7R9sQzKsZPp9zL5Rv5GG0U1X3RqVYgKC3XoG7aq4fj46
TPYm+hxJ29EOcbZUPcTm4KycuVSGSimNQPePQl2xBQPdCzhWG0Pmq9VdZelQse5knEPmtUTDk8j1
A+MCuw+PAZcC0vYN4+fuka4OE82M/iDf3b3PXqd6ORS3JHHZmxBBRGD8992Ax5oYqY/vUJsjMSwI
G0QFLnAFxuXgDUn/rvDsE+Cam5Q4bGTm23PfKP/kuoaw6ytSCBuyQ+TTPoqBI3GTXRf9bTsKSQdl
RWMD5di3bXEcpRbEyRuxO/VRbvL5rBnbYlkfK0Zh4TBdstD1Ut14mJEsb4wo0iPbSxTB10dJZItq
Ga4DwMKoqiB9LIblmemBGpUiV5vGB7np4XwqeIudhspT+e74XQptvtiFsdxATGXBQZTUin9egX5b
3A6/5HjzND+fkncHNjady2zk2n5H0TqIfO7MHUOXhP/zx7/TsYQolJrs1tWrKSiyQBI4h+J/7qeD
a0GyZg05E1SxdL3ez3QUDkUWqBs1OZAmAcEdILfJIwRvKAEpHhJSogUre0YuEZM7LaprOeHVkVEs
ghNReW0Fcn8KEoDEdl5uTp4nZKQ3UhHlbaEtBqRkOkyt06/S50/f32+W8MaAsIo2tM1ZHd8v+LQG
yHh5NAmP1/+6nf3ZerH7vsHT05wBfGi83EqVOKvTYbcV0kE1DxhMTdwY/QCnxNenYep5NkEpZAxS
uEZ+UEHj5Wc3VXuS/As4XIiwgT0QVqrLu8LYqq+Mhgrxx6FPId9kf6eSpw0mif8xJXGhvQbDNhHW
9JtVj0QWZuU04jApu/WDdOGSAC1hesrEBKVb88WlKHjWbHmziWaB7j4LIlmmkkVfGdiH0VQYkNXW
sN15gs48pDQVGzkNEeGrQNlSSMlL3ybD25JEI4BwA1nTO8AxE45hUrU1mhHL2tdh/+77hDRWn+y2
2fJfTaUMQDKBsPNmvcaGOtez4oily6a2Ye68JIm7KDHMOWy9AS2O3gWGGp4iFMC6XbxWIl1czUDk
yQ7p75lA76IWSuwbNPj5BH+bkO28+aFRpnrDb00bRQHRDsYduGH4L1OkhSbggZKuY/yNormY7Ssq
UAqjP5j6jVrxMMjsatPoHZR438M/TatYGXokOuPHfYsL9oDTJHMly1S+BoiOfZEPklG1A0++kBjy
FzEZgamxVNyCQ3aK9ZfT3bZev5PSzs6g+aFtpxVo35rWRDxF+Loa6g7/gA4Woh+S+fbYqnKwSDHW
QcDXAXcPIGJP+L8YremBxKppx4QGnr4bmbybQOJqYvWirgha5gSsm0X97hSehPlJv/Lbl2iA2zS5
Tf0K9g3hDOWX3hLPPbq83YLspvSPLZUKkyjgJHwbz34zzn4pQ1Tztl5RSeyEWbDPi0p4m1JzBfpe
UE75SNoaoyVJTMnNr3tLjTHbXH1ejA+gMCKwE3NZW9etbevbiLzZ3D/OtEvV3qWLT6smuvW+nc9X
X1P/b268EZvfVj8BE+f5YGjHQyrcQRbdci/tyC2lhLprrLTcLUN2GypzYQR8fyAL+gad03i+App9
Qy1Q0G1sc8+fPgXLlZ9kjAOP1qzlEbBM3/GhdYBqMMjBzROUq58JJ9QWJPEe8VOatElFHM3fYfa5
9+SXhSqSxSzsHdaLoL/YIzyWb8X7c0CvwD4F2UE/YQXuA1a+ybV2b2rTuRLYhNaYUdJi7O3Shv2O
uex6oWuNFcV7Qnc0GdsgJhqKXT4UWbs4XTC7ezwLBLPFMSlx7RBJYSAj8y17jrLg/2RcmV39G3/w
ZKOYgb2O3g0YBUVU5gbplZyxYZ5GZhXwtG2nB39CIXti3aoqeH/RXmp4ileJV4FbTmogZuNaPKlu
ypEIu3pvlk0VdRY2eJow8pj7Y4fUEdXbEBIw+OcBosmggUTVbCUNzBZNy9W1qAoTbdAUx8DvR+HO
Q+QFM0dTi6HxX1idAOk45ZkwmKR/VQye8v3Fq/t60372Y9uSRseNEQNgCMOQ3cHV2310bXrMB4qc
8MFYFAZLKC9Vtv8m10IOQvl6Viwe1G8EAYq95Y+InChR4Vt2/JDWqdHZZ9mlanP5r6X+Yfwez9nt
8zXGEIQTZmL3atH29g/5nVe4RAEXazrVeKlhtXEmXE5B1YW01ESZkadaQzDNzMQQV4leO0FleNUV
YITH+ZSjKRXRYYi1EN1B3RSEwMZRadX5g+Z+T9eJbYW+827mfeUmC+glDS/Lxj4YibZOgo7IezcD
98c7sI4xJxflPgb4SGydk/Fs697926ehAoEwVhN6X2JiHVkK52sq8HXeTY9ykeVqkKvupqaXHCTz
tC9tnspezejLHUDmbbBXFY35Gb/CZIXM1/09TBrlFH/oxrby37K+oCjTUQzULMvIo+GLRwadAnI9
omWTxvC8MBE7LUS8fJ/FbnBbLrJUHkne/1QCp7rYK+rrOfB/sTBA3TOBlMogXXKl++99KDXvq5pl
Jo7XFmwRY2IJT2Cj0FWye+ml7UEEIPDV5fKnFfaepXRq+M6LYQTmfGcRFTKiobM1x5tqU/xi2nYI
RZS9pjxRjKhK2A+znoH+nEoAOamJokkekbihDAfKm4Et+dYG81yl7Mf5nhQcWTTNJtLVE+m+t7p9
JSg6hbmRivDPGVhGP4BbnClmqPuznqYWjbVb2bcZRszrUk3nglj1APmBMoBVtRF3M2t1vWj79LdY
Hmog6oMVg1Pu39yw6Mj3wHT9pvzbGuAuiSAW/j6fKBnz5CJj7VLpbl8q9MUfPdo18g82/30DxCwU
YMKpx2/Y1EpB+2BAnm1fnRBFprQzlmxwBmTMj10F3L05iSBdc7fdVx3a9qOytP5FcEKCMt1iYYLl
3PD/oHggxlfW/fHAFF++yTlfBzrr8GsnfKTbOqT8hiL7FMAWQdHHBEXgY+4wyrMY+F3NteNNC+4U
I3DnyTbAYH8nkiucoBt/UGidNhzrhb+GUdzADI1g9lIHCNoB7YHsXNI7p3oO56N27AWVrDNFd1vY
yD6YMatYezWGwzHSRPA9cCoRW52WEErPA2E3ukWCv19fnyUOBmA3kHmFjzxkRcs8iNRjtw567y3u
lgwhcjkq8D/vUeWMWCkQQYDFhijA/jxjChEJPKdxbeEh+Y1Zf3sIBBxriLmlpM76rRgQu7yBEQhg
F2gIdEbXCqpGzfG694x3YBnBK3hECUS81dPkf0I7qaZwk58FZKrNzzuna2G48/iVu2u11VXp5Sms
qngMeFLIcRCz/rMT1J7Kmc3kxF1tnp1M+QCINjg9WJPkutz1ORRMrjQ6R9M988YXG0eTUxtnQCft
CxjwhvnphWqPs9Ler2kxxmxvsV6lGl5DHxJKVwFT0911tX08F7qh1/62z/GKOkruNHCPCBJoAuNa
iIWMva9l9lq8AjSrY09tKV5ABX8bSKLb41SZ7V+JW6pNd0GzTnlUPRQX8Su2uxCvFJDDfP0ZAsBq
1cU7WAzBhKFuuviq4REhswyYH4g6jwOTba8Nez88UaJeLMz5vJ4IiO2mt12Bg1ZCp/rcf6Xx1+6g
TSgGEVZZl716xjuziy+GpxgHJar7Wwx/R1idLg4ew+J3+t3YKQwJpT6WBGuz4Ts54kKPBGisJzHV
P6z1iJ9TM23fb8YDhY7RI1UaZDfURTWpqm12BpXZcL2vrt+zKoNe6ZdiWdEm9MtVGg4c/So/bwvp
guAB5OLtNtb1xHZ5qeXdBHszR0mg/K05sEYHIGbAOunbwG9BU9+b56fk2CPfK34kVdDhXTQM8LTk
8bHVezb2nLGwlZJV0ecqQ5EzxEU9KxNImBLC5kwJhBpPhaER8BfpikAGXTeBksSoflxMZrAniOlp
fo2c+zLS/55J95bFJldDFAi6fn4PaaS1dkpDL8S86WRSVbC1kq8yxBEHLCDWmttrqfzOPlDZ7CEj
qKPXB10AzCLbW0NYiHKDW395XXodzMaQ5NFcrC42IrJcWOrjtZobk7IAw8yXqiYKqDX8LUR4Ovo1
KCHh39iEYPsCoX6Qsc+g7RFV0Owyno27+oBrn06Zy7pZgd597mj96yL8uIEzzOJZLPtBsiOxdnRC
tDatZ5OXPc62WFUeBX+xOlu2sT6jUmBQOUJn9+XaMJ1C7KAYQIYZ1+jcz2TXm974eB40VJgGjh6k
2CczE0M/fvfIMwiFAQtoHQDjzd18Hsg5tX/4avYhDj8/ESJTXFCt5tCXexeCk9naHHd5v8SirYMH
/JLgSuUMdfsWrrpKLOLiGgfDO2usi1jXU7iQxTbQ+X1obMdldpEbHIRtRzzQkWxxMkVe1mg6wpAP
iQn5sdcbB3Mh5W6RRt+KBFamWol2CZOBYPYHKJxkxTYghm2sH2jTma2oWKWKkPn0KLxWMuxbVz47
Fx1zHNOoAMzSZVMyVseRl0Tvgz+WLLpnbxB1muRsk07C8uhBVQOfWfa7wxPSabIRlEo3DNE2M0b6
ISv2w2BNU/LXfJc2Hf5333ktBmf+3+9oZDGCAvQ1NthVWJQvN4ndOXDFijujDzDFT3WtoZtIw+98
/7XfLaae2rYDomM81zbTvRPVL+y28rD5ePR21GcjtNNVIk4Ne41SMXo9lloLnRS/wsoiixhiUZnh
U9qwZuAWar+Ln8KcQ4LP4JXIF2NGuvBmku/BmmqInkfLUTRATpB2vxpkimoAZhZ6LVG9llU8LFD5
F7reogM93tXNgMAeCL7oRWXzuCZvaHpFTPatNBgKyNkKHHYwJI8JjaVlpZeXPS3JUd6GctUwlPb9
g78tp+DaeDT2Odzu+HyNB3N7zc7Lat7Dufvjsh5wck10xPbZAM1jOCZCqIbdZp9KZPhVG4HnsqAl
i2eSpL9JUGWL+dZEoAqmeBpfYg1F0waZvPLXyQcIxgYu17Bfetk3WDZT+KgcpFTmT8bIlBkT1EOY
16NJVTKVeOHxFsfxIQppWyHzNQyHw65EJcrCvFdgPDkY3Rj6STDJO8Zuluia1QWP9pra3yNYkQ7x
koo+0/OCgpdvloZC3E1rSjUFaHVvScBm28BN2rmL4ezZuw2JFSDjYej+QDC9hdq0gVkOBOW9ihRH
2sxvSfQL/cDxLR77v+EZrGa6pIkhFHFMj8lLDCxinMGN2J5paGhxBjuh9Tx4bxriSD27dcM0sWcG
ew5jWFTeNadPmrRQ+7V2v15LkqPCAMeGreyWpCARBIijZ++JQjTwPojt0L0f+x6A3doRhg9qFMI/
9ZQUPx47TPqsbw8votB8h28vNoDtNB7CKT3dkyfwraAy8k2SDaIuK/BZjJJVoHOJv3pWI+D6KExz
JWmdiz0gr3Hev6su9KZEpyVmkU4dJrmZZ2huMR/i5as+VNd+Ocq8qWq/NMBq+2uK6kU7MrXqwCez
/cjpvSXO08Vhhkc2xHgRUE04cayyldn4AzQaPwmuZG/p+fLqmebLQ6jCaZvfOYQ2IekAazwmkHwU
qZOfJ6h/Gw/gB5gDyL6QyZrzXuzkEIDHjx8rrY4Dnx6Dt82Cw4F85NWgCCxI7CmgZIHFmVEA/ysP
Q/7IrnUgbdHPTzZePYdzDEnI+tbUNX9NmHV8Y0husazElLUdmDFwYRUsAvjusMNkqNvUXxV4fi5X
doQ7V5iSYJP9I3L1E7wNA5OUAj7uC7wbOBri6Pti+qLfgd/Aqb00ik6MpY2ykb1Bj7O+v0i89O13
/theSjs6+YwJ19k8DfhzdfPQZulz5aMc7CghT3ZETNWu4KFla5KayurEcyH8OH8NoxkLLlDyQoGA
9l1vwfZhfQZCOlooSQok+jnWB9y5vWJohGSoC26mLAaWnzsG8lZ+jqQL6Oa8dOmg/0//HnNMWaVw
15OivVNecsEgSQ/5v1pCT/25yYB+SxjPC5J7Cy5/SVPG9KSXUS/Id+73Js6RpZQya7ig2Fm+3cg1
IfPFMxa2eIBWUrI+o3VWmw1y2IuUTPJg/3wrZQ2TbdRf6TkuUa1vIm9LMQaMDIKhqCD1PIDOkoO1
4/Db0DoCwnMbFcRYOB3DoGB0Yg0U1cN0laeBoBkvhmzDvhAVby6h2zMSIrS82NY/RVARwnipBa6Z
/Q5sYuHOHz091zZ7UbQA73rev16gOLDkmELE5MlzUdhfRf6XYLn2mgf9OVXaK0MrheSamDggW9RX
QDZ7k/rlkTLUD7OtHyJl2vAsa8WstB4DXAHy9riZPXkV8gIeR+fJbXRdihuEvAirDAXPp8cfBfKX
RZ4dButjm7WOysFzgAUvUAe4l2xMcF2bRLEClbF7saPkQAVv2Rf5Y7lLCtXm0qtGPiXfdEK99pMK
oFizWs+43dMeIp6dFCyspGx6AF6aIbCAa7lALcMcE7XKWrw07Q67ZZlvbJMasewVqUOfVvcAswW8
HRrf+NpHja3xIMdP4NblwsSQ7ElvY71ikYu/n8YHkRiKjnbCyFCNOPg5tX1d2a0ojpejIQ7JOqkj
+shHIuYQz46AJJt7pkhgT42o7v9ayc908Xf4Og5wP0ec5WAE9YbyrLi/sOvtBESm+Jicpl7MP3yt
UHY20oaSia+98ZmDiZ+TapH44oa2/Pia6w9tvu0jiLdWbVeA2ATz2gkuKAQlTFz7yzJZap7RuOfW
jU1CMurljrx91zWOuIQJu5Pj6DrKQb4CKTZNvWwS6ydl8FqjFcoUVmkBjYVxzru1j2R6nKO7KV2S
k1L3Lf0/3X0FugywKL+mskAq0yScUR221Xt20I1X3rYqhOoOlkwHL3oG8JjPez9b3+ANnCMBMgPw
QndFMunI1sA27tOTWAOLF2SeqXRXQdJpw9yrFy5EV0T/rYH8boRh84owhYK6GeFYR0QUTThPSv3Y
9WU7N1VT3JHFajZE6U44CkFqqfrgpnbv+RyifBHZXMZGAnzbtt1VaoA1rxL2QUs7TG84fAc9/wGP
ex1tOMO3h79oj/9OokP69D4CDYR4bt5N4ciCyG/l5ka/qkeTf90u6LBG6KVV30hbwWh9x+AfncX/
/ifsCu+CaphdnKc1cOC+Cn4l2Vr3z9TKY0uWaFUEklRC1T8+1AT4CiJrOji2EdkQqExzEslgr5Yf
VhIGLOmqVnGoJorYERGmNZFspYRpvyBv7c+/ofoXWAMA/pPFS37nS2biinwHkbfS9LtXnfYbxwRD
Q2SHDRYbEhQP71hlQgh0vVPxyPoN8u/gU1IGbG5FLwyqx2hnJeylD3SrlRcJcRvgoZBc66xCXlxL
cG6shpvwg6wq2YGVZy4SPT/5o1VWHl/mxajkXYfTjsvcTx6ED8015tP7bRqKqp6qK6jEqsCZnbeG
gSFc6xnQAJu/iXtZPdbKrHOjHR0+ZA77c1EVGpeJkIdhd7kwLQ+2ZxhdsbIXV47gM7eJvJHEQnAm
0JnelMI7e18cVIUIYl8hsSNIrSD1JvD3mPPBdp0G0EkvhTPLLVN774uoFLjb9vgIz4VvTEWwOSFQ
d4n5ZC25LMdWBDV5Vxz9tPubtWyIDLfM3S1r5K/xxRfjGWVVkbzz4O6H2gj6lZ/jLEpYkwpzV+F8
rUTodVte7PT5rA6fNfrBF+pe/HMu7ozanC0NdQpZP85TijFBa3NtjuqSgWP2RIUWN2UxawKMdjjW
OKWtJXm06tpbjuwI+iEHe9NYEZn991CfH6ATRnzUE3DY0d5Hb+r/jTe7OHYrh6R3Ld2+JWegwj4c
MQkaydF3CT00y7S/47mem9obzXGNIYbtakN63aGSVSfcvRMWW4EyLjGqlHKl4Wvv63t/1E4za9v8
c/pa216KH1ciHlfP0IZ8jjJuxxFJzrh7sjV8UMFpHUCaM2GJJN8TbmthLl+b2iYB0IWWi8q6q5EP
y4EkEMN2kivVPHWGHnCXc26+bUhuLB6Cb34nGTs+K03ntIX9oP2Zei4bRa8+BybOj5efuQpiRhWm
lvLlxBOW3JZunXCmFw/oBT0Gv+RylyLokovstFeUaY5f+9X//y5hU3T/WYNMfvfJw0KHfnyWk7tZ
ZGDoFJpW+jYtH/LLV+Oje47KGHzgRowO2QURU45nHCkKbV+bQzPAC6LknuoDg+0vrlc2KlT7Jxd7
h98hyP0KeMAf6mnsNViJ9OIad5h7ViKkDYa6Q076XfElpogX7nt4rp/lMohg0MpBFDYFHFk0d7/b
Bdqwg0v8vn36XH5eccU+TEwCFcRTCVVnJPhbO3h5gHIkzN4zBS/vKbAO/TyqDXOhTlh/sX6l2ZE1
DrLGHYLNKfcoJbOs3e4URQmOroVXPHniuaXKhx46DgWadj8JlpEkGixBNHp1ugeQuVqZJ+aq3gkA
qHd3+S7SSTGRjFrWB+h+7LwquCxdFX6CwTVV/CyIBnHJg2wivVoOlwAObXDmlGPdPtxHcQBe8JR4
lqc0UtmxPZG7YgK8YXw8bmJlHkN3Z6+RBsCUFyADXjUeQCQhWFgNbeYc0ZX72obF974pH61DdgHF
x1X2zZmLU1xZoTdGfheWIQZXJB/B0OHRYDYlr8npx54hCVZB7avR3OFjwuvuiKMBzeIVHgkBKzCd
aiZ2ASK6Kro0jlwSO6NZs3bcwVui8faWf/oFn+xSz4CSJpTUGVWfy9mWgydbouMqA7VEGTkpCCqP
DoUng2ExmGlAp/+9MKncSSsZuPpAwOMVFGzd7vEk9dfPMzuBOL7HJTpvmkZA8p8AETuejay+HnLm
v4IVps2x3kE06zL2qyuJ4qBERbV1Ozt9L0UxEVADi1FoGDw3VTqPTeFTSr3POW08I9szQInkOWPZ
JC6y9rTcmYnEjhS1IpEKz02ROzos1FoGf5SnejUavu0XIfv8qQYftXuOeeh8rbSxtHfFjTnBAEMX
Ig97OwNaxirXZxXYhgWbtCafvdb0gr7wywFAp7niH5itM1unA3EociCYsUtAeV/XHP7Z86KlaX4K
Kp8YbHGC8mw/m5tOjR8Ko3RFgM8FszZKTr/x8UslHniS15Yc+YiIC5UH93dDA/2Tzk5WHCN7CeFr
rmgP3F/sY4pMeb57u+c7qeIBNjwtgVNlYAwogXhXtecUUED+vIugmWxOEJpA7hgud4yRJNfYgcyG
76KE3IfzbXgRgMRJkgbSEam3lEofq9CE82oR4lyd1Yit2RoU7J+9BDcnYG9ji4kiu596Ufh3ek2e
9KV6h9QA0zjoV2MbljgXRLBt8VKMKLuQkWyes2pf5yIf9nd9o8fIMiaVJR2iYFMOweRy4y7HIXN6
wG2dAWAp6qWRck202VeecB6ef4YuBsr5W0zXJVdSQ//0iXuNYpj0vl12C8U5Bp1jI8U108s3FA0t
DT3Q4Rx4VlNch4WQw579I4N4Fk0pLqE0hVpUwupycPkGwpT9SWntxSg3eYLSPajxXU/0os3mAbqS
dJ7xnwGp81bBXpKjJC/V3AUIcqcCs+y067goJcGPREvda6pJkavyXQ0I0Kv8pKG2QxhiwJ4rdQTI
6ZEPJXs+c7xYKoFnbuQ+ZSgBYPpXa7hqTsSv3GeFWdkLvnV8nnpn2Olem27PjvVUq9AqAUT12G3d
tmK9HcJ+pQsYf/AcBWN8ZVv003T86xbj/cLbb5RoAFm0RN/pfR9OU6L8wRZMZ4YmzZxq39iMx2kK
LCOeNJKMSWUlSx/IjEl3ptuRHoemOkAtXtnvd66AmqPReKbU/0H0zoUp8aZL58qQTpGfJ9sntAzD
llL6u5MAYMW7qXV7d2K8I+ach8O+6Z0Y4fZFWk+JQZUGb8VU+U9454gDa4PPDxZCGpnfZ48FipYy
hopMtge1+zE+3DXd9RsWuGbFt9feqIjtolZFlFf5Cbht+oeJY6GRfRmIUOjfXXWAKm/3TJIqi0Iw
TqqSS9fXTlcPNpzPXs42xu/qNdr480WaE7VIg8uWfe+9VBesB8Q4mKIlCvzQprrjbtctWgcq326Z
tnIdJHyGfrcPPcxdOlxPu7KHy3GR4TudBdFJK6gfXkNihsvQyhCVrBpTmDq9CNLByNWSpeBroDVD
fSs8u5mfvZWU97r64UHtnstY65p85siNUe3aLcblDlGhWP/k0is0UslCeTmAqZX/TuPmJdcTnb6H
H/ZI/kaX1iFqvpOoPXQjRObkmfn8/A9UASkfgqAZBeNAfYv+mmD+4lvgV2FQEpstb+mv5Bo2tcSU
3sxnxzgx1uyEGnP1GPVbewbDd2vLDu4XdaAJh31t13nto5dV+Wc2wTGeUhcJHVL/CEGJxhr6HkQf
dWZDOwOT7vDEPnIxHrK9VjOsoOysAAc0QQSkJfr0/ez3P8Vr2BJZqtIB2hxzuoBqRK/50a9StC5a
6Bts+y1qzi01M/bAaTq0cUBkwSMHf6gdxn3RZ44pYpfAhrSg315Yzt3LMjltRfJDH9PCuDsTNCjK
yz/u+540uARRZpQUwlYBzkpvdS0YUptmgrRG5j/8yzBMWxFZqe6iz+j0rVQoXRWeMWX0ShmITdbx
4uTCUOUI1umi8DKWLpK7+ZUQ1gk2kb3GldDuKCF9Lmo7n+W047hLAsLXHh9KkMKphwAp45/2uCdE
U6lGg+EMfO6aOUWh6W4H5x/+XoHD5evFmuxz1Au2cB8VpqXhH/zsR8KVY1L5sif7z0JoW+r4BzI/
o756CVE3inKl1Wz+bH4BKdQ78PN8CW6tTnjzSQw23o+evmEyb/9xCe6txqxFZPPFMgwMQp9h8NFI
rBzIotwFTGiGrCjuYlUar4M76+FebhlTXj25ihRzAwG383wrcd42lNXA1WDes3ZBED5NtzAnM92f
eUHiyaPwYoxgQL+RkdfUA4By40ogYFezfXoIf7sWKTKHi94IhmTLE/FR1s2SFi/UFqe+gcV/wYBE
KRUytndGoz9GH/xklQNVwNqlVtFzKt1ccZOg2kofVg/4Rvs1UF9tfYhQnr60hNZzrHFZOfy3Bh6U
dPZfEmm5ezEGvkq+PAo/1D2l1J3hnmJRwPdgT8KImjXpB2bClrcQwRo4oGnTlD6dA74/I2IjJoyT
anrtIuVC0AH1IiFbxFwigaFANT2n1Xfp8WgKdZaujA1hS+tweDWVmOA+sTdF7jU/s3wuhSgvD29V
9oqYjGLiaFKsnRt8bEiER1KWM3uxTR7QQgV5ewk9YAhXDDOYWukm2eHAyAtsOIIIDLzlMdK7ROIS
fMnttBv7WxBejeGdHhyupgpLMguLo2dUDhYD4HoaI5d1LRtDGPhbXSdtj9uiNjY3PTs/pSBW2iVQ
ltIPn/w+qjSjvR5SOp3GX2SsP3k5fuI7Vpfk7I7jUL7WMIG5YJq7sEzgm+isR8b5X+uZb3yg3aht
HO4358orI7baT84N7qFNOUVeyfs/Wl/DTx16N+YSn76Y+7/a9cEbJsSeI43OO3/5Tp9Qd+Aubfw4
xZV0LeulvmXK1x9eiiFXlLNQoQ+JPo95nZHJE8atbfW+1mM3zcWolzWLNTiE2GOqD69gOPDMiZ5d
hiszRO4Y8uS5ZGvkMJ9ECEUfd5VQPzP1+sZMpSmuj5QCBP1llk5xXaNHC6rLOiuchmbLWMYR3Sqm
sim+ZZdNCmfqUGDhHrbTJxLIEgW/+3sb5xzOexjn6QUgfcWdvY0gWAAX6f59b6JJWXiExRbctRiX
Ja05zdOpTa7UIAYEadxJaADklg30vjyGVWi8A4txeR2+BAg3x0SW/zzMYnlBTRR/TZbJS8GffcVg
mwNGv66g/X4vSL45PfmMVPP7JMSSCW0WVHtSG61ypyCiovZeZK+j5Xns9Z3lt9xwnvepTIwc3qbH
RtjJO5kjSRcIJr9hTgEAeogfCiAza/7Nl3HjQSt9CaOfx7mIVFPwFpCmjlmxX8lV1OVOykC9T1KE
W7o3ggZGobkiLWBy1BrGIWmhoAjnRjc/zK7JeNPLGAQuMIyTKKLNhsWBPmG/IzunL2e4i6Mb8Pzn
KVO7ryLTBf5Mx5G82fqqf7M0WWroIfhCRPw5iZLct6SsN9HiiDnPsaZ9lnS9nDtm0vUiA9SZ8On/
89N2VvyXQ2wexDh95zo7iqJKRuWl++nmayPXthHEdsApBgcwcEaklbfbNXIE1IxO1l63QyOFzrPn
CiMi6O/iANspij8cWnWpF3t2mtP5MMYQp/+EQVwbYvhCGwDvu8PhqxojMaSXzidS5ONDdaviBRn6
vKqzsjtghRH1V1OjC5gLCBUxn99IAd6LV/Zicj6pQbcp0IcfVhYR5sY2FiniepedUacTInmbWUPK
ZBKP5p1gUCb7H9BmcQaTxW/zacqKEWr3fX67LZ87MmtVcfKQmpr9cfZVDhWESdJFdfd1v2Hi0ZlK
rsDJCtSINS2WqOvlolD/ny5ooJsawppBVti3qvIDY8whijleexTVc319eyeECWH4GqzHEWyVq5+t
M22fD93/3w+sPuCybnEgIqjWNcOqGFSK+vWI2YQFwfZNDxgBikqBmFxIV5owQ+XIecv7LdQ/MzQ9
2iypCqgAtTaNtF8nyvaKfRkX9o9166+I6WHDi959KLx2YA8yRzblzWc79b8Q5OgI+m4Dtdc2i0i0
UpSg0j1oVpzvMkLX2/ncd+8GUogLGrpygoU7V1dAaBxdikAd2IsrvO4l39ZuhWTyXkdaFk5sBczo
QdJ1RV6CLCm9sU3JFBWDsQE0ZKjZ8UrvHoUlKy2QJOxihTItR30NKhL20UHKlBPrIHhfRNTwpeVC
cIFW3tFdbjuHk/jy6F5LNJNhLCZIG/k61d5I6HyoplW7pZFTwjDcLgCnA70JEp2Rqs+ZhT5p/ln8
4gi2xg2kpD3S5M5y5xfYV3HIhEaBCp0Hekg11l/UMNAdWZVWY94l+u/JMRdL8oF5hd390KsV8YT8
m2BrMIoYvDN49oyL5pAGXbl0MFaFbphsE526eu2sseHXgf9avGuQVDW3hprAmqoKpbQUEsPPYZhu
qeMRGR2O939tuFCN0TULDwlAG2at8HPMSoDy46JKV0a4JN8FkTZy7/Si1BiJ6ULZKSAWO30+Ldi5
hSv7k94f8g+iAXP16kPhBp9dandYJ5Dq3rmY25gjcWrp4W5t5jnn8uVOcQaJXWd1GP34WYvh+e8b
1vvdI0/JtxmtDkbBUfaKDTpNPPJ2lzxFqXnIXppD3nr2rmuZRSmkX7Df3500rd/bgx/o0GCEc8dX
8/0Wi5sW33osniWc3peGszU4cQDrp7T5FpoIpN5c46BUP8nb1x35GsP2V3ix5+NEm1yHiUCGGiDo
29UU1xINuXi9Us7uFTXPG0//sYC2NGSPrugdjTYCEU/EdD1IxgQirQ8UxApnZ4WLgcJziTPF4uZd
r1t35yxD2lASHtlokJqF77x37tVB/JRzT61vXF/N5mMWO2/hu0YD+8+E6QIJzOUmZLm7IH0gZAee
jDqDNjcHzLKOT+QK7ymcWon4kCF6at1MZ+yyKbG1xqOPU3YM5pH4g/URQd2EhuOFgdvuuVC9u4Xr
0qI/6e12E+59FgA/5W7yVMn6G/2wZX98DQBQn02I63rqho0M8kizj+njD+ytustcorMG0atHZ4yD
DXEQSiTOtX9F++EssgZKx313dUvkeeukBO+UkrjuswumOpVC09+DoRQXC1oOfCMFCgI0Xb+cszWU
tdm1f65usai9hReFNk651Hk/+GAYtF/J98kWAzFwnFeFFV37eY+N2BiUpFFYEgr9QC88LTULFyEj
Sd+EiqIVLwkd11a/wk3upt2rJmZASIq30r1RhEd+7DJ7qyGkpQTtGRYTGfGVHKqym9w7OUemKXMn
v23UEnZCV8mQlXz7TFcV4DHxs2LSkNiCdcRNBZwvfEJy2P1dCxoZGxcagGOulHiKeLv1EUS/9XdS
2/BrhUpr4l0rzYImMVOAHpoSxDvtGitRCswtlF436T8FV2bHV+UlWWwlbAxON1UTviIcU5lESR/m
6dk4YIUEYACobKe14lmFkBYK4s7NzlJfQno7ovopLplm6E+/fQ8dH5vfPId7YGZCKDAHqqQ/HLSh
Xc0I2ytYpMAJpb/X3JTAmpt47WHSGAmbgPr0p1ZnWAGI0jZKj8Yv19B/8cT+gC85FItTpSwN37Gr
vRInukqgrr8T86N/w4uYXdbU1/Wq0LkQBs35NJW1tgyDkJiUhvRc9dJ1GrlMbVmu1a/G+PGwhfMv
weBgrIDrir8KXjB5Pbe1wHaVd44f5LR5i2yy+EMo8qnm/dpBTrSTez3kaQoeBHGeghvo7UcJZ0fC
ZQTZt/BUEFvyEcLaU5/r/zKxe87pB5IqJ9fa+W7b1THWdkOIsTc545FwosZg8+mY3wFsM6BC7knv
Yp4WtdtxQteEX4nmBQqAzTE7eGiA17+3+CuMQr42tg+lDdeW12TTU+GNEeWepglbIG75RL2BmnfS
G9Eryjn/PhCrpFFLHWkdRHGo8lwiw5qMO2B9pT/+r6LH5WujrL96yJZvv9FxFeBgO6mbNcsYoyNt
g+mvA+bHrTNfyl0AAh5BfFe2uH/Kq4ifzl/lYV7Ghntq72nzFfo4tL89j4Q7tINhjnCI/jvqZI0m
8UKDoeJBLSf8Eb5KpGSwAD/aiSVQwrvf19PbI5fXdFzv0AeAy0nVT4dTXWj6b1rd1nFKYoyuJBv8
f8OOiE0PQ4k6jhEdhbe8bZZeLGDBqBZIxRkfWnf2MT4TDGRo/Nz8c9tiNrhWXlcAvxlQZosMpQzA
JRRMQZa8inZY1xcetI79sVxeOpo3PPyo6xHl5R2C124qH4T1oKI9IO4cgdoGLtlD1g9a4gBDObi9
t6ctKngXj1uV5DhUgiCufIHaY7xRdkhp+TSkEcyX7mmQIVvVHKw8OBvVJNmKtc9USmM7r0tI5CXx
fc8XADPobKIqZTKupLoj5U0ibQLNtEMQFC/6XJv59IVD1wn+UOpQzs8p/+JpmRQZswk8odGu7afM
3ui9JLAHKS9LRh05wyMRj50k+srIc/Z9vAkhBe/PzTCm/l7TjsVNlUjoCTlc2+cxcw1rK92mQqgp
qynfv/yJyNE1HC4id1Z/jj/0OVXGS0Dbwlimjimmva9OO4QEKuPr1016aSo1TqiAVAhhtkHDKQIT
kqZ2Fx/R+dABrx51/RcUo7Bs3fI1IfbsM8+KPgO91/fkr+qKCFQu/NpOAeTukME6EQxOMmFFQ54o
Pzq9pVH6+vC8tMy/E3uKnpHHqMVZAy9BEc/YNqF7/dXyAkaQ84EsNQrGJInz1dobVutTMilaP6iL
YVM85L/v5fjDzVm+Iou3a8jRdyf85Y9xpeAcj0wzkbrl8tJC3VR6hjv2iJodu1FOTHSeGbEfo35v
w+rprwAgZs4CDgJrSTfmak7JTNlflkTACnTuZ7x++lr2wSO9EPLNcjHb1f1H8zeoMxWaJAnQqon1
RrRfFmdVTIn4q+ukUvL6Gg/eztmlF7yqPamkouoLBV8ZriKyaJ5dN28cDA/6s9ozlG6HtzjEa4Fi
p3J42dy+eGuV7CLllxnQeXl4Q/fHnWg5Jk66TnfdzfVKb0nQ7dZXmcS3tqZ2sYdh4Jz0WjmMzExD
2VdmJ3jQXfq6bEQ89+9CTF2qJkFrqUoaAERGGiLtptN5dMA+IObT3tk9iMmML7caP9310mjTEgY3
AcgRoi9N1Q4l5l4uvV8mLX3K3EKFL0nDUkARy2CBLAtKiWkwzDHegLcvWbm63HrDoUZRKMP0Zh4l
y9dHl/wlrQyTPgqIkSGp/M+i5UllLoOHY+fuyNVMDhanMbwFyCq72gyp3JdQOA8MwQWV/P2YOb1E
WfZnH8n7xX5zHaF5apZvZRWit66CDtxQ/LqIzXGzKzGLA2OHDTHO7cSVSDpu3vRi9Evf/ve956Lf
jVxIIAKHKdURZA1HjBylmuPri2lgCObz1/YSdg+/yQVYkY0Gvpwf10fVi89FlXkmnBE1dCZBT97U
XLPliievbn6Bp5g/e/ghAkBUQfLgJAJ7dvVOVydC9zb0oFysXdvVO0NelAnlI07qS912U97lzeEp
UODcEuwV/TxGlln5SgxLBticwPFKT5sh85R+eIeEQLj1IEA/GGWTeOLk4urX7SkYQR/uMa/BQ5d4
4wNCcKG97Qrq8Vas0Wir6dlx4KIWg9Yk3uB0s7u9MVXKrIHMOREKTpUHRhLN/+oOgN3R7GSp8BnP
c9IQEv5z4+I9Fnp7/0Eh02EbPnp6uwzXbwLg3i+mlXZ5l1WcyHWP81TaCDgZRHlFP7Hu7Cs2aTnB
4TpdOd2MS9freDKpXevJ9rmuQHX3SbT26wBCtsAyrGm7qQhjK4a5dvGK7YefQCKipjdN/TTFZ1YS
WAwwpgp5vQfYEuVGPX5y8s8iDqXpH/5kmSpKKXQvu9z4Zr45v9CfoEStZt8ZW5Oj/UoZLBX7pHPd
aDxm3EXmKROdWiUd763vf8VVQArhGzdIcn75cAnlpji1QIrLumRJpEi66i9kOaTKK/vf/c3CY3al
jV+C836iBP65h/BnM6uf/yGFZEAHZvUpPillKbwMTz7N8x7Y2IOpnGVxTQ/pQIbI0zUEWtvS9FH3
3RheRuWTd+uO/+DCNX/ucHdVJcxyLdfmSkYByhmgcauOxF96VrI1iKTgClXzwAbBx6aodxCzOQl1
OblGIXrite36TqjNodfKXIx3G7gp74/dhCSkHSMYiSb1W+6g8suMc2Trn0OJL9C+L7KO35hxKgkH
SUXwgR0zeNFC2uUBxVXLmvuY1RY9JNlZy3lAYrYMmBbYHzzUzOIYHFA+d3z4f41xVPTA5pCPuRI7
z7v1rtqgKAJBR4MqENbYXVkjMFWMOVm0PqzSmBO1h5eTubcOnscUniVlu0zvdbIbKKQknVT1ogj7
0MDfdjwW9A3W7LoBtq9f5r0I8DK0lXrwht/ieJPn1YELNIITVsSLyAICYSGBO2QJ74u6sN5ZLwjX
FtuDShZSO2q/ifYmfedATmSgJX7MwD2GwOLXTYIUxY77G7aQ1vf04ns0RFUF5SkmsfXl2Jpk3kl4
s7hkRcVeRMANPM5DHUz8jK82iqzghwPRvx1lilB5iSZ7/C7QqHbY5GEUnV22QPxYY0Y2MjKxqGgn
hKWcFrG/U/M8rnm9o+CnJaLzGcxdJU68lfOCSMGNnFF6oAybvLZ7SUAyJ0acjUFW6O+KVxxOs2oq
t/ygSEntZf4WA2O8jbQ0T1vqAMazML1BKPxYTvIx6jAT7LbbiaMcQvP3IE/G/C358QgYzbWfeAjc
m948QrcycIC8nnrGx/+PlWerPCvoOTwuCx5gU9DZfrsNiFKXKmsOQyXT02hhvaJxZW6lN36372fl
AjJeZmxiQQTEcyXLRRQQFS3Q5dyDUJS3/ybqMLuwI2xhONuUhtkN/Fry/pc2T8U1azdedO9Z/CvZ
iHVWrYofKzSJtkTQ5KiHIbVSBPrpdbtApNCu5BVOFjYDnlZStnZI3ExXhz78/jcqJd+Vl3hGlze9
7lnD16X02kysRXmCvocNtujGce0GnYYCwmD7Vm26K1SG5X/4gYL3t0+kg0fE3sLhr+YVjpo4XS0l
s0ew56n0461x5nyhhGEhU63zPd9JDSRkeL0Zazm5Nxvkw2D+SziPEIV6GPXTPBFtxY4bg3Bbq5Ns
zng/L7NKiUhjIMEAeQN3ohZA3CjFMExBWQWpIA5i9Jo2K8jYIrYKUZhSIzsOaWnFbHFxuEb+3d7z
8heRdx5CkjY2LBB89UDeqwUw+/bLNUL1JuSJ7Lsh6T6SJh+YF4HzmskEM9ODKOkc9VnhN28eJTD9
JnSPm+g52qtyJxvofxahKJCBx2DMm8szcHG8g6zGF9R/FsGnaHMResW35iUCCZkvI+46HYsZg+CF
MTZx3g5o+A/emSgDYRahFwer40NV5iiiP5YBKBEjI5fiGcXjm0cj93sxrPnwQ4VqV07ffMf22ngD
uxT7zzF1XzGcKTAyeSalillkoId0s8w7tzwDcD1YpDGL17OZIo5STNA6ZkmonfAcyGa23lTmnrkG
stBkXPa+Ve5kbvj0YiZL/xqCCLal7sUXEnp7pSSvpzITxL+qaPhIV+AUAt5E8bq7IUSWcbAiKzzw
8XA8ELovuyn+H6Cg8rWYBDUdROUY+Ph3Qh97I7HGE+RrRcQ6EHWhjiU0BYdxWt+abdouYG66IJFD
o4k924lhvCYwG6UCcNdvakK5ajFica+3omkLhxfHg6o+Gou5tvzJTzBFLh6qC8Rv3neTpdiRf1Yc
gUCfHm0BdTx48EAD40lTBWZmyMxDSk1KJz0zzjZVcnt1RlY7yD29A4rYcXIOZaXYcvA4pk2PFz8I
bU4dPOucp5e2jYo174xNVY4Vcgn6Lqq/J9jPCbX40cgR49VkzJzRNnhmjSAlj1OUQTblEpQjslh8
g9MC/QuI+5iRTmZ9HTvOurOIB684lMykqRQn5+iFXd5zSwTUXpj7o9/JfP+b2rBINNNVSqBAGYhp
/5BMDm+pDUC1CCxSdPtVqCmoozV0xc30QLkJtQAwAtRsQ1+tD6ATjoTwBz8bdaKjXV/ba1QJLk+V
5sVvjqjFOMCwg/52uuYUAGGBCe4cxXm8mWvndS4YFp/7xGKl10cdKQjHdkOL8EG3kDvmtKwXM5V7
7xsBQjwaEHR3+ciQOaATUGHbERSTUZ7/AvCmOhIy0cWeuUIrChQ6FYgE5gtBmOr39DEV5EIHzpf+
z2Jp3Sn5AfqAi6YbAQmq58uL8yZyXmJuFWzf9qAVSxB3XU7hh3YhBhzAnuoNvvw3mOBEdFmDKopa
YL+pCq9xkE3MpiLRWhV1c9KuJ89p/F5egc7Hh6OlCiZyDX3DCsItxwAAC52VCYjQGGcl98UVuGCR
Crq1nJKjrZ/CZcZJTDhhTsxdm2AChYnFtqFRO5yTIMQmlgmNLVC6HinHrj4h1Qcaw0tOZJAVJ769
jmO2RMoWiCKezXUzx+llDQhgrNHyHIMh7GzyEEjoqSjk81PtCz6qzVlfvWy1z0vUVnPmmv80cgLw
36IIapav+WsgDV6j2YgNgNu5vFC4TL8zS3vzhsDEEDzJAop37ilGgjzCBLK63XlIbK4LzNep9S5Q
u/tRtt1qhQXUo8n7kkzyN5frbuHC0rrs6P1rSPyh/7uKtsm6qqIY5VJ1pcZwuATbR4yDt1/9MzKH
+/cwt9Dda1cvn4S2l35NJiQ4uzVIYaLi4IsTzJQXjA0tUDAjo8aroOyCaeOKNIqGjFTM2rz8CXgb
Wen5ys4jtiPWzMWaRNANiFjrVL0KLmr/lDVF6meEF2uAbP6WmLqwCFy8Giz4WxxWSni2O/WgKMzx
PU6SG/9dl+nQ0egtz4/OFakx/GkBMqHkBHbHG2jOukxmrHywfdkvoMachUA7zkLaapdt1s9ulQab
UtaK0UM3RwUQocsKdDqpWZg7WvmCdzQLYEkWAeYfkrpguETkPpoQHCNx67qVaWkS9X+N88V8BoGQ
K+UqR/LW7PeHhAjCPtVF47MaXswVkBmhT6ZhY4rbCf0k9hkgKJrSmKAXu0/xz+dZOQ4mi1N/01cI
xxUs5mqhJYtoZAbPIkFXMxmwEZH/kefX09/FbwgAaFvh0hi6WlU/pbHRBpsO/F5SQJ5fUAyPVhTe
Ut1S17mRWeY4mFkZNaSo6bY4dxuQXctsh9Eo8diJz7H6Jm4QXuTk4tsga7DO5DighRB7UYhsL/y9
LA5uRsGT6SwoYT6FyJtH+lH4ygGCTnfR3CA3zpJB6W9OBsTwBCY6w/DHadFdqloI/2q5pyPdS4Iu
UaDz5BUkBJm872VlWoASiMQwDMfEPtBMisxVEt63AKmWpDBTcFEHgTzRgzHcPoXxvHVo6m8X8FWs
hdgeE6BXewqA8ku5TcTRJq2jP79dU7cVirH0XeicVz3+vmbLJj2QZmdXqbRIBb03M0mwYlh1w0+f
Qysq67D8FXq3r5xK4vciEZX9XvvH+nW/qqmoLLaTAmTN2qXFZGMVmzRx4Shi4cMnTf63hyGMXlJ3
FR98xbnZRVoIqPAtoCU+7FUT5ccunnU0u4GreU2L2sXsov51/tlWp30A3gRvUoEvQHcz0zaISrf2
3tQRtqj0kIE3H8Kb7/Xq9NwJVS6shrCN1Dev/TnBJ3jI5Nc+VHpB7rMNlToTd44YGKBdVCrhCXhf
VasrZy6RuiOpESqTwHeE4mJJPUJKoIhGkyppCyup3W1XGd7cS6KBOf659c+Kq5GHgH1GF080c7fB
vvy+lcFs385HbIvyWnByPuKX3UFP5C7b6DrMIno4a26EsBVrYe1JSjjPc0IS7cwNf2TXJfXI4RM2
ZEIOPComeygRG9jWG2CLGjjHx+PYpH4N5Tf7gdtsUyGy3/9gCpt2lpT4N9UAOlJWQDM77F5ssKqH
LXQcfM4JRjkPTEQM6Jz7y8yfB5b75qWRw8bI6GfrJs3uWQLPCQcZeHbs5wdnJJT7YiIHwbOFf+Mn
zVbwSCLFn32LFWbcE4ZJcImlJXxqH+dTipBTUXJAEaC4zOhZnbEPtsq8DOFy/cYu74ublqcXwqwi
u31ZlcpMll69EE97sNSZ7Qk2KaWCeXbcty2FQmSQY+cpWfEM8i59nyfs1bLy7GjOUvt2uok0uwEP
9etXARNYt1DcIPfTxP4FHEJhvY9O2haql8HbKn6szSwfsix94s/brqkTNmcgDOHiU7hwe8KU/hXq
sjP+WIXj0fQyxXe1N4qmqN0SrGWVFHtBiXmO782NStlTKKpmi+fYplP2E8V4vPwn6BepYnxmEutx
Mo+HLJ5fvXj8B1kv0jANEHJtPpfli72ptxjLzH5bRJDKhsVIE3KgCZzlDHTRbbPfaN9d2FUxzZMz
vkkaWgTHXKXBhLSGBRewWOY7pyx3/jJJwXjaYsDyqpS0F9nWcogVkJit/EJ/AEdFJqBX8wrwh/qY
cE6NlelYI0pXc3OSU2J+vEwNLGXvuUMgZITUb5B4Kn8SDDSnQwAnn3V9t1eTxrspfArS5dbvNJdy
5M4eb6z4wDq6w0b0CbuBTVbkEZwxbKQUDOE+THCIdJm43N4Zc7Cb0Zp7hd4Pht8zNZSv1KOyqC9b
0DL1eMJ8CeSHJoEthgF9Oc+HYx8ap8cdyjguABSaKVc4XxENQ/cflseVO+GOUavxoMBzaahkHyLZ
IaKzbEz5gAp4z6z6MFb0wUM2OPH2CNA+x89KWLyR1q24TiB8hiAvrGUX4GUZcdDRPZ+SYCCYXfMc
kxHW4GU9N+jR8qx92d+gh477cP1Pb8MC2PMv6rUqNh2aEXOk1SB8LiZRjUBswHDcDFCR1N8SP6Xt
gwjRbUEwQ2IXXivrpm/XZad1zHCHBDCEIN299SlqFKzHIGGRuzLBTvJ49Rm26CoXuF849eWHdu8R
5++BkgJSvYSiY6oHozc8un68N5YiF8VayYb/nPCs/6nSK4axZWMqD5elhLvOYuOI/n1KiwrcTCPg
bg1SaNUOO4gK6dFz8kM5u99Q/H5X0IYV6wBCCRjMK8DbxuoE38xz/MLogSERaKKSgr+WuaY/AnLY
QapGJ5z/RLL7cg8dMiheQFw30HpdU7Fkn90FH9rdRi9/04x6okpqzGMvCYW/vo2jrS7x/uLD8tvm
uAi9GIl5FexXaWvH/Xl4MRFiKxr34TboVgnDQwujA7r7Cvls6sq7G+QjvxYRo6y9I93bcnvoKYjq
fop7BpFHB7Sidy6tVzGaIQjZjabVsGG/yzyC84bjjd4XpUB0SBdNbATIVHoqSsvW0illJuOBuDDO
mVxJoBk13lUOA6p+RVXP05Vuaq5QYVuMsGvNfjucGRxAlFKyknXNO1mppkLZZg03tXo1GIz0qNCJ
bp0bvHShn37TH2J9mtN8lj1l3Xj3uEJ+LQJD0i//kP6SLfz7QK2yU0OKTZagWg7XVD0UQ2NbXCcv
Wy4At+LBlnCOtlx/PQ9+C1ZbdxYZiwppo+ON3/qUCy/PXcBNznzsIdw3ITVw29Cn5zYA+AFsH7If
JA9fflCGIHXaq6WXtxOpo+oD2WGzcewRujt0sB0LDMJgTJyksEUTs0ceNi65rRoeHFH5Ycd1mVYV
T1iC3xtxcPBGzW4J+M+bgT7U8LbZx5x3967fkSykfpGUjeLuwwUV4IHlABiPmNzU74cFYgw7Bpjm
4/p4Pu3ersZbf80S8r09VeZkcipi9gnGcEMGj+jLnjn/UjqlLLCD97ikUwUYk7HtZJ2Q/432htq1
ZV15FYnU0gQUF+KdZbcdfdKwiXya29xioiV3cRewirfCKym/NMe31F26AruDjV6A/YSqi7vL9JMB
BdZmNf9oAmcWPvQKUMzq/4+6N64gb+UOYx+8BfakMW/QE0xpM1qHMGpFYXU24x9rhIlOa1CkRSdP
aZydMfF8jHJR6q1Avp0/S4NlITPl24cpa+clIhuAgKP09jeUfuJzZ5ysRGOchhRGR7FYFGlSdLPi
Vznj/gP+jxJI6rWauNyNW3Kb/4aMJuz8D3T34weTjJuUt1TjkPE7C4+cyBXIg9y8OJJCX7FmE+oO
W2cNwm94/XWmW9K4ypeN/RUiUypi/mGIz4VfB6FdqLIn0or4cI7CK1efBl74NwnMQ85hMjLY7/BI
SEiorI51jcag8CPFnN9/S9fEZhIFem2atA5iGe1DZVEo+swHynUUkv4BXDUUdmMrm1T7DatUkkRi
4prltWqgaVWLcO1GCyGfPfxi95NYNhJIBMfr6rSRfKZlgbTbVI4PxBNmm08DLNEMTVv3M/04/f83
H53ssFNZE6uznUBQd5jdOaxLuBP5UVhVF98zElkvrre6fkDvNH6bDI/TclXTM8hQ8GCMFoaR/1Vz
cdGw3IongWVK9jfn9vFqIaqpJ8xLIwt6VqPsB5D7UvzNSUnUJ03tZnxg+F3AQH1YCLhW0+P1wbVs
mPKs87hdaqmBMgvDht2ApVOL8793NW9R3hO1f8Ckc9KQrGaPrB5lLHeS0imDfb2Qnmvred+MVzBN
jHY1n0P6kzl5D2O3nFSAgf9DJY5qMQFnAOcKetkfdRZeJsh1SrBqGyQ7061s0NafSWCNIMPeCH+O
XOFbq8jZp7OVdUMqSOMN8shgj0KC4cXZg0JEg/jabghnfh0BtHrgA/JKmPf15WFl3+wzr1lOc8y5
ftO9ZRBor47uZQPeH1VmTY0EH6tbXHzYBJ8CjLaeI1Hhm86MPwCbPGsQFa56yBFOi5gem4pG+jrU
NINVqesJI1GKEODDhVj6y8uZ7BOb579Ob9uXjRO9E7xdBgpFAmNDIBvX9mq5DdiKOuy/I+9Ws218
BPSNWAreAJnUkd+JkJ/M+xPZ/864t4osEtoM3JifqBZJrfsJmxF3oXBjL/YKB9V68YA0J3wE76vb
4eBel/sNt4o5y1IRTZVoJdOFGguW3d/9mfCPOb0P78fQjyyRakCbyltwoDQZxjwIzkXaXUsW+hQJ
rjSSm5sXJLQSUhPvxi1pwIuPoGbl+/5hH1Pxrw1c8ugmMiW6uvvFBYnp9QoWRAHKnIXMEhD+11cZ
dq3MtSlg6WxMZi75QhDJXZJGU2BSDnqSZ2QjdyR+OR+ndtn2s3GQO4likH1bquQ3xirLSpAbb7Zx
qd5fqXWQAlxKX0zwhbe19CsnKrVU7DW/nLHvH0tI2cmfrbJkMsao0B4EgW7EUytGI+H+71ZdDEUw
8Y6Sh0jF27qe2ShrhRw04w1Ma0A8KxQ/BFgnBdxHBszkL2NiP8O+0iuphxOonq8WlOVnktGpGUix
KMSXJQDlswT6R9zSr0QvVAEwbpPvhxYLKvJ5acup7Q3FikAwI0NM0fLCsiw5VBLeoGGwjqGcjibw
t7zYYiARbDcA9JCOQzszDFmFKuHDxhNjhXXY05UfyBVtdQiUAbSl8FvmzI/yvWdoTEQIoMzVB8MM
BeogzogEd8WI+10Q5FmHqM92eH868kXg+PsfABQSs6s2SYzk3P/9QwExZTJLQnhUtpga1xail3T8
vSKoJ+4xPmRIB+0pN294HR/KDGqIJ91/9Vplt+r4YCRPjyxfQFt6EM/pzJ4hkk3euJRDTKeQBHm2
objWev68w12/EMqXTuMrvFr7sVO4NFLW4GrkxKppFDcL8djiPe5SUbX94dcm4pWKlIAMeUlazHyb
aZE6/gPlfxMiUnpjYiOgK6Ufp+H+coal3zM7WM3pwh5kEK+pPgEpUrmxSamBJxso79FBqkmVWmjQ
YXTZBWeDEMBeLaJOUeCwHAg/32ZBeBxPAVJj7r8RUaMTwU842x4Yb6mCbLY+wz9mj5BIfjZEHqFT
EgxNFvT0IcpMIROjodyhvrkelNXk+CuPpWyDpXNfYR6q31K+TT+z3KGm6qDwVptgcNiG8wq5BL6u
jUtYYjRlK0l2tZfhk46HXkQdHbE+wNygaxMRHEQg7gKDoM6VvRfA/Opi/iqS9Y3gmlTKthA123LG
Qbk2gLMX+5bjrBE1UC9e1+PMlAr+e1lOj/03iB9jMwK9sHCapUDFQgZfOQKWcrRv6i+zFKQWo+OF
jPmAXNpwzCyfRpRsFhr8E/eeDsDDnuPoOxgEjTXI/u7w4bhIvE3lo5V/HR6yLx9T5CNR0nGkgDYW
kWsg4/MUA7pIlrxm8M27Z5SzRLpJbsoZAH6vXcpdZPOAjZ4hfa0H/4N1V2GgHyyQSw12C0/IVi7e
9ruMe41kn6NotKL4hm5yym2C3jDLqllaEQ3iOhqsrmEfE6bE8QxyfsvcSEpglKFz9yawjlblA3qt
T4RwtGL4x1hetaslx+u7VIJUWPt4hBjxS+/rPvdhCe4c+tFMiTt90cS9xrq8GSBfeUkWUcYBLR+f
1Zu+0fQ+OuuceakmvNbfo0pcXIGCYcq+gozDT6wNDj2nOWUDzcTkTvOoh0UQplILS07HmrfjPmxB
1TaIGy9E6pTvzqS0Sbp7f9/AeK2u5HIszdeMdhS+VwEzSDLD6TekNLECQpA2OvJ8FqE5KE00NZBP
aziKuS5YjudBzpjUPuQClSOaiWtZ2vbreLuSF76nsUyHGlFK2+Ispj/5MVSWBuioZ/qsyaBJsRdr
daysHyypaPaCGy6cJ4TkyCdQj8F89N1csDjKLH6T4sqBaiYyVWk1cuWsMczKv2BvIwsfb9p/AFcy
N/1pqaZrOtNPSKTPaBypSnRCaU73zXh9IKNySJczvr8GvihYpyAVzUvcjz3kLEfGAJcIhEC6YsPS
VRfVgEZOmHF1OPJ1pm+Cm4tj7CnItBDMG17EdzsUYZOH3J3bnYjDgKC00ZFJvhzB2xFs0CYt+W9e
wf3gPsx5e8Az4tIdJvTIQuXOXjkvA9BLh8IZ9qRBGmJyjAlWwulA6xh8H5j85+SU7yZnAOHdiB1y
AXm2R8woOtB/o0U7nrNOuz64Z9/5cJxLOV+HjYmIxbCfedfrBEqWR0Fh0mB7OFuOku9qyGKj6sD0
oQ4r5m1QxMyDIROpDbJspI0iuGl1jRIoXfNljGVCWBJhOFcQcS5FhjRIrC92HYJfMF917RiHBahD
M9jVyq2zliksf7jSmHuuunrtRC2PPatPt2G4RXGZC4hiGrtXluTJR3faW7ukWame/nToYyhPg65B
dZcY4/D2hQCm8rGpAeVk8A3ecBHpmOhLkyAo0ENAGlgRKrkxH6yOutbICGaQ9XbgKt7eSVZe+T/u
GnkS1YnsoHBOoicrGgUf4Xhr26wBeJBMjSnE4wS8u2qTG9Seh0qybcX+Lbwgj+7V7/HB5zLub/WI
L2+uUlZf0HOTkPJQ1nxHRDyq3AdnSnZRvf23YxQvU23AUGjP4K+wWJU4J5Uw9EUkFhTuSm4IwQ7O
5M2XCUhVsm8tJVYDqvXKTi6sbSfdf/Hs/LZuzgG88zs1qvh+uMckBIEtXNZUncUvAjj/z+rH0KQf
mqneSon8N72VvNHHzmdmnaBLqU7RSoCmUeETT+O+I0DccDV2XwPgs2cQy805WEzdIyW71oSlqhJR
xsyibmCCGCIY+ie9SesjkM8kOpEiVl5IdGqQBr/DPM0sjIdcYxDxV2/9CCMrDVm/TSTe/DMB6gYP
D/bfD9kbHolklJIqiX5WrXlRpvTOtJSoOMzHOmD20S0ZF+2nf90KH8m//GEPkQdi7xkvvUXCNY3c
Dw5TQ8ljl+38AXtPUIzf3Wxbb7FMLwxs373RFPcP4iV1OM3Hmk4a54Fcr/5HUn2WGAuejZCzpXhq
ertpu9Pouo10ZLWt0Z16XMfQuT8UND9IrRPkNLadeGkPGa8NToJSO1r+w4BMpcITkT88275xTJYU
Ts69Bc+3zhVA90BIobmAN/ispYPmAOYT96iKH2XwZOkQqQ1lRlb7EfUzbXa5kTi8ltll45Py+fyl
QvCas1Mp8o9XmnTMuAJAMf9+roqeT6pWmhaL7/TRZjvUvZfRqFSQ0F5DTGfUCvWQfM3AiECMnIvo
l90BWU/Dr7G5K3ZMjuXGjpdrDlo1LQxDV0sIYeE94FhT1AU0zqzDxHwyGqN9b6sGeJsj7WZ5NSsF
78zuRe1J0WRKHZ5s/ha/oqdPuff/CLiZkPhLP01Rs8DqTzaH8MkdyvzrwyRKtxrYEX2AwH+ua90n
AaZNsX0WNcbtMbzrMgLGLLRO+U/vOofhiamPfNcFojDNrI8onMGcQDt6wPj69+zEMaWuF47MT2tt
L5J8VzFPEotARQu9aTNEGZXqxsnBSL+s1tZNAPBfcyC1nm20zyb0T6Drwi3aN+uk6s3BBMquBoJo
5HwgmOQ2hfYTZYlRg55LWTfpheqwAPhJH2s405Zw7vfc9Tk193yAQVUUNGTV9cudI5cf3yHjYJm3
hoiyDlyvlIzuA+X5xi80eCRyNKJVvRZQ1TtM3SOVLFRL3cGkTM+KMl1A6lqJ5Ssk0fTZI6j4vkB8
GxxtvTLgno/bEGha1Jwx07h2veQIcqPrPbsUXsIYd1XYu/+Z5chYdR8d9PEqXhAnzibELAURl0qv
oTAR43cwpzpEmkoZae+0Cnuq58mjTVBGRTUZXD58BmaMiwZhA/O1+iExlxAMb7DG9oxLkWGDv6h8
J3t/izvYxLCjixbTOoJpDtiBtWgrqw512zA8oS3Jez26S7IELn8yMk+B4jpB2Q3wSAU8l5m9nMyO
gpSMZXpHgfxtNSisXs3uApz5ZG3m6mYw5X7/1MlLb7ga96Hn3t5XPoDLdk0mLSsr3nr+vKGxHtYO
G2ASgXKmug0dpaH6lwImSQNiu7UYP9f6LpDP5Mxq+CgxXsVmXoT3gENnWcjwKRSGAf3CrphOm96R
yIo73L6eCg73Yt2KZ+NikObvOQhJ1fLxyR59NagZ4n+QXH/va3gVvYbmoi1JONXghcC7Bpt+s4fg
7KTPMAR0XWodzX5RPoe2ZhXbQ9KcBe6znkHZ12jXg44FLFu9c9uRc+xtzeyFX30Ev6fUROeMx098
i9Q0DqUgqnevwOC60A76Hp0VtD0YGJBMuniaBMnacc/DrEf6lMzhxGMGLx49WXyg6Zeuld8JPTkv
lRfOb3jqWHot6zWb4rsfowtl3C9WD6m8DsyrQ+3gDU6GgyD8lTRxFO5KqiZ7NkIjntMGRhsrH5wD
zzva/Ah0bMRw/xxqkGu03FQcH6JJE+PIgDutINB52n1gtyiHRFNACP9AYIiJbXyzHhbK0k3FKsrW
i6BnpRQplMmwRE1ZHTAcmB8Da1Jr8dUTtqU5vpV8lbnE7JchdiHahHL8nHPlnOw0CcPINx3/ON7A
mIA4Dm0kLgXMwsckB/6xPB9sEZ4jannmoLShlSW/mGQ5i71DfaAvfZZ2OnhjMkwgVcuUzmtyRTue
5L1L7/C8vcp74gmIdXvjBuAtCQ7rVcdghAwTCQyknPkeO2ZX3QuQNisXTl5+FTTA2jv1OPyBNJZ+
fLDHamUGU5oahqnAsbMOxk/TLvQ//IlVhDM/TvEeq/ViQDypCp8hrwrbkwdNMZ46vqw1ypKh7Moy
adDqAVilaMcwp1myiVxTOg6ZKAOjQ2Ce/fUMPQoRjlfzXgqZ/PsYpfkMaBK9yVjJczPIMMUFW+y4
c4Cv6bBA3Z64kx7oLqwpxptQzswqLj8K8Q0S3hPpPesgryydSXAXbJ61o2ePJT74e/uvbDFViem1
y7nGMhTxUzHJjukKVecjltJmdsKcRrMz+dhi29hqO44+6fU7WuZxqJ2dQCq0RWyVGrbsVEcCU5Zs
IehX8uQQWb59RyHg/U1v0i9KzWwsA7HxG8WE+qnbP2Q25VhmGhHbjhubgrjPn6w6AF3cBeaAPrs6
SuVF59nkUJ6UC1KaE7+Ks4dUbqge8rE/07NEYQHfMJzt8t3AAaRGzX92nNrIsmtqSEoMg5E3KyBK
xQCmP4jk7BUIMYDUDqv1vZtOaw+TEfNyo6DYpZK2qCBcXD5GRkiKS/+I6W9H9fzIR/g7L1ceGxvz
lHgZscA6YNh/wMIdUeAoaFKDiRmH7De0AHdaAGrr+fr0EH1xFfIY5WuIvXvfvLG9sjBDplPsXs94
2OeOerFgEr0jE+3qR7IR/A8ogcO3zE2C+pv5Ygd79t4iZwjgwftGCNY8JrxnXOKVdeTdpPhJTuqE
z4hpF/ueujqFOMsO2fTnwjMN/rPB/8ZoDKp0OyIwQgII6KjrbnqxuKEKeJ8vZ5JnZNUkwVGdp7nK
upMIUcY0076/u0FT6lZdUH6bgoF+4inu56HU7hsk76QbIa53b+FaBpbk+M3YDLw5P51ljllul3Bn
wwbxCNIqU1U00MdehTXpHtsQTaUKvejCRIVRQHTJiLetAMAyTO6wsul3hUQtNoq7Pf6r5TxKoHnY
SZmi113nDXToyX2xQ77/Oh6HgnU9HGtTm8MT4GQmr2j2TL09akvR3Mr+2YzdKUlsfobHPMPboW8Z
90dwIuKwzQ8T9/sbSF4LO5NB7+St+CGKBkF20K5xcfo3mkempM81+KItF8FflpWvb1lUc6oKY0N2
KVAInTW9vJQjtwPqa3373E5Ngbz7/zBDRBfNWViS31GGBaMr+GsBf4ocQRe/iIwmF4jABi45MVle
+2TgX9JsAuz6H83zWdhNPs1w/qJPqk+Spe5K9VPCO06hKOGKWz8056e6Qk4pZ2gY01T+vP/P3fsL
gKNwFS+vmtQAfDn45j+kwt6fs4vNa9iSBpd9bX8ojZAT6d6CnFEkWn/3HiqNlBTouKVkhc6Ivitt
MAgtvNTUsN7gDlbTVqc65Blf4w00ZyktEIa9WpEuATneBz73SPmCMUADsXhuGc/o5Cu0i1xCalMt
xfMgXoJO6O3t1JaZw8Bb4Ork+3b1jEkfmkwpo6DHSc0+FC9Xhj45sfwtr/PSROybcRwx8j7W+u9V
9XQTF2nJqAI2Y9WGZ82Z5OHCeglHogWnOaN1rXNyLikJs/slYHzeFAB3c5V50p4bZXCNSrLxTt44
OV5gVC0twtdC6+W6i5ECdU4SRz2lHvPO1o7rb7tL5LsetXf+6PmIbjasO45MqY9xNFNjwfUmpTYA
O9pOgUD0yqjJflEpEw3jXuB7ztf9O2DNqK0mNudUxlUpfNHDuKPnyYmHVl90H8p2bCxf1Fw0hx0g
t4xyiYY0yWfatp2UGPkqfY9Qr7JCO/GS9zdpK99rM3KA02wEWChqzbW5SgnecdaIoTpPu9QbmDAO
1JY72898O/VJNmBEVmJMt1rayOmYWbZ8KvJ5+abkqcq6Ltc6IXDhaGFteKvT0PE60PPWWgeDBs3j
HHltNAritEjqSMAyCR/Ctm6J8g24m91zTiHwAgWsyMpc6Vlp4e33QBJ/FfaQRhVjeq72ubTCR5wa
MUuAo3ndEMSH/7l3Rn1veqxeLPmiMJ5HYtqSzt0YMbuG73Th+jwxKpOY8Etmi3Xy95O8lUHDqqLe
nJM7z/PR93ypcj7Pw3HESDNiqT53DFpBeo68MPUhWoL5j2BH1NeVwK3bleTkM+VC/xE5jVbWKWwL
niRfomtOVdahG+5IeqYfjGGNfw+xJJWV23VsTUf+5n0Q8/sKwtyxCKeopdhu6uZYFSl9f7qUgHr4
2JSFTGpmg+nBc/2s2Uu2+1uQKkmVNNRBxjNlIibcLIZ0uRz3ggm4et5JvrkWl1hvadrc7u8w853c
44i/Ip8OA1LWCURKBq23ktcCMjwJLLhDq++8p/uePmnNQUv6riZhBE/8LdpPHgFjhD0e0SreSIxa
/igl7YPtOwHByQzXI3wNSg+b0Rzvmh535v6w4HCHSc0WM0usM7CBG7tww6Uz88JUVauaEodQXEyw
Tb2v4sK+Q3RaAnQ3githfg5y5uhQ36qFxA9slhJv7keq2Nv+zgfQMvboaPkSOWQvlC26mmQJjjRs
OYCgOZvCkDfXIZEQWFwAb2JZzq3gsRnUBXr5R4akV1XO/4Fwn/ubDNrPXuVsafAvVddHeNqh0I0I
+G/bvS5Nze+h8EetuZHekRSlYWRXUpy/JOWcmg/QFNPfxuH6MkHOCA7bAjbnmWdjIOPmLxQf1+hY
4mgp8mXZS4rKFqYIJyvTCoRbUAZz6x/1HXvhCtcHfwjnNLfVywff6iUS6b/CBXZEosIfuPSAyvB3
3fJw5fKnAwHqYgTplVYLfWVqQV6apLivoMyL/iKHXqPQ05zzw5AlakTX1ljYx49Y8UWdWwnoU9t8
hfrydhfkhOHkHD4cEmgMfy6m4nWBKk3hx7zWwK1z9Rsx3xNfG5lKmU3EgHNsy06riX6xiSwnyn38
geusUPlvWkgzbSpRIgm1d8RfziXXmC5uOign/4fapbHDW/8Dt9qubedIHS9uuc6QINFzEI3EnTWF
IaePqgTTjkuOyTymk75U0mt2v4SuuSMSfJX8RFGadmCxEWtO5BxAiV4+JGOPUAadPWKZc8ZXu7Nv
bSjBUSRq7wlFeKLwEd0Xr6mmj2IEmsRnMOAyiCzE9crcZa2vkGS7PBD+OLtkJoZbevO1xhhH8hkj
B8FjypITV5Vg7S61WesH4+0CJLHoXEF3yuqxbWAYM6VLg1b2YM4clZG7IcluH/fqO/1QkZW6IF9k
yPcg7HcI+5v0cBG2XjWpoyTDXRbxS5SnNOWLSRCAktVNl50JzAYRlIGpJXMYw2CJgqCu6jfL1A8j
E6fw1bnD8QQ8l8p/XE/1W+mTMN+qfnT/j85O3sXhLvS61KmRlyVEZcseOoT3qHN+n9YGWgmrH+hW
IJHmAkleFcirQN+mVa+M1T3wZGmHNWmFBDBq/U2qyi1BmOT6vMoBy/xl9oLjMqGF5ApuPFlHmIo6
p2gvBB4zDEDghqUcRiN7a8bGV12OHkYi1IHy3RuUc5HEZ+5X7mfjqsD6fv5EPgtZP+t8iuVpcemz
+HxZZfpBKItO9rLMFxqDXcIwr9UGrywa4Miv6g7l/Vbt9+O+hC7ZAmIISwWTpYl3t8cZFTLTtIWB
PeGe1818eOMYA5kw3Bjz2wKxYNy4UdFipl1Mt8IGXmgll3sJ2Vt+mroV3ZpwwS+wzSsnjPy/JpQ5
066gZD5S1GKDPKugvcJ87bPAu+l4ZbqpkO7GJ1/iu0117rSSyPeBeP19WzJfedis03PzQ8DYt/CW
hTI02nULz7I8vRuHyjwLc4GyqxzztN3axHioC5lWoezLozfvD/aZsYNkvVzTVunsXq6ofc00YNdm
Rov51zEA1Kb/ICvizZjP3y9i0dEWdR2y+akH7vGV+gjJdObzg+7vwSQFLFU7Ezj0mUh0zIhzKfsZ
FcY6O2S0zzVvv4fO/JtmQSLRv5kPr67zhia/PcbcRrDXDp5J06LDwtDt5mZdvkrNZc2uc/Aa77+L
AWseLyWa5yd6T9wtO0vtF5hR3eCVb8B06XbYWBFDZXkB3jCfogc5aSqIZl71P6SzwFiVgCblIzBc
dWe4GLGJ8beYGxogCh+2eXB+RzrHMY7FqlCL4+I0D8Osauxr9fniJwmyfV91ij0jMcTTOt57Gq/y
jfuqqdzTmnmMy6PyhvsQ9Qfv7uBZnGH+RBAvO0oEormGadK21OyA27HJ3YofO8eNJi9a7U8ulXGa
qh4uiwDQ4OYOmjymjXzRtA5lTI6eEUjMwjVgIWLOjMSKxGEQL9rOT9AC+WgKQAkYhAzstZF5iD8A
FtzWAfTk19L1QwM4TUSAxORJAsUfDgtxBynzBh0ufA/EVZeB+tOA87Jg0NDcOP1HbesIaEYpexQ2
1cwmYVoY9cEJx8sDV6WRWLOmze9vs1EjK+NxlGPhpLtRtV99ihdKpPTOzW+Qxo3JJgNEW25lnliO
f74W91B/q/1Fv4Fg4TJn1NDj7TkcxlAi2R86JHPFs32UKwFEvlQrx35BwmJqfX6/7ZyI3LShHzvE
wa/DKDP6ygCFuRhDp88oAGLT+LqoElWMjen3s51Zu9IZVVatH9XoLRYsvHXpAg6VbAQt+BP/EwyQ
iGH8Te7mWFI8DD8UL//WTZWldpmAlkmRUDK8cBqGmysetS8lk5r/5BGE1B2AgzzyUmkoJtKWQeJT
Jvd6fLb8euTE6e/g/07FTuNPvWh4Pju3W3NdHzwlpvD+7Y51AWsC+yBarlDgE8oZAJFk642Srv/J
FDXUD7b9V/WZwe3DUwBlI3EfpjlABrzdCziFvtAUylUEwnBVa7WCsAPVLx4GAM7oMIst7PStH2E/
SLwmDAFL0FqLknZlc8GN37qvp49PNrNr6kD825XQ7a9UkMPKDFa9dGVmY4GuwtvP0C76AaRIGSV2
04OpR4b4q2vLAoQHiWCr3cPgtpZaRIBYFYxXoxH83YWFldombvY7Ohvcv6f7pJu3ugQffIU8iRqV
aX0Dbpw7TtjHVOcnJ0bj90ZlnSUQoKb/GHWbBjdJDP5WnLJNOIgBSv5/Z2ELYX4CSbep0x8883PH
R94gOKmE8l3VSdAgfysOC+PJ4WQKLposDRTbehuwG5sQGN7W0sZbXZYEjU8GCu3MQO6E7vJzPsXL
bCErB2PPZDrOndJjoo28c128kQKdOw2cHYV6MbK5LRdsBk2NKyLPWHlPg6TPusMAVi8FqCcQe9MK
IhcV4D1PAgxWI8ZBF7zq0RkakWMQgP6gg1VredjEfbqFUuFG3y/agQcHMLHbVEOVXOS+fY5BKmGi
SBhoZSvq/u3+Ml2bzzGW35VwcNSoPpJRti/kfKz6E4BzVX34FF3j3hWN7eNJi6wCyUHqWRJKo7M5
fYQcM7kec4ZWWYEpx2g6un6y5iJCvw+X1V/3IpPTZ+x3ymnw3e5vwey0/0YZpkq7F5P/3lpAHAkX
9XxiGI6sWXTX80n5clz6AjQZvgGVxC0ok7134wTd2gxyyVbJ5ju1snYHZfeZLo9oSXHrvet6aVVB
lMo1czHkUQx87GCG1d8SBajP6IUEOatFsxX0vsGODgWiOJVOgRuIJg/Ua0P/ozXmmrhENjwSK8lw
T9SkIlzN0r22vW3JBP0igUUJMtLjZRpNSuajdryKXoIOloNk6G9fR1LIiogFKPt01W061OIRALSO
4gEP1DxdruQy06gxTOXnxJNpmOtQWn6a7dJkGXWAFiDZlbyAzrLZLhLzUhEOIDQwSjeoz1iruw8Y
OqTW71ZDQ+f9Q2kG2bImurpht3TGMWZiwMJmHs2b191UY7CsbSR0wgtG5aOfTELdzlIw4DrdhC4C
yvm9AKhg0jTXI/nGfgnLCXuV+peE9QPr+lfyr71CDjR97y4USrO4HQEJQDMhVHAK+TvGATpqGL8Z
brrijb9ShdG7Teg68LCi+3jgK/d+/zfJagqOqSa0sy70hkvcf7jXXFU62PyxuTQ1U64QHz9vWU/8
nviuLmtctUwHDa0yctAeNYR0TC11ZCAd72GX7fk+vteaL+S53TLEtkwO4c+3Q378AByK7cXQp0jK
rkUFcFFFFXcc4gMk9s8ZqmNxqrxPVQj3Z+LVZZBJMQs634+/gGZODnldF5A5QP342j1tEUC12hBA
md8GlnOUOSq1EQ0HFeb9kBR3ugrLuWJPvjnXWZo3kfgQYRI96Nu4L6JbQycDCYkaTzvoOJmx3SHf
77cR1T2taeaHBgggTjkz+daedrq0aPMrHfMRgirKZ8eZfw1+6DlBHePwSD2H010jPLQe/3NXKisP
c7X3fDzKfxT7jGBy+mYX/fZy5S/xIOI8sKldvSHBUE4LpQNROl+Z8P9J9WqxOSiXCnQ/04lv8Rpj
G3145HxWbocLJxmtwEbcDpyDAHu6WOhYHiTxt8+dKrFVKAKGsrU7JONrRrPfsSYc916ZzwRuUtFY
mgquoSipJPGJAQFKpp46vW/vgEau0priolsPBjoSMS4dgAl6PyiugMzTWgLbT2bS0PKgr76e4vRB
ujevG13hB4MSqx4fK/Bj7+zsbC3oCq1F1lxBfzejLGKZdSt8wMuAOaLUnLs6FOHgvMO231aDMPyv
yRDnDK1UE41fS5dpoEQEy3GsCSrC9atFnKP6EBx3UbmdMBaSuQAPm2IbTlQd1w3OaxypiMZSdAUp
Ags9/QeUxaTMmYuPhCd790YcLCRsLcFWGtcfoHRbyyrIEpYoeskTi2JQMkYARkSKlZ/tZIqOwPdI
G3pxY/Zy5LIIjKPG288UWdAj+h/rTbot8MoXi5cu6v7azDFmBnaihxA+u1aWCJfS35RUKAuKrK4F
FSYI2FaNN23vIzMY9y5zBGArNqrInBdB1JA8Pnpbj0VBC9zG+XNu8XtrIExTM1bB7kl6FbqR9PoT
JjqUWr2EHohDLaxjHSZsSgYR+a8ZlA1uHTUsXhSFeKOa2O7z9MNVUNkrT9ZDyQL5FhS+Y7w0cjix
6RiF6T9hVKQxi+P/PiWbdP8mMmpeNZu3JPEahGVulwxFz2GqIlearRmN55280BeanHoiLjwDDs4Y
nNnLBMBfijaFor0nXGuUvFDm7u86lOAePXVCG3Qg3pGzjb9znePbsvyiB2wcbb8syxa1lc/69sK8
CcgIwNzwapoZjyLOPjz4r51HsJpJfUpH9cghHV4IeP+4CuhtbqnBTsalO2bwc9qC+qqzpQT3qnTt
FVibKwMYo0eVgzb9bWYDtQ3z1GWE/MG7Ao6jxmY1UvDODr92N1kxeZQz0Tf9jSe3AwUxfSXvaR4j
fV1njli6gVbpntVdRBrlCFxRR1NBtzIRiP0W7gum46n89MRfl+SSWsXnFjHeS8MgL/6LxVj58weY
D5I7SVkR/Pv89bNpV5iWbxDTg23r+1jgc/7p3QRc7zWQME3m0RmnGbVSbxrd+4WDCZ5vRtYlXIXR
mYUn77Z1c7RxkyN00C52BEF7i+QNtJJVQoWBxKsO0RgI4ywT3EJNpEX0bDCDXT+jPNdCaw5FG29C
jB7Hd5KPiCErZa1fkd91sGiUR5cECKpTUDXWYuMJkpCT2eFeb8eYV7zRyYiO1XIOkbLdWF4FIVst
VPzlJOb9nwLnDNQAjmZQrdq1ayWuKbvuS9phwUEYYQ2GRmFNxGBbYhJvf+IExjCjrg8gBBTjkf2X
Oh4Wu8O9ug9D9KlLvrQ4xSyFwX0Bnb9eCOUO7t05H4id3OvvGKU/NS4JmeaUiUuemo54UlGQX5UN
CkLcvRAhLlmBzgz8d1GM1E9opAvgtZPRa/w9Ulg9nAyTiQMDChZyPyyDsI1SPqGb7UERYU+Daa9B
1LFau3XIEm69cwA6K4yeMJYRHeas87CW7bFtjpwFLTL4IWRjcihcFwNvH+JuBkXjr9G9H8ie6DEB
TX5eZAzjF6BipraLi+PcDfAQiZ/llpCOoxJ5JV3lB8kkOJ1XykCFJQ1Z6svBbQQkjz5NmNbDEdVG
Y3Pf2+RkfZtIcebcvzD6Dikho6gT0WnYpinK6wFCh+7buSKaXhjsLOGSXi6my1vW437HBtyc2/mY
HycwNJBM7w5rJsbgCt2Nm/DYFBdbE3JXIktUNYsCg7bJsZ+S8jb/VJ5CWt5Cmr8/lmPaRuXO/v2w
ZybDL2Ge7JWM0gRRM7aRoO7zt0Gh4iQCul30QQJ51cAClbbLWT3MyS4NpFQ2zYf4W8IBM11WsFrm
hPxVBjk/WrOWbEi1Z/dvdN1fHdHfBLUkIumeYK6w0UD1h8hMcfe7OF2HsJxYsgnN8atuUq2l9Of6
rg5v654OnQgwmEBVd/cLPgea2Ef192WOP2CWlB8rLUh26rw5HnWP4/TKAiz4HSAeOEcQJZvcT1LC
RpB1tK/p0eocvvNI036b4W1KsqS1Ydkx+PWgqcZuLaUPNin9iaxBSCQ01hpICBbun5AFSXqNehXr
JrfH4zY/swb6Om38+p+uK1Tu05YZI9TW4DwG6YsGR+27BKoEU0cEATxD+0yrPZSdBjZPAQHhmCqG
Oqa5mQgeLVRqEJ0qbmuIEKBVQgM34z5rEBUzbbzuWnWLZvRmfNXpxEmG8aFOAIB6opoqqZ/mqlc0
QEZrFEhVo5HoGbGc5tFaKfxkm02loh0zRr7bYLEokXjFn7pizZGbqlPCjRWywDZOa1riM8ETjhi5
TW0x+otLy3dum5ED8PKDJOR+eFapwoYo08623OlseniBzpxXf255+Tu5ho2rwbTsO5Abd1q57V3g
S00pEWDPStarno7moMgjREqEunjLrKu47mucgH/XaqLgciu/V9ovpLOrc6dJfc/aKVAxHWvq7oVj
1azAGU57G1N5BIDOxSIcdkqY7Gxjd7PEk/3AxBMoiBBOeSFoWQVyC80ErSm3sB5/4bvSQH2NyL8n
qc/uo/oevHOpflsxG6R2zLAjAJ7E0usbV3zGBUtp9VRnXK70OQ2PX3hqvP/GMzM9Kqwa5tc8U5gU
6hxDE9qAJfsKN2pxTmS6F1gOOqbaR714YWVxY+EcGQECLNTyjFZ2LgxfMNARHCVZYzMS607OJOuf
7OdCB1GEllEXrHqJ0ALADiaHBis8smog4Am3ETZ2+/5Y6vVBio06Oid6PGFpyOSi9jtGpVUEj/rR
ge2Ik7Ft+xjnjppue5oKi1AfAfqCwxG4R9Iwl/vr0PVUDg9uvZ+MTKBtxY0pLpbAtv3/zNr5to8D
dt3kYVHrODgngptR5oyiLZ6GFdMj+cuVK2XnS8flpGCHgigY+l8gLxVZVMAJCSZO794jRc+UC2QJ
JiRwdg/YDHcprSdozxGXgBj8ljX7ybyR24D/R3ol8FcTFbN6H2wMZarzg2UtGdmiLg1mqEHKFOjQ
51UHPIEIqgztiJ8o6N56HhqI32rwPHy8u6rcQoVuKYzHZmx5iklzRvsi0XIXiJo4gd2RoT0xvjHj
IdBTtfOLJmBVKG1v4o/lj1gzLpcQ+NPyNsOf/GHXXX0f1Tgt0u+RSYV7c3TEbtARICSiZ0vRAWmA
17olu4jk2YWxHtJi/ymbNwU03DTocxjF2i/OD5+jfmgkicKSO5bS/9nEIKWYTH5Mo9KZCK8KF1GY
oewPvTJrqgYXShLbqblHKCjynzkWh0RyD4lJb3uAJzfujLJ102IjD8ZQvFMtA/Cbo8uH4FoXLgSg
riajF7Oa9sbru7tgwuFSVuJoNNysltVoOAfEGjAssPUb2nthIVrl0FpYLF2QRc05/q5Hevp7o9AO
obnA0Y5ZWtm/4Hr8RnadeGc1gUjhAclWNhABl+FndDB4uaWpgzIZfIomqf0tu3fP0YC5sRVKnG7s
bPPuFlVL3VnzRC7WrKr8R46oLiEOxv4WmZq+uX+TFfr6yBEpuw/Um0rU5PM0EBFeWsAIgapdiUnn
k/xZCWHEP1jKMrgbPCRJ1WARI6nYVbRVaUlHraY53QnLOfX7Yyqr3ymLMggY5nyinMEjg7PdLV2L
ctXjTaxSityxAeBx44JgvxzpNICCVLXtMWpt5AYCaIsdIu9GbN5nN6Y9yY/FMop+xjY9NzCXEg4Q
9v/YbcVclSrdd0Fv1OG57dgr2qCYp6xVWQ94CwEmo4s6lIiwxPF6PUuJMUEETeE1fYFdeWPiEpJD
WIhLvLk8BLc6hzzsdnm+nml4mdQsKhOOCZPu5NnTzOAj+/ODgCWd6ZSJMQLu/kK+Jc6o89Bf1xmy
H9mLABvJzycNjfZ6CwiZDEYw7vzUOq2Zhg8BuveDcWumLgCzzNxJkBE7y5hAIy97IFwHDT0DA253
GMn86+wUFPuDRuW9493R0G1SU/BoNQcQccNyfsvQ6mxFTiRRFgf15kST0888VMph7WiF1/1W6d8X
k7EaJTQsng7E+rFueEiWMlC8hqIgFXf5MT3jSFjaCwsoW9R7VKwW2MlNWC1GdRIhsBByDlbMGPwE
QhbK0Xi8zIk+Foiwig8Du2X4Panq4qzxMKXOpv1aJvdBVEN0Pbn3BHB7Paf3JAePC1/90TQnk1PN
Z7UXrVHd7+xxKcul1y0Joyw2MrjfORHqD9z4ySEqSz6eGLKtLMMbiNciQ5fxjlZALQtNHNQcaQmA
AEbYK9ZRIe8ktiiH0Mv/iSDwtQm4KMkgPyJlRxl81gwTsKOBGLljMsThfSv0SdBzE7GLSSm8soUj
WEN1PEWlBEiBSF0JnA4KRoN+8kyq+xYS4v4WyJtRXqWcfUeK0x0R4Kq3qvtc/6EONsFFcQadGDVr
QAyfdhmmCIwNnbgywTWYE2uKIePf6ibNJt4vazuh4HpWPGlwN8viU/j6RzVu7GqY7nha1Z6vPDOf
MvQdJBQZtxWtJfQ6eYTLOt4xeCqL9MCgkiZ6HRVxMAA1Qdpf9XAt1Tx4f7ZwJPYYiz/E9v7ZGm5D
W7TV5CkMeuyT833/DzDJ8aFg38O/+q/jALPuH9NpudDu8oPMshuUh1dexn/FSCLBD0CQiYLgR9U4
i3arYoLqZL56PV4OcnQSfW1zKcnvy2BawhCea+JO2uzLS52qXeZu/YFqtlBzpacVZzb+V6EMLd3l
e2CMkK3KvO51A4pU0lB7RvWZ0tZwqskjUx2iNuK2gga91kL9c9YiQbAloe5mc3bw85fhDl7JcHYX
lXju4hHARmCdepkrHo8m2NRA0qRKXawDQqpjPyFA4O/VRUCYHcTRlqm+geuiry1z7ripKs9mOqt5
eCyaVx1iWOJ3K1Otk21qLyZ6CayUG6q/f05CVK6BQDRpIxC89IahRp1JP8+33V9DDG1xxc92M42r
WJUSyccqKTbn/AYGk/0MfjdIV/n2Fd1jamV+z6S0/c713bDMvgCfLk9UQvkpLNSYKLaspd3lGXAX
1fT/pQpwFG9lXBLucrYbyFKSDFPRJKjMBGNotTregpNOV/chf3iFjXBCMw/5E3Bulu3YsXbRUQU9
BlSrl/rbZiea//XeJm4zOtAFLDn9ltDQygsvB+OKmby7m0+cOeyfa4QKBiUNwzuumCtW91qEHQAb
dAEM0brAiE+ULI7K1i8Fu06oiOxQCXxWjX0r/LC9PhXaWvcP+fO9fxBoUVrpu1SOtsIv8H5LtSuQ
P58/ifajFX5+f7gFQDlJql/qzSfzP+D+PQQD7wh3gfGMCya7afR+t/wxvEPVkmlbOut0byu5zSZD
jVIgqQ++/kWHFbgW+i9WQ8tGrigNFzdoBB0ysI6xRuR4nTrWA80rI5XcZesD6hJ0TJ557L5LJp1c
EKKvfEAFLEBz8tVSCYT5UEtwQEIzSZQtLzUtKb6HbsxS/vI/1SlTYcFGnFzUsSXOL6hLTCUktQ8J
gfquo9EC3T1FHwbec5NQU+7aJwj7E4p0PV2KcruR4iqOQ4m93xxgocyIPbmkMRiJeq80+NmK5Lbh
B5zglZMj67+l5H4Tndy46k3B1O+kLWKayoyi/o/b20Z11GUTIxjQNwJJNPKaRBgg9UkmZK36dRTS
xbgo9QFyRbNHpRfxYGEeAooV0gi4bfSaAdzeTsnz4SXkE5YS7RlPI7jZxfHLIfVczIP+azqPawb5
Ov0iG+sT+JNxHhsI2innOnwBpDo/IGbIs4kN7ZK01Oa+D9k1kY8rYFuYKvEC6pAwEZdgZ+UYEoNf
noeSYz30/qVmW7ciBYYh4koazGVTeEChQm23GuWgeGGaff8Shwyc48wlaIG65MNoMojiT1narHlW
D9o+y4Waol77HfepVJbszM1rpmg7ovH9BavaN1xtUMVeKluZ++DCMq2Vw2ikFy3AKOAsVRIY83qk
Pjon+DFAM+WK7nJQ8V9zHSSiHyCP2Xmb2+FDTANIu9xpCVQsKCw9lJrDG3wle3F4a9wnc2mK+oag
g5SHbC8KQ+fGs70onBj9DADeaYNF/Zx6FrdTJOR8h/apRNogHwFaQbxx4w86O+16kIxR1/fys1n/
yZssc0mB/gw02IqxE6TyNKn/cwYpJ/9Fne+PJJcCwCgcsMDhP7ME8lAO6e1Ia9PcCmkTqkIXsKsz
tATo1sCD9jUcpIZwoYxB4RYr79nGiUw3VRelRyC6Q3ARmNgk3V5bYTiGMD0BtSDJj34KvhjJj7Jk
JtRRHg/JGe6DjRJrIlKFEkErHYJFYATC2l4zfciUOzjvbMbPboDCZkeonzlKi1GDd3Q0c1shyjc7
lGLqpFt3KSVPtvNmpgaeujNspjP2wB/01PTeMFzzL9/1b02grNco7nfOS8AkfdfSp79ndJUE75Gb
70EGFuVuVLu/F8VqvV+2i1qGAq7BLlap33Nv4qjRpcqCfUHqpvgdLHm2zjfV8QsrqNdIV9QGItYM
oFwga1klsOmXKRYHgEB/PRekBy4PdyprMlilQHPjsEJfzgTpa72QT65EN6cBPZBGsgsVKNIkVUe4
UThR5zXeDK6GvNyqUjU/15SvfhDsfORu95Cg6jTZrg2u7daFJbh4awAKdVZAcjFsH2zf9XkYd5+F
dc3nEn8925jVWxqxYszA3bTVUS5VA8lINlxlLY3MJGG5ktJiO6mTMXbXXSjKtuly/PVk06N91jXC
kmKSsr+ajPNRqtkrWNfqZ40hOA2WHf79fcjI0p8286ffUjJKVs3FY+3hQXYed26Gq+rU4jn3U0GL
VqCDNb4+cztbeey7kiCLxHQxl5X0MP3Qq7KT/utA1Laik7D64HUqCOn7axL0wMZ3T0sy0kgULX/6
gY+hBXGhYlbf6zgUxYrSaiggptV/57/Ul9c4m8uvx2KH80G6d9CWme1Yj5OXIlZpGsacVIyl6xCy
+mb+4sq2Z5kt17NOaRnrLoN+/oL2xRkG0xQOVVlMr46Hjf2Q+9Sy8h7UfM3uelKANQloUEeDwN8L
YcuszOfZhWsRn6V9Z7xalrYXgZCILwgT1lz3SEH73bv4FV2atMEJf+34KsM6sK461jI6JJ1nWtPS
jfMPQwZ5zl2YEsKXD8khj6eV9ElYD43YgjOWri7N2YUJhgtGSOuSjez4zeH2vcXudV1ZnQ0NVL7W
IjDbvqFNnEz5vrIhUsyWYfwC56lVM1vGdF8msjWpPSg9ixTn2KXFs0c93akQGzvDY5TQnGoFIhaI
5GuWbna0PXu8cWOo33FagKygpSz1nV8SONaitJqSwf5y3beysV4GGAVa7AYOOzbeXmHV3QBH9E7a
nDCq3chXwABRrXLexM6QyRHbMqJpbpd7uW0Y/DwLm/1U2XdD7FA3YQlZsizBkCfTI3IP8jT0xC4R
YBh5linjP+35FtZ7S1fZ0vkySXwvK+x+Dr0AviEYEq+OJ6BrDllBOip4V5Gv0qE+a0xEj3eiq8JH
24uwoFecESau2ZudCRN81gcTAapx5jHbi7kNAggF2+RGi9V+kASZDQc8gvDFEtRWsSE3i1Ox5ysi
Q70zWmXdrY8zDuW1dpy4jyaMeLUDj9Q5QEQrT/Nd2dWXIy1Vs9m8tzol4644PneB3CCN5Lr0g1vZ
aTrkzhN/SUxKXM8wB3G7TQnR77x6gNQZVddVXFn+rmzEtLx/7r6cFvZcqCNKvwr+kJhnNgfBdbQH
ApbpgRYleBXi1DhuTHfqeuBD4Zj17qxKZYNMR9xOGn5XFtf7sUluxxBO6WpGWOXfB6F312qEScCT
Jrnw5ph8tFL69NBUgtTIzUU7fJP43YPGDRBnHGX/1VZ0PjWFQU4BJ5kJa8qlYF3lsyeoZ+Jhm605
9r1Y8/7X+YKtg4dAaYfZu2IxlAdvRiRVskX4UWbQfWygVwNysdMGJuQhEYRhGxfQYc6vHT6DdEN/
sdIwOqj23ea1kzMRHWR0WpWTg+j0mfNxy1cTHmh83x1OorWOja2orSfdfqKQi779etw777uLkxiU
Or+VWBPzXikQhXrBiQ/ccu40jYi/FcIqp+dyQyChPo57tUjwVdIj/LdbySUlRZSBSOL9r9ckI9r9
ohPRe4RRBm83fIoa7m4PH01/7Jr41zzOrH+SbgAokpWuRhJbNcWlLktkAfH+7OJmktPCVBJ3MVoa
ZI+53uoTKvsDOrilJl/ce1uyvSw5WXD9A/srevGOTV1syAAzbCZ78lxHq2PEBDgcjEOhvnLvanFz
PtZWjvLGaDwMbgtKqdY6wLY7yfE2fvyPeC1qp8EGmZz1D7xly4UdEH5M5bIGjQJr94NCtRuecDl1
amecmLJCTLGpmmXe5pOn9MpW9/ISiqgmdV2+pbEnqV4JwDzl1YOpuMhNO6kCK7FYVG2W6o4Xsbtd
9T2FbmGwZ3pn5UyPzL2+czeLbmGJO4hhsy4stmR4hqu9VCEGqhAj0IwUOYhQrywjY9cYqTcOAxhd
B26hwiExoZL9vZmXahz4rrBoQWkHGmDY016T4vklV+lSmyrmKb563LKJadf7R8sf2eZjyUUwydgI
rGxXGwvjhUXtEih/qFC7OMv1TTV5726XNGdDF9GU70SZxG7MXd1N18RmWkgtFDnI1EoxbPjncA9S
RfWhdg/CVh0d0ljHU2i9ZzxRR+KxDoYjpRn3FCmj+rja3z55EUqA0ojKtx5FimGycrW8zHA7uvXS
0enWR81zmP4pFYcGNC8dQk4q+a+QmYd4dvXzPHEodI63qhDl2iVPxUEaD8Ju6gHU+++e3D3iVGIO
fiVtwzCRrRvju5QyER5IsAC1XGIjOuAFFyyJRtlN5AHzmClXwa6agtNTVpwYemaqFJ2AsNYgv2wM
GnpjM6ep71OxS0c8sbH8j7OYS0EOXp7SsJrPsKH4RskXbcZLkcp8V6iXCC6iY5BnPaC+KjOJWWcg
p7uqCuBe1a9vn58md9gWCfPByK2+Mm7HqMpMZRyn9bb1jT6RXEuBPZuBWmkaDpER2M2MXf2Dj7Ak
sRd3vRybfpxRBk/tpPzd7cv0DTfpzy4Bo1fOw6X8rtOfR7Zs/MQ3BFBjqF8f3gK/mmW/EoyLHt8N
U9oEGBLYRJClZuMkJ5/6jsKEW65C6EGuf44+31Aqfc5Sf6WHBTEvnDgo6O04eD6sw2XQa+lHrpld
M49DC2cNLl5FXOteyFVHdKKXse2vOyKDibhkNlGXuuZPSV7866I1K30e+oDaEg44jB7+0d0+PaMZ
NgjV2pCpypz9cCO8bEsUpJFquxqA9O2hGrrIhqOFehKeDqr/2sDycotpBfCciyfBVZg1YcsuCHQw
U2VybtqMcjEVSs6N7ieLT9Wl3wg/jq7pxtaB3zRvQI78Sn2sNcvEXqMEchvl0OdHF7D3gzldoKQG
Zgog5OGYr984KGJi52nthBxy9BU59weUzpUgg8DuOXrveVthpxEapy45uqhySSF3upZeJKD/nMhm
zozOh50qxGZmhORdJtpI6L4aRX8LzrhzfkKMheconVi5e2cQgL5O1l20F4Xs3gYqtnfRuEwTdfvG
1FZghTopJvXqLic2pO6oQvrvL2wSCyQBqZFYO+BpmofbqXFH72pQOMyTVTjjDqWdCErCRBzbUq8N
zX5DVnfm8bAkAgyIBxmgZD8d4odavo1AYsxZN7ZXyrOqRGpoMsCGl6cPuCtLJ5XxDmN8ZHYwYFga
jp993XrTqDdkQRy8vgQR5wwKSPuHjdamxUfz/wuCiN3VEmZyoqdrU4ZLYI/QshIsr9dY8gvBz15K
H0WaEFA8dt9lzarasu3PgLP4csx0T6K2D4ujJjWUAcvd1w+rS49jN44Ly5UCD6iC/r83DMDDCeWO
IbgS8QPw2uxpcnEJBnc2fnIPLabOkSG4/RfmikrsmjWTlIxgg1a3nccA7DoA/B/kAnWihwrg+wY8
Y0SYc1IsmJuNyGO8RPJ7Ql0Yqg05YLiR+qf6PZNJwJhEwZsmpzxfk283sXM4ciB7zEcs2oPiOq+u
5Ak2QURmfxUMfcnZEdcsr3XnpGKvGk2657P9keadHzKwAoHzb5IrPvQVfLthGe8GAb6GANG14G7E
BKW+Vvfe5hiXLB7eHvLrthlJ1+xzFfpOPxm4FiJahDvor7SuJINR1FDxLPz6g8VeLpJoaL/mA5yu
IGn0qesJPYgr5FwT3CeX4V95drMRq/lPkhApD3AWWgyvq7KHKEqSA3alfAQsKon8SSUJqRU30IZ1
ZU7A46jTpkuhqyg+rA73bxHqd3wshtukkljB0+WM9yWlosKqVDwvfWyiXd4W9/rUDaGTRpL7xFGA
T2K/ow+YwlQTyh/eUmnEVht7UwqXL4/ZmynmxB6KfMK+1T6HG/xZrj4y1slmRo2fTE8pecxKLsQE
CdEbUezQP3nRU4I8jI7yfC473U3q8teS40SZQBd7tan3C4Ebo6r1RRe3fw2PfOQn/pN4P41gLvWP
0433LPr7yYFBgldcluwMHq832B19wKMJJ1zEffNqxsjDgmatDNoHK60FspDQ0B7wburCndI6G1nj
Mb/saT/bvK04/zoc9l8exTNO8kW9whRv7h1OcOSthc9IFML7lLC8cWsphjRoLW6amMCO1QzcKbms
wSmMMheTK1Ju0amRmBJYZjAINND0NgODIgk8ulim+6+zd7jGprh3AadXJTkr3swjButzANw2JdAY
lFANXAjC6JZFjNPvjJHcqdrZn/y3sZdP+NF8MWdd6rA7ec1YeTM8LuhWdJhaVtkKFM7Wg76mP687
kUuVVDuCpunVpA5v2xXhqbmLh/zAgKZchzyCV508pt0VoN3Ci4lQaeuB/8/u/YkKsewxG5khWm6q
OA3mgCpOhBiKIUKr2M7zCkOrxtiF0cmkvuoZw+mvbLMAentRpxDLd0dcKQXtwvQve8wJvqsb4nGV
UUCffRqhHJZ30Ps9HCeW6qd1syQeeXM/s/FmztoFD2BQfsqFW4y1QRndlaRgcd3iyzT4WPhjMT/+
bbcVfwWP96GCl3XzX0IjDvd5zT29dji3zt37YjO4VjkIMkPV705X1tmGy0ORfIjQoTKTwQKNi73E
jFXhyhammQ300bW6YmyfrLbhIIRQ+1d1jN42U9EMSWGdiaSKHgAPeBUPIBzUDMNHjvDnQcmr+dup
vqOlvj219vEqmczocX7WJbucHNN+UNAaCGRYaONDmlmFbZ1DywyS2UYQ0+JBK4YF5u10cFot2+3R
5u43xE+t+b2UJCG9iEOwcrv2/gmDl36YU1u9ExQKkPBtaM5KXIpVfEVwmvwpDvLiRQm6LuV7edAa
4ZB9COaRkp/4vO1OvH2W5SItA7iH4LsJtXzW3co1z8IDlkxejihGUIr3pJNCtpavhinKT3akb5CN
D87H/uBmri9iEilCdpp19Wxc0D9fWVX98MVl5FYlQzptS7hBIgg5CgtUtC1wagJK2C3hv2DweKU+
2wtv3jgaKcoc9CxjojO7922wPEeAqNENTNFV8HMRPq92oDuQurGW1V+3FE+JdWpI8GXhwMIsO0tB
hLqxhGy0XbIcy8M8VGH4TG+e9A/kvMgawlsBkBq60OHMaub5UGCBk73na1ktklndrS+TuUisR0X6
LD6nAQTU/i4PbmsL0iQFYPVEt6pIjTLD4P6cgnX0cDncUppuL7kY1YlmEhLS1tM9VUG+pc6b6A+P
I+fAVjUK+7jEzUMdkL8XDolQxQDNz10bkDopiZbDyb8RIYpMRdo1g/OH1J4jwRNNdQXPgtwd+LtD
LTc1MI25FB+qG8QtwSuzHst3f87dTRAkjDFb8bhY1hoJ0nfntgIFjHwtlsszExqmkB8n21aq2WyR
f3HvquY5z3+nsGNAF8n0EeN34+/aWs1jqP4njDw97x6d+0nLp0AXUtA+RVPS3+Rk6H2XocI3B34t
/06oawn1eCjfiy+palokkOs3ReJ2c63MDOGCeNbd5ZFWTQ5Uex9TCHdUIPynzGaUjZvfy1AjygfK
IZtgP55cXs8eZXoxtdt9XVKxpMARGGQXRC1Y4EE1P/qFEc8mT2t++L3o5I3oSiBfWD0y+lfFygsL
mWMF2mefkG85Korx6pBufH0gXrF7vgEGJFnkUZMpfq1m4zGxqvRzXR7HnVcEttTsq/hvzQ7QbrY1
wwv805FyxWSuMq4JSpF9alyOtcz73FaRfqsGvNSxVwRG5URV/cBHdfkSTsGxxI1OsvS39ozRzODO
8blxkbGsVltR5q4zETyAV3Tdqv8dosTGi1VHu13OAnIJsUqh5ESM5UdHmqf4M/K1FjK40+1luEst
KViEJI9Vr0rQ2FYorZ/TLF47Y2MZIRpWXXsixizEaMUrE5EcpzJKFCOEoPSFvQ3w9DcrwApayYYB
wr0ClmEFD3KpG71dX6pZU/8gClx8ZZHHMlFhNtkJIh8NwE1jWGpfv5Bg6ix+sre2s5XAv+t3uEDH
8TI39pxPJzgvL0Azhzk+QzysibA4I8YmmZBVoYhwSHy+TZBVmSTvtihCcoZ6qJSx89/tlcmIOUbR
Q3/LLogxtNEEMuESc5WQ4olQh8TYCYhqU8cZ1vheCtgtZe7Csfi8DN4iWeoAot7CJzrQQEVZh5ef
HkX+E1P2FIc0NhE0LripIV4NQn4ZmF1tAmLBsgE49XWgWn4KnzgAxU3rS1Ew+cV7cVdlk1dnBbm2
Y5CxQKo7BOthuNETIHkqj1BjE446aSVIVZgquVIue4xUJFs6GF1uizEvm0PvCaffkfv0BU+GyvyO
tEwVpVSB7NrJeVPEkxorpRichMgQlulIlMqWH8Vh7RJz1Fll5n7lavfmDwjl7tyk0QzEWeJFOPtK
tm4vYfA6M8Yw4NVVys/Vueivl4cYpY1g/5lPPA0CD9RhGRI/WpAin7ycKWcpnID0amJs02/ctpr0
cQJyn64rw+0/3UAisF5s9dU0qps5CtaXFeBtkcO5rfAPUUx64IG8DdG1Q+1lMRdicFSOiIiaVDy/
wPWW/kgoKYeliEH/4UVPTiJcWhAUNNqLFVK75iyQQ9RrSulamAt8wsirpWyXkSG+JK3Kam8Oa2dk
5gyHzpxTd9LkN1SP72P4ICDX/cLsVdHtQTHf1s3wZ3i1MB2C5aZfnG048rk+JvaoOcHw+qhwvRFx
KYbajdyJZfhhHXHHDyhx9RgFLIJR2jnVVKtsGLbWAnqzKBG8uVnl3dU75UvjkxuaONGS48WdqRHy
xchIEI40w4iXhU63yLBfb23IvGeryZmkyLwY02ihBYIwpenWB2bJDMmhWS5y3qCN3qf0YQN6PB9F
YI5nZV2UkE8wQ6GpiOJqbh1H7zh5lbA8Rh4oiNNrqV9dBKKvfSffyU+1tHJmQZh3/vpQnPTmBd4R
WCkOY8cLZ2dKoiwP5EWc95iXyWCx6D1Lql87JNS9l+x/pjegxtbsUcrCZ9YZMp++4qUkbtEtktAt
zz+1eHWJjpJ60W6p05/iRPjPGh4951I5D7ykWj88DXrk2ZhbYbLsANA8SAAEy07Icu3qo9rPSaME
kJg6A0t9K5VyEKtBfenedL+2nVgDp3FuHajARUrOieOxBoFll89LWDX7Bqx5K+sl3/ss0l06KbLp
fNL8/f3PshQNdSIs20w38TzHaes7K7jHJ2UtrFC3i9qJANsxi3RIO31nGimpQgQU9pBKpNQ7e435
vRgtvH9ibOWknQHxG+/YRMf4cs/wjYyV0Psn4XTYdPBZJcs8gRnmZDAVKVVsSQXwmx5EuC78C5O3
YqvqNL5WkaxrbtfvatG9Ax6X9499AytAowazHMIcri+HL3eYHTyG+WF127lkiKVGYDyjQ5GZyBti
GIi+Ti1xVhYCh7m0C15/bja+8EwOt3B3QMgoZIBvdQmD9Nq2n/P9N7HBUvtf4et+valNCHPWuAkR
OLnJO3fFR43RJHKVZZ1RxT/wgNEGFr9u6001LngK8iYKWAc5boWVU6CjkqMc+wr81V44N1b6kKUs
Z8mkgzN5jYkcw8Tepc3yYQJfPOoYvb1c0t3NfD1UBr+KTZ+pvuLtU2AyB6O57ECdCl33GrFHYVKN
kx92WbWZ6WlS9Qjydxh0CjJmbgrD4GewnCVtuq5n7eGoYl59F9PT4iqM8BKUWdSrxH/GZ4OkoT/p
OWu+NqqzOhK5+081GSMsOpsbOyOeuVwQWp0RlTito3DSzoKj9hThJ0MiNZMsy5Hj+bVi5tQ30i0L
ianSdZaDqFIn0RnmfFpcyccREjs7f4+GNFhs8qMlC1lxukx+oHGzYS3B0dJgKSElioDnj4hfS5cl
768oBXNSxdfUZKznOOwHvnSio+bKXY/2Xw38MaRVKaYBuz2adNZ4k+y27qRHxy3iT+VtH5XB/G1h
OGgkAZmi+OpbubcDFqyZm1iXy9yVCUj14NfhZOS8WT65hpG/mytom8gQyGlLamTMh7c3r+7IRAQ6
rYb/gmzwjpOCw9+6z7tDogg5R/EKhDOdyKwlPeqS6H8Bb7u6ptTS6tYdUX7uG4eIEzjDK3BdvWvr
M/yVC6kprALbPLrT0DMFBcZFOwttpsj4TIzn73xjje1Pm1LYOF1+FArdoTLQH6y1w8Ykd45lKkHZ
UbdJT2BqRzu3lJHgXwyNm58CRdW6l+Wei5SPuaVpkbChgBluBL96NoGa5HaRzt5a3s9AWs38mB9z
g348OVhH2Kl1V0GtbjRBk8mdZWVPidhB9C3WxwPBFMg1kJBh2qSwLKJ9jEiTrzi38lvIngjzk6HF
dgqwCNhGJdEZ1lDWq43bViMlVaA4l5gH0IFjW9dD2uOMuidRoAhaSc4j7m9XUueMAprdAMc47B9Z
E8y5sRy7VcwCOuy6suLPeZnX1rJCzCiLthmrMZEJZPcS0FkbS75NJiIq4tWfKIrlDGgUg0nt5yS5
iobgGHZVnjUnkCBvJP2eEBHIb+zmjeg1fQAjGGaxyTe1ngCOdPjeQ2MUliICWGO1Kipm80thw+D9
P2chy5htiTWCd6GPAwV2cr+9r7LeL4qnCidEaII3gDt8yJ2tgo6IWd/M0VEpiNCan+1pqRKgE3/r
GPPhgW9VIzhjI97QYDysHHRW5S0JuEO6FlOdZHiKMVa2wuOdjqmULtCGXJWK4NeDQkCCcJg84g6m
7SNXlzqxl3aEeQSNYU+YLfTxWlQusu6MlrsF4TMBHN+MjWAao6ZtxG874gi1l/ohXGyk1fVrdqPa
xSn7HWCrklRdUDXTx4pE7PzbQCE2b9uJR2Evxio/5b6+Oo6kqncEL+cXHDO/dO45rjk3/9nGJt4I
5WDOauhNgXJeOAqnyqD87pZWWRdRl5FmFjsuUADJ+4pYQGged/Y9UQm6IRLfNMnIR9RyR9weywuv
ovL3HZsDw16goOOJgeCUl3/PHORIMW8rtdQgo9Ls0K5itz/MVWoSacSe00BA6031TuUr2d4ENpXP
JqU4WV3hGV3cesMm/1qSHkFGtQhky2xVtWxUbPgr9yq8vxqvmUSXpBHJljSpAYXKK9vTk82+zlYB
ALdrlNdLwcaDRYFpz1xbEnK/GaFXYMf0pnzP0K6BTcfduzuGUjdwbAB/GqhPu6FPuKZOvBlQSC4l
6fWMUrRMK/Lqlq/TEqCuIQewcGuiakjIpYoszArlMN2dpQjNmgNBpcB5oQT8dK/12ni9i7ReBxV3
oFMhfKoCyMa3Kq6Vi4e0ygVsiY1W7gnO9lzIKe2MclzrAoR0bw9AghPeaERZbuSufE0UlH3BsNpH
DCQMrV6A3R7GuzWv0giv5KgThb7SdOM2kCsP/aAdLFXggsue2k0Gzy/a50qBNhFR1Q60d6CN7jYm
afamhkf7hZwHAkTe5oQbMhGnpmvsCMisTJAtBBKgKGCIbT9knQ0cR/EZhhk1U/8qpXD0XJZCjFda
dCYd8IeZ/veEGV3H3WIc5fXcQM/BLpu90T6iUPP44l2+5LfQDVndVyAQNmr8kuriOvKq4BAL9zND
E8yQxrQrLhWLzytbK0Jw0hoKf9wghd2yYhk3YR75s4xKvRh4/DTfUa1XlAuixK8BLPMx0iARHo//
w7e3dYru2/XuqA1kHQQ/jzDjDFjmQ54YPoCCxkcGzJBK6+G1Pa4sUep4O6J5fLUxkM2B3+bZgWeS
+XyAs823Blnu9iHbqom7ErhfLZdrZagCRtnf0MpIB5MYu4vJXPRS9Hmyk1djvOFXnjSTq14J8nSu
Ajnu8ANfhnjuCnMLejVYNbRA+70TgkKNLnaq8HhVu44/XtxBZQyUVYYQ6y/CGoLmg7d6bxwNbTfi
wae0McZ3Q1bwu+L2NHwAwGrwNv/H1O5oFIGajqqc9sODbE8GaGr9yAIZrzdBT3oHowgnLjWeEj3V
ck9gM2xdEW4/dXk30K2n6LyKXQCy34LMcSruipxJUjUlaLvurHIs4jvMx0Gk9v70nyodq83I2ZFb
+a3NfU9E/vpL7V/Z5uj+0IioMHGTy0+TpaeJpGpLN5u+CQncrSNY5pW8OS1Wecouw0zKPjq6Acti
irFXYH/pWcJTYmJ9TbJwhbDK3LAVUourESQWWA+qvhXYcOTa6pBH+fkNDFDzrNOo64Ake5d4K7Vo
9vKcDe37dzeM5zKOETbWLJaIlotWEUQGzD2Tvk3jRwoCaZ6TEMI/dP9eVDFejTfI6eN/9ole9iAO
gjaldgc3wTFbJBIfi20ft41y0Wqci90BsjS7AujBbweLwh7DAwYZfyBZbanVCMr+EeMBxQh4yfk2
mXFDN+lVkQrfn+UsMo/NKxvSJ3mNtsWkscqLeAHGbrlXBoRnBRrkr5p8boqR5oreaI69YmyVpip6
ll7kbPlL1bjwIN4zXEyLBZRh9gFwMjUJOTpsqB6eLHrGKncCJsW7e92KSft2KXbyaOQ7klJiiiqt
qdQJ4ezbas5mPOlGBy68n4nJHErtOj4Fje+gYGUnJcT1EXU3ayij4QWToPVQ3agOpSUh3k58mlad
cVWpH6zkspOvagML0y18eQhVIZ9eTMv6UYw2o+Ps7lHmZFxkjO3hgyh1xQGnvjFI1KQkgkK6D0L6
xiBxH3DwuiCPRznqkkyBjgHivUckP3X1aIZKgFmgpDM+rwk3usCwtvYpqw8oYIdonCGKh4PGHagL
cqIsM2vkS7UeNqwmZFf4/AdSpQ7+uwb8zwtghWLac0a9WU7h3H+B42mIy1yzMs4q30+xJFTFnstK
I9WBPmsFC7x/3ISSfS49+yUeGnlVm5bue0Ui+XgSVsT6vi2yzJ0BNjZTZVZ7spwQkf/rR3gdVme9
TfYxU5oPCKq3GZWgL2zxbZQIXpmZ/7XO6zXbDF/sefaXFjdlG1/VGYTGPe18/hzBLFY/5HKDIAFH
gLw5UQ6h9ekncUEyhx/ADwFQWk21OkmLwwAiq165GO5ZrQ8sXGFYB0XbdE9ke9YY+uJPrENSfVU9
lN+D4whF3q9P8C5BfiMayZam+PT9NmCqUj2GU76gVyZHTBZS+T+40HadqNrZupz8EIgAGfnOsBpI
iNAtJN1YEBhLz40/AZTAjviDFL3jPaE4cip+qxgBLRsL5oR24OFpjl1FKO55mY1MdXkDQPUyQ1M0
hZnphV7QqVSROxv6A3TpPGZxwoc1YqWmT+sGJcV6fi70+/SJ+BOxQikTnJb3j3oLqNC1+qUQxEcR
2PDkslrzLvhxd+HOOkTvN1m4w2Pbj+xfloWvYN0rjtsCBjSj8vmZvdxVC51WBPjBy6G7kY0xA+Mk
uHzW4J+PzW3PZg0/5Z6kUH6NQtY8wLUvpB/+OUKgpxtcxywi4BjQ/4eA7nwhCXNCeACPo3BcjOdQ
Ldynaq2K6anTAj11y6k5BNZspLCXRfI0eOhvVODq8Cd6q5FgVgeRGUXE9X7/X/UbgPTjlFH3z28f
44sFFlH9CxD5mmHheMz2M/aTWjhVp6OPj4sA1eDIivq1uveDUlW0qZUPEyfYzNfTEJyVgsv/ull4
gF5nGq3J/A3p/8Xto3zhIxO+KU93P+QYvZEpIe5WElD+oRNDnbqY2RaM0gsdI11a6YEI9gn0AEVm
pzP9gVSYEPfbw7QQYE3mWe0TLveMQYdDQ752alYO9K3ctlhdSk6kJ4ZtEngy32TKSEjk3G7w38AG
whmYjoODLMg6YwiWaC87Bj5t+VwQPrFYSfu6wiam6GOePcvO4fw7yGqDPeeuWDsOB8AwuWZdGkxY
U63mcP6DxGzh7Ik35DLg57+E1v1/19/rztFyLZxVPPtVT3hFmSFLRhlv4BzR0Gpk0rznjZu7C4tt
Ib2I5FWFTrcf0NwCnZVwNjac1Z+zqBrIrDJKIgNiIDfsLdrQmOsW3fYpA75rfkf6XRr/oyHxxCye
Hjg8vaGgixBNe+0S+VKc/jo3wzvbSovmqEVCWnm4K1X50RurnguHdpPXtAut5XbrrNKPLP+bHEkp
SAcyAfnunfPwtvPJCfPmEekhb5eVM5KSTsgrnF33dyIM5jERTG87RdqsgR0HyRgSHB5aeVbrTcVf
5/U+M1c/gRuPQzQc5yMmwp8/9LtJXWH9Fio58RTHWXO/0p0CoBsPpHys19yTtb7L4WDwMmwCHviu
1ACnBv0WxhvG1SZSriF/FYses1Md5W+1ez/oGD9llP3gkjmT/SBQacX6sd/WzY8x/d58zysFJ4EF
lLXhp0nKQvw1umwNybsuls/fY02FqdlyV9jnKwmJUVyCtZFpy2u3CAEz/X7mKb6xTcIekeYpzOBR
tG+3o8DN6YshBvWagi9mQiUd9c9kT25CmDWQkOzMKFOPS8v0Jqxvz2VbnGLriHgqgvZJnDATj+M/
JuVPzOLqD7MqmO1h1Ew38dYHQrk6okqQxQtpmglmg5jJxSlRsNfQWkj/eBJDQfV3spdgnbOMswXe
ExgewTj+iVRkluFLYek4nM+RQYNjxJsTQmNpP3yaYsrQTpTShyjaEZ/GH8MuyjEoI/YNui2erhHP
2C3sg7m9d4QECOHwnvlhLTyBdNhIjTn9hKzZA8zId5kvp2o4FedvhgP4d80FERQF7Q+rhGpTRQ3j
8cb9VN2twXQITVSQBGyg/1+Y2LFNeJUMcuoIhHXYt7n/6IqC3Qt0xWH6hQ3KTlvLD/XpnLqd1nvi
V2sSJsVjrQEWcuUg1HSOHif7nI3LrQxyGEIVNT0ko1hclVJQ8NA5O3CMNmDjFvjs+EhXm7IzsoT+
VXA5p0iRXQqmI+EH+Gx9ME7UKkzfwwl2gkA8tDflOibAdUcf3z2IfzQsZxBPlkrmOA0pWAfPeldg
Cw6fUccdVIGp3lDFKD52yk6wvKeMW9yxHHp6jjdJauga6s0wGK4vTi9vqhcZ2RRATqtvxTCZ3L7O
YS9VlIprGoDW+E42/oQDTbwO3yFMXRgHDB0zx9GKZ5kBQxbMQ1Qu9KbUevune1nGeQjhchESYy7P
VvJ2sXsVUo8EMW/8nbDV3OsysLYm5xR77mEaxL0IthnK31kKDrQAdhh3l89Dhsm5Q80PTzgxm+2D
TpIdh35xmUcPddDU4fMZ/c7eSuMh8itZqK4wtHWfOy+Vkj9jLsLGW0vBP11V1XFjAC0sSXa0o2Jt
hOJFqTkjzDpidysyNVEfvwvj/9c4KcsL0bUa3ZZf9uAqDI10JaO7pGtTMDyd81oXD8I+5NSz4AOB
nUTcGe/MmPWBLJuneNd62NVuoUdFANvoXkHh1ANbAx2MugNfessHwq6ZyklT4+K7m2Wg2Xj9+4Yv
uRPrhGS7cdNdNWFL5CMnCM6G/0QnJZDOBVy2bATUB50bg4ca58JnIdQm13LSK57hMz2kvbk6E8FW
sNUojZ+n0jnRCJMGH1Dzx7p3obWM8gdPnev8g41KwdUULt8cCvW9B3wqC4LmcX+IZvnVlmYZ12Fe
9mldftB0InLaZ/j8gmv6nDcbqxUi5mEUBQ52oL97uIppeop+KNiw/cXK2yHlJxr+bfX/YZ6SMZbM
lMJb0QtHuHV8bsLpNIlInngmk/xLIt/G07zM9uv525Gk2CVW7So3idxbZE/ubOznEXfcHCkQj8eE
T1x6+X1uGPjHBMSVrASTJ2smRWs/IaUVvAuNwqx05OJl7Oqdfiz9Z2yUiCUaIzdXCm5jYt1TC1AQ
+dY7jVyYxrQZwxUPbUD+BS1RE3u+WoPW27IBz8CPXofJ/PihOUshNDpre80eIM43nXssJ8NmK9ji
sQCrxnZa9okIT8hzre6giy2d5Qb1eBhKk9rqc4xh5T/fMjHjA6Pt1uF71f67ltcW/mfWOPyhBIMb
2bFp6vF3w2/IVC1F/S2RtgLXOUhulDYjmYGoCN9tIPf1p1FUJXE8R3/4EA23MqIorbB5UvAEUsui
qNsZvYGg0WBqmoHYTwp8Z4LgLCnbiPIVyNYmAjPjwCBetUmPkEthhLwR7+liD/ooLgj2FajPFHr8
Z7v8EoVEApuW3w8vnJfJlZB/XPhlzbjKt6CkW8efH4xSCO7BYf8DjspwvQ5jJHBkjP6dZ5FGRtom
oONBoHzrFKV/GN5MJeKUFLbc5AYUXm9G5r4TNCrzPpoOZmVHCfNnrDdlMjanTn8JPdMBWMvNno5V
SSMekgYdVYeDzdG3yXkT8UCo2BwSgJfZvsHDazTSTmoWOj/WjeRMsNQcDQIJ/abVSp7Bp5rNsdBD
ocHOJxI7hAWWAOe5atBrKBxPY2agQyhC4xN5S/hw60Erg2RPD4kCGwLWVez3UDin1KqN6V94w7Tc
9CiBq20Bme1UP0eKZhMfgmFNEL3CpcVR9WSjvu4Nww5mN2bBc7uzSHUA7MNTphXvTamqvtjU7S4n
Rf6CZV0UHDzE7x/CQnAD5bRR2EKGs6hUwxX1Et/LCTwSwhuFk16fsnn5fX3IoJAsWRfnNw99dsko
m9TukNEqYVY1yv2uuo7Dr5t+fWlIND0lyO31ayNM/FzruVevuYpZeUIvrtWEUmdhZ8sP1ldS2eMf
/AuCCGb/3H9XbLsMLroOOXZfiKNG2Y40m2VtZxQmUzwi5NVvolL2J/FxtCPdSU8w8AMdxIdX/QEC
e0VXMS9QOnPpGDTDjgi7LVfiXKaBRwLw06DV0Bc6zyqLjg9jSTFIQdIQ3Ln8Xy9ybcBHxT3DAlNG
xKniXmzvvPUJgI8k6M4g+iRDWPkrgzPgk7BY1wkfZ3DwsABP6Ysc4xE6qROdBgghx2Zd5VUXVx7e
ItpyuHQtly4ssI/Xpifoln0JM3RqZyuol8eM96lgBaBz4ATFTOvBSpCqMF7pnEaiCRY/R6Mdl0sH
PPEoGWbtjkf1hckm3HNvVCCIhHAOoysxIiOQGVYAxrKxdjGmWqUCQJk5uGwsCNrSOs0uZDn+foqM
gcPaJLHg1a0Q9dgT1f15fiQyMxKqnS3gQykpQRhPD+Mqahjk5Z5q/yKfWZpXQatOObkWGhO0ea5Z
Z5GWa1PFOWzyJX7OsN13Ix8FiLGDDwGiTfOVUrXSqxAnqJEU8zfekOUsJWu7UGCMf4ZNgFHOwEjL
rOVFEwf0y8kplKUUcGj15Fh+S3nGSodrpVlQ71ftS2FJGKSLLVO9D4X3PSgSMp9EeoVPhAKRNETX
Qa+7GVeeUf1nllOc4yBooSb7bKPPCZIpCkE+P0KUTsIdedx+U0j/pTexSYzjcxNZUhtWbBJfRrnn
UlAHGxaek98nKCJwgA6yboXgZg2HMDgHMl384DLbuMPsduLSD9usrBOxmjpPJsG6qIryLHqS35Ie
B0ca3YxbsPfUvdc6bgQPcPf+tA2GMuGig1hdixEPX0qYXAO9ZdOhhOaJasXYGO7LA1NyaGoUwt+V
Q6IA6gqW0wFFMSozEqpBRnAVd9Z78NdtlCVIrOKWTmDOXGQtygaJH1+pUFJsMyOy1xJspkyqw/kX
/7LbSDuRPV1IZ4MTJwTv7hiJtYnPvcGHYZ3VTwIKL1qIm0kIEJYooe4OcRSGYYq8zqrI7riAsMfn
N5GLWS2VfesCp6CoGf2PX3BoBaHWrF5qILkoAiCZv2Fc5ub2/QJPbTWtudDrzDtl73jt1f8kn006
go9PHm6FYxRSFM+3JukwXUWAsarllVV7NlHKc+CPZVmjwX2p/y8tRg6kIk1DHQ1KnYFhq2yhoHOb
kEpZ7z+Fqx8u8eiAUDmgJo3oZckKRi8tNgmnTmw1b40kLj8ds3kzB/SUj7T1TTJv6D7BSzoLbZYx
a1a5lnAvSk0ymORVUk0omNtSdwFn8GscKUZnv5hrmngyRcmQJCLBad2cnziop/7Xd9Yt0lss8jsI
oP1c3p0Z43nklD1ADVhqLX8eM8rUvTB/NWCV+x6xQ5bs+2qxzisgCzuWc280fT2wm8G3O1MKpX5A
bzNzSf4nMQqbjWESNG3yzBQshkTigFrW7VZnQJkGoo01VXJOwPm3BvvXdFn7bqZsCrdQbHvki14e
dbhWDXNnA22tWRA0D+kZuQTtehRzchcXFl+UU2Wvbl+Vf4RMWXsgcyPqQlg8lA4iS4WA1C1TqEZt
Y9ix7+EDBWtm+Sv6XFaEPcH/DMrfhQpa4caJCasMSRgNznyNEC5sAQlsvOMGRPftHe6oY2n7yG63
8PeLykbhmTFnFUJAfn0Nmes83b3+VMAVpKTrWPQrAsQjO5LzfOcR5iMmLVJpz6J+rTIliM103/DW
w9DVx2RzCcb1ZQRu2+bucbs3sdgmIwvQP5JzXbntUWX7+euR6cyCLanIfKm84ZYiBrE9x9Idt7Tl
wSKB2ZUPvvG01ArPOBAt3dkw6Ez6Ldu81WjQ8SDApgACY877PX6ZYnOgnq4Bnd1CUeTwQwMLrHaS
RRxsj3zReZ4lis1ou4JOaAZBpqvr6d4c8s44Afu2NyhnQxu+wVuiId0KLqK5gDK+DIo9SZnDswjF
rQgLvpT59zucMSrDllFlck2fhnBZEOU5SJT21OGTbh9EcMBF2atjCEUMtxd+UixveE45lvyCazh9
FgmwJ6/15dWcQ8j9ho3rd/VpC90Klm1JSTbUDqx2uRG/Yzt62M1RLKruFxtxUS1AoWAY+aI1yT9k
cFdTv6ZyVrpJslTH3FyVH8zawGbuhCWgPpRGZag9Ef5VroGoF/EFqTUhFQenvbLBSlSHSCVWhKJL
L/GjkExf/7+dK7FEuPRPnD8NvpywS5d4D2v1zDH1ygcNaWtRRLIWibNYuLcrPlwnJr1uf5G2I6oU
CgOBI+dU5r4gShqWxc8RPc7aQWbWFRFnK5YgsHO6y4TSVSD2dSiLOHuwGeYnPv/yYZuLZ7CNtig7
xa3IxQb2DWnHybpogS/VJ4zBmq4a4qzYPMISKo3gMgQ4bhFaWTMaYRyA0UoBsfi5wJD9NkoqNLdR
b1oDZap4xrEMP/FVr/OTaD5UCXfbBAfrDi7RS00o5Ru7b1QOD682Owa5/5WxLjUXkRxMvBL/lcq6
+1rt/D8nUG4Y4PvOtslEM4Fu65mUD9sDvr4fxdpE5zRwQvXURzmDv7EqQmjyEsy1oulWyLVuY5iP
6Tkw5QnOqd1EOBTlWHNxfdcp/21j6CBArkdC6B+Wf6n9SMQvXMlmro1joZLK3kphvbUH0/wVRKw7
YtZD/AlBTSyKxTBYvFHKO7Q1jwcyDDmIeYiOSiv7jsUfOJbpAF2e4hi4+mlJoSU2H3EZSpHMgy6V
v8Th3UWxzMdXDk67tUQhRlVqW0Gde0i/w8La59ICUcn874cSZavvkPm/DX08DaRx/y/KxFXSfdIE
IpUjIwl8lf4GwKq3kN/HtRQv5QGgg5X85hpHDw23BCGEXiu7DDxha42TmgZrvpJHIMDxQxJT7p6J
3PqWMmJAq1ZfwqeKx5QI4AYfTdpoPJpBDROi+TIbmWj7zGPBU8RfjhHFwNnqnZHHYYXYpGZhfnBe
JiKJXuJ1tv/pGeqq9uk9mjrqTcduLJZLnStoq+f6aYN8UqwEupbogAKmHM4Pte8bzl3W71BnhwVJ
Iq8XXFszgzraYarv8hGHUXUGN4YM80stAAUxKcbWq2khoTfnnBBPJdVKzSywgeE/0+DkHrsdECdE
Hm3dKW+bRVQb00qqSKOXzmHhOU9TU8z1URSB6mEH/nuV6dnrOMJl8aeAzPuDOzuIHKgFcDIF8oMG
abESmIBoa1cC0DAExSwvM2D4q+PtCRtRrmDYN7ABdM5xPsYLDzThSXZOSVLBlzG7mpHW4fcVHNRD
scDnrMkFs10ojKGSQ60dUn7VQJUaon4aXNRdgxndvpDvjEpwJaEZLU/27cvV/Rj7U43R1YRzPpfE
Qi54jN2g7NImrTiBm5YaXu9Qpj4bsKT1jkdniScGbISOwTQ5Mo3GVlJaAuHGwjwhVZC5338ZRkVp
kRgTZZMuGtxLuwHTkMFyBRT8rRLpcTrDdjtE2VC07z3u/olnx8CH0JG4WyLwf+9u/EnmZ+yVQbXa
4corPadBocvINKWOeigE1ncPHWPsMXJ+eKw/HaJIFpmQVtFi3FqGCf/HmgrfCU8srGRwXnbYbCkb
6Y/rEKS3VgrWf9py5FfT3Nf8vA2JHURp8/hyoZLjuP8/0oc0K0FqCLfQyO9lr/ndsX+NdC0mZXeO
N9m1pwpsC0ky4hmV4cg0w/ZR+k+DGDCrL5dCZ3tIQAUsIJh4efwtLBayX3sMCLla8EQPAI/uT8+a
S0mbWkrZq0ICGEQ3AeYs2shv1nrmYBc9HKpUe5TtOcSrdHxqOhHUF1ln4RuHr9J7v0/Ijrt10DW6
4QHsfT+oiyF7OhJrUPCUvFLSp/9GIMi5lHm0uXfk/8VSVvuNLS5ndfiHZhQsnDBQLAybKl+7pgbD
sD5b9Rlr3+FRTSV5VCTSZ8AlZsWWHwUWepYxoq+xAxYB8ejRq1hii/9zaTh3iYx87RdackbwsjV/
c5S+dU2fYxYYSd0j/DuCZzLDYGp6mGtzO4ms0mKYDSWGPnrNvwJQhMc1Lec6UF61TJo8wl/fHMYF
UJtH+niQfxGgsc9lKY2T49lm5TruebiCC1XakLGGJFYA8/BBW0In/8XWlbT2mjKCOSnaeWcb9yi8
so4nX/XlnmveKpG6X2D/BQqLgoYYgfvXbnWZiOekjXDveWykOajEqY1EmTixMcstWbB+cIpDDmh3
hmAniD8pFjeOrNsG0+giKwIqlpwnVYugJ5pFMnkAyuRTuytB8j5j3fmDPsnzNR6tbg56fsgdDdiD
SNCeArlxme+KzB9sjq9QFxuRCvAXyABBdi/O6Fg0bAxXL5IBre4MW9A4XvpVKPd3pvD9TWWFh+Gv
uJnoXq+CMKIrj6qhfSYCD48bCQSS9Ix5OP14oIX+CFN0Lixz/Gqo9FgPo7Zl+8Abgrbk25C3m0YG
fMJ0L0GMpvuaa/W5rbNl+PrEyZCBKnW292faW5xmk6auPpJvKvqGSGajmmDHBN0WvDahMBBoUD9q
BAxKMkPilCFxH+rGebi5Xk328+/m1+HdCj+49Mu1glUMM+W+vEJKrux/JEl/zB9alg8EcAGp7CVw
bS5dAuwalvI7aVL1mvaKquXVhc9b4i/0E6CRXf+OJ3kfgftOsZmt6Lyk42j2lMiNQS2dcztmlgYf
6hUEf795f8at836L8/q/2SJz0IU60IQJSyCVcIR5VUJnssRYMHDgA3ERn+ihhUdKDcdDrIDHc8XC
T5aoRvaag8c5AOa8zp0Jx2kmo76wLWjUUPm2g2MlSpbokcRbME6yV++8qDdJ06GYpu/gjIs62fAf
DA/S3UfQkcpISEnmfzkCWufDeJK25ZRJzPvebaxWl5SzfQn5gzJ5WmAlrpqz+FiorJEEItcK6Yj+
rAtSRyzj3chJ+JstQBFn9JQMpHEpuo3qos4dKJvOiZZU0IoYoqEP8etEoOi+pAlYos/c5oKYxeJm
NAjr+yovFUywYsSirZwplf96reylLnwU6kdmfez0Pc4HAw2Q4x3+DIy8qQ9D9207QjfpfziejGlm
bBN94+IxTEJVPnS1JAympNzXm5M2shT3c2NS9mowd/NI9nkrBBEns/27SRDzGHg4bEirpzNl5EHh
8Xr2wQ87qI1qdkYSsK+cyZyIKBf3FSTxakgOeXaYbLjptGF9cPP4ra0enFLdaEn5qglFpCZnf2jC
JKNAsRx1ROPdZHvGSwkT+dfe8dMhQOmnVnW4FBl6Ql5biGCx6IUtjG6f4bgsnvrdXlRtLfFU+mYJ
i7nKNCCLxm3VPPUEH3pknU34pXMfNIsvn96J7bKoXp6sUcuaPrMxnHbchNeYp0pgTE4mPhPcPihV
gfyfrczOG9iEJ2S2cInummVtevSdY3jHxy1ceeXKHT+yLUCPGqpw/NxhUpoNDErDOwGmgZr4tjpc
6wntYK3Nqs83UtKHnvF7btLzEEhU/mGtLSjBf42uYqPuQgHbRDRjyVk8/PxDVqRXVaCyf3DmK5rc
fAS99gpUB+UwL54RVWroRjJh2MgSRwU5B2C80ZS7ZHRNuwoKlQmZW78spzwZsfL+Et/aFz+DuZcp
QlzG4/Rs4z3xh+LY0lBgqT6wrFORIA9rz/425GMIlPdRl4RXe1dGETx8FLYPZmw2xKGzOdWxGSEe
fEVjOZrgd+cUIwie1UUjZxYsX19sGq1cgEQmn8+oiEYgmtCYuSvz7Ck+pbVoGSWPw9C0jAAlcl4P
FHjC62fy8dmdCCdhytt5ro3UkD7CAtH8lCAkibzo6FaM3XvuqUzIVJQVB1CLtCUQtFBfoRDon92m
SLuErnBgJig5e8ryh8Mi8zCmkcw26dAMul5GpR0u9GupaBPH+zV+/tNlFj+5onJS7faycAj8+VBZ
EKJW15t93oAhS4f6zNxH3b97vxwsnu6zvdbiK4+Lv/ldkdSjpnxHV1JIqBifZn5hfH9wXTOQ0k4M
RX9FA73Ji7oRtEqArzV9iGbaNuuY+2pRREmkXQFS8fFhSDvXIJH6YP4IqdyIT5D5q+O7p789mOB1
OL4nqjZV5SkufYqk7LGXsf7W4P5a+DOsZDBk4uzTW4KlcAIA2PIgrViufh6A4yFHNsTOyjL5+lZ3
S97w2MIO9EV1OvY8jFYkPF42X1vhUkJbrfSBwMDW/IYXbVDOAAACVdwu3URE3VG/G8mv+lQo1JMp
r6iMt5zCOTQOBl5iophYW64TVY6ns70EDXWxnJgJBG4XhlRymQyzffVXVcUcvam+5DS82Y0ikZbO
ReTUKuIqWli0JFp5WFOZMVKXuBW2MomXTniC6tDGz4OGoznaUt1EEbPyFK48URds00HEibrmdGif
O79Txn/BR9QsC5D+AJiqERnoenermmEJ1tWtdb5u1G3zsHs4R7W9R6IFLJdCQY2qDFdEYuDlEr3g
2VPCxsnOJEpf6VgThkeRsKmrISXE6YAm1FO/qmEDq4w8fMWRxNoeOPn2DVD0TEkFKR4GWQIZPge9
wewJjrTDTSw/6W5REuyEE0Q7fxTh9hIO2lyQ9tS6FTm05Dm8oeJRkQStnkCH0YD3HdI2UYmF+vkh
Wjl5PNniEqap5kCBO8seU7Kj/r/T9xrvWC9qiaCWeDyvcPo42rWAUD6xXcQfEeEIge5K2OhR/YAf
MZiGrLh9L+oorwB4NfvR55RfrhrvVXhTwUGNEFFBUJ8XNOoV2X7khtwzernqvhp3YIyy7r1HXRTi
wAckhNrho/I0DFsgDM43ZuX767y4yhNbnFZkp1+fqsGXZiHtQ1wY0Mhlc6Y83pWvJvDM3VyaXBFk
Ajr96zSZaAuuMBEicrULNc6T0ipWWqxTO0Kfp90BXCmwJTT5c7YhIPYjH7XaFe2zeHcqMhbl1GNS
GF0gKNxIcJ1YGKjRj7UpMGGGpsIEITwz6XJtjXzopUZ6lOGskL/WCUSwEoGXEYVHNvlBawthNNOi
CHr4O55YTqj/FPjVJnnO2Vs/MIqRB0QXctPeLe1LMEQiMZi+DJkYmDY706djB42gdV8ZCpYUAnQV
VdHVsxXkfz7kPW2z3tR54SF7tjXftJRJfa/7wCz3jMK2XJxWr6TXdBXFa142SrGzuGhncnrgMj3K
sJID4mI2i8I+V80wXduXIfPQ/pCNB2GpiWZhAsNDSy/QY947zhsM33DZoqh9kURW96LkELMQIwrs
9jSJ3kFSWJRISjp2PpgvoRfLxgfw8IDbBQvRtQAkpPYKCSTgGjKM+oXegHoUgX5pSmbB2kHVGYnn
eprjqh969xuC5AgjuvEVaM8/y9VvJJqdIcM75R1rg9SebB7buDWHulwU9/3ldgvEbh4nkR5HTGeq
HLhdFx8tkXVbL0ldN5BcqIdiITXDth8ZhuBDWVkq8XsqWnRm8doCov+fUJrArInnf+cN5TbE/kox
jhXmg1p5Etc5EgV1UjPH4vatRQERdsvKLb5szX7dqiO4Mr87sCcgcmquMoQMZMhKIQ4+ktghkewV
AIBRdf6TbbD/LMLJQmVufpjV+skRV8IoDo/5qYIvgEFxniN4ukscDTKhWnwUo24Tp3jlQ/WV55Fq
Y8xmjwMYatAmW+Y3t7Q2D76IxXUmr/EmqTKtzcOD1ECYL795JL6zSq9SFF0A00JdYhPIi1fiqcMi
xKAD/Hy1v5ypPneYgfsjSbKZmsnaS1hH8WhP8P0ChBNGmBx8oDJsp12EAZi1O4+gTQamdWmIrLEp
8CgJjOqRYA/ICmZRRK03PSuf0r7W2T8MIK5cl8dopLUFiP7dJHcRxdJYs8sJamcdBOV2TyGdI1zu
tO2TCI+VO8rKolKicbpPOqNDXu3jc6vdHby3VdRbBqVN6kXbaFH7QYqJfsipdEudCyOeRa77a8Zw
BY0eTdYQXIJPm1XTlvRlRNlyYfvOuOlV4CeDJew7t/4RXHC2zbyVSKQMCdEwKEKPMbImuSF5nGhR
gPwkhSrC+8ICHe6lAPABpGT5bVSxIgLk1hJ0PYuRhTHFUkmb7TuACYHWsu5H2C+T9AE/50MJ1Iic
W7PXKxTWBn08Ad2XAWeKCapvLEpl5W1GU9IXg7V3zu2vtBoc7AgrjteafdlV34jfh1d08a06boTV
AljIxXRvF/2QYXQI52e+DLOwms17kfJxhN5F9Pv+tt3uq7d2DqfbyO6X8FS29V0PRGoEdhvAgaPt
YdgTQAfl3wv0dL/ySZ5fBYWZ5+x932ozWUFXxRImMJxZnaOg/Tdw/Bsrp0U0T+lGYl8BWRxfApGP
+8U8FHWkwAr07dn3Qsz6kDENzDPl8Z1vZOk6XiEDKEcVzF1cGpLxXgb1igYDH7gxuUfo9bePVFtz
lb0V9Y6MWHPxCZEMtIuRYT7aJT8ZAVEOCjWJ7vjlWoL7Sf0yXXMMSTZeOoaWi1OsEoF1MHaSz/f6
HlJDQPu+mkVO82n8RpQWbZyZRi0n/zdJo59gbKNrzrDiC03/PkDbJi+C1JCj4DxMfmLFmyYvRkG3
jZ4OlLpe3Ppi7L+tEQSYQrf+z1PSYxB1KznFNxAG/1jOccukCBDJ8oejjVts+EuW4GCNVOFrU+DY
ZddRuZl4V2fGCHoBzAm016eEkB5DTJe5mTNjwVN16FAu0QbzE0avC18JclNDk2v59rsPLWRmP8Pn
diYSt9vRuUr0h5D4scgHjjtsWqRD0gcRZPrMLVm7kyNSgFC++oNgpQa7UCrdYRNK0r9HX7Xpgmv4
NaBrI+Y4MyOXiGmRe5pxGDZF3sBceIxOQg0O0j6rj5yekLPy/CRp0XLtKjz0CXFcsP9nnJgE+D8L
22GVsk9jSHIJn6UoJnQqB3YFj5seNR94CnrB5PrCvv3JulQ17DR+lBz8locvM7Wh6u97h64BM/pz
fiFc0DmNkwFaFd/LNUZHwaR8lCjcZrCgbi2LuuIx8SU0UjnaljdMjqCefYrCiiyDLQ7Nc8FDol8J
WpmnRud3T5NoReUDj9LEvnvyES4JN7HmoEfpoiT29J0ekjDPUr324JFlka1xqGaU5WwXgJCVPHcG
6plGgaopHV28rnbh6nbStAqxml0T2Z/VZvD7tX6Iot6jyslNAWPTVT7ZS1iyNaPErMmhgWFoHkYo
tPBx4NVNGnrLECutvavZHPe+EoCFPtEBwNtpkKKcTmUCix57Fyv+NGmyzZ0wLac+CsexudUWeMb0
7VTDvaGNSL2+QKApVZF2Y8/ftdgHHsPiQLAlPUNlcvu29A0+Pw4ZvHk57r0PYRdJEcbp383VCCbR
q+E3RINEJcRf+Ondj5+NTj6bWO5AmsKVYPa+9hJmzTx9wjrO1oXGpbC/Mb0qCV3ZKgOyHIA9LDG/
N8NChUD4rg4azBZjlWNTizniHAT7hrd2iDlIkb1qUjP1QHMLX3lDcOH01DFNMlf7MQk4vNiYoj7V
OBfIpybcxBxGi+XV0Qc6gdelcp5lBFwayg4W6ovG4l7Q3jWTu2l1tVFBBBRgt2uzmQY3bI5wJ1vQ
twMWA7vSA95v1TxPu/wMX08wAzS9h3NkHMeoigwvptr06ABS6Bzg9Bw3vUCvAJUw+fTPWR6uO4j/
RFwg4ch1WqVCTsiPQAq6gbK1KwGR+eGtbtz3HhYTyoPxiOLWuX5pxVPYeykIHtfiaUnaYXroC7+d
M9SkHObutI/WoyDsRYES0YzYZycQ/JCxvg4o9msSJxfrHsYYJjN7vr9cyY6AucNN5sKR0HbyVrFK
D3k3cCWyM+k413kC3FWrQwDTvY+oPPtCODjhAglO564VfcVI8O/pDOZJtyH/aXTRXwSRPx40KmVc
3arrBs++oz3sgL7QRLnb6czwYUMBCMho6AFpfsA0vreFnnsvJWplVf0VTQfSPNhtzXl6xTgQOTc6
5eZZ9XNSdI29XQUoBAY3yMpDriq5VRw7JGyxc6nxDjI/iwKWyZk+OQPJ/ue5feRDlCfzgEb0dlRS
BC92hl/tJWocpi73XIlcDxBrJ3VAVip5HVDCxSG7SXMvuZOBKYL0oWzUmdjGPC++kzXuSjtfpMy1
SaT7Kknwcx4Nh03moMROOvl9O7U/Bkk/+9iP8MP5htWTWUeyfn4Pg8nZvbvQxwmP1YeCsQ6HSKUn
D5tQ50KpHr7xSb2Mudzu8mWFCeLNjI04GvZ5A0C0p4750GEpJTfrNlLgIjFC+0t2hln++/RN5kfH
mjF8g1UpjWmwtXVilFkMHhR1o61bLcWVlX+3GaP0C+ZyU3cXF5hSUm9vhRmpUMTeMBf45JcAs8qo
0QaFg/SBpr26GkO/3P48phmxdGj7ojJ8xp40LgaLMgxkgmyeV7pF+o57+q/nhLtGDWbQEJGyZiTa
VPrhi71o0aTk7atIqEl7PZMqep3DdvyMVU2r11bODu4U3McfHrD/kwANzCrlw12Lm6wpgNy+k133
0KHI4q2zBB3bkXOqSt2zwTAAd0eVSJz+GO2dbGzd+derZCMX5rSutAnvz6qzqSfbg+JWs1dcaiY1
996GcK/UHXRCMFUhuOZE3yWbJsDQUEIkqtjhzmHSEJb30MDKHh3urb15xCaPM1tVAsiH4A3VfRfy
DEY58pkSThAKb+tRKPKaxSofmhRWJPgGu0JtJGGTdZP22ui8M3T3EVSYoCRm75RpbjWnE+wfdlPd
wK1jOGLHNagA+WxZSnpyeTs89VfE8Ncmg1SjHJZ6MV/B7TLVQUQBTGV75ORBjKPyHZx1v8Tc95Mb
jBBFE9flw5WQl3p/qVbaUc9HifHCfwv+Mr8+FUgLrrkrBBYR/lpxeuiswE9vbis0qte5Xaxrgxmb
sa10ZPDZ9O47W2GixHzPOy6LnOzpihMuFvk/ClJzBq9fGThmCBezr45Z3Or1n5x/wmCAp2hrGXP0
EvUGKrN5O5whYJTP2Oh4wwibav5//Ybs401kD9aWMx2FA2NAqwrBaZH1iFg4UZjpHw1PHpi1yQ0W
IdDhulGw95MXLW1UI39PAjk8O/X6B5MjhBWg9cD4liealt9fLDrNJ3LMxWEQUJg9HytOvzD5nmjI
uQMQBuXe1XpSb5SM3p5H9izrYXGX0SJhEZLAEu72EWgCERi42HVTHjqWeOA530AA7RW/rU58BwFU
fY3z3DfrTK3QAdSAZtbLUUhTfgS7zK7T6lqa2/o7JtOs6QqkAd54U5QmxqpdbfuPHTvofD0Ya/uq
zfLPgJwvGq3Zps0D7RMTAwHDG5KwIsn/Xa2SLSzhAd7tzlhNuVFXKYU2qI2yD6gheXP9NjoGU85Z
w1MoAKIe+Nu7o0T/RgElj3WjyudaSdkX8IU4DfpS3Fcf8hz0e/p9dKE43aYU47BIUTw7XXM31DlD
ZNyWPDLZiXUuMHx5MPqZ/IC2g3zYNff01QCntoV+azAQZx2ZZyek15zNemjyt3XU+eSlkBGetG3o
Y5MK2nwK6DAG6l1lA/p++H+M9vdvgK0qtkFhREfpFnShAihWTceDH9Xvoh8KwbiKSxlv2SAhCUao
8Od3b+Hu4UA2q3Zyi2MSx+eAf2jt+gN3zea9H5BwQVKwbdPBeDjrRG0WbGdnCY/UIYJMZ6hOoiq7
PLp5BaQFqbtwiPIlWYFGLSd2jL7TO5Ar6ebP3PtSw/0uXwD7Y4+i4619f0EclDn1uT3a6fa4TC6T
iHNsdyBI8v1qLIAdkT6XJsK7bcQUejbguEW0eqvDyDZJ8vPIy0O8ZWeG2mnO8Eu1yThlO3cnKqRy
ivLntTg3DJFE3s+w+NRQK+rlNyfsvy5UECJ1Ce2gYvmqZi++okFmS3ibOI0KGG/v4URWRJmJoNOy
jaSg0uwQ0u3gIC0mLdgmRc3Q5k296jbP9C9LXLahDY/5KLNegBkgX8bh4MEF8D41pr3ZT+Z45UiX
rs7EYGJgOBmxX821IoNJdOBWEI2gr3lN9tYQqhVe18eicTgzSuLmze4FrYu3iVMyWszucmleGLku
gLjKEmOOlnherJvZOgW1m8IWBbvnBQe9fvKufF3bNMXVPomwOEBEhaHLckkU8n2/dduwT3ikgzUN
hDV+9iSKPQDGLuJzglc5tBnnFJFGcQVmexRvQcVYjOiAio2GMxlr6kNBx4Yv7vTUBocUC7cVcxGS
iT939LaTJVJajb5WwQEuTPvknus2xuAj6RBZyZTtv4SnCMEnW81DqU4nacy38iZmIPmHudFmNKAV
cvcFrS8SymFe4iTMeDflvYVdLfc8vLLxrn7Hwjn979WTg44681Ne91Q2X68lIzspXV4lwo+1+onC
2lUoCM1qwuGJO2pZk83FSJczmBQFGRm1xNF5oQId98x/cxT+irosyDpYnuViDn+ZUReI6chltiwf
gnwgPvt3HMsUQHG8qKTqykduH1RIt77jIujc1SMCfe0UtFyH9ZA6mqAbYHkIGQiAtacWjG7ywdBe
83bo3qc06dKOF/IYAvza0ulDKc7bZPTV6Nxambsk73exKa8BdtmP3xgyYHySYccxBMEkfF3ReiMd
k1SiAjFIqdZzpENX3qNwveEvKPsAjUoXFN8e+h0S14Y0EX22LDIaJrjKRBaOc6JxSuOPdXXqCPzX
ibABbwNwRK5h6/vGQAgqhd3cgS7USz7bhoTXE1Oitr6uSnn8b3q5VbN4Ti2vg18REAKa7lDCH/6O
FLe79o7L8uGyRL5qdsyLKKAsS3Anp4eO/ArW8Oa1/jolFiGv2Hfwq+zCM4t5TYS9k3W53whA5sxN
dHJzyHcl6o0bWmDs05WXTVIB3G+knzNmZGcsODwIJQpK8DlWf+LYjjR08zpyVp5euotynyo1T2HR
6VeKA5Tce40oIb0K83QF0wfJswLUqm/Ka4kPSLAa7fxuGLmV30+O7BdcSQT7V7aQaqvrc/5jDuN9
AblLSEurA1XSO2o3ySvGVaW25Zdd34LLynURDQW9YDCPAf9gvQx9GvVQ87POhMV+Rk3GUH7k0SLd
yjisaUcTBhUtUiliGBn3lB403a99l2HfWEFNUvpaP1cF0LQxn0h8lip0R2g9jXI2HpfJW3ALEfje
/vXBpe5pURvfI2RIQprhqnF7bJ+81q9+mthVJPcPyKRctA1CWQokfWb3Ag2tfXpRs4nTm+L2APBZ
Dx1oxpy0plBc1hfU35Ntp40KxJYOFhLpX3gSPbus/25mfN8a2F/1ydVh8h1JDkX/dxXotRms3d7v
YHGK6FCdFN8hz18XfWJK5XM3aQzQ7tdLtcN/2k98HR5fZ1HuAeXXhWOnA+EGk5lMmEeKYA04ycCk
HEiSmHPl349GzFa+w6Le6Z9FkgAlnXl27f84aGIzbR0exmil6h0L3aIHzeiRCNSTc7bxHLLXdX7D
Ea05fzc76czF8Y7bzfrrVHXPeQ0IPCqB7fQXjuvUyjDZnpxe0/6knmemVygaxhpykXpHBdE03c1N
3FzG2kJH23vZrQJSBkIckIRb/8BCWiyeZpmM490tfDaxZnSk0qRckZJDVMsMk1n/5UkzTxkhUpup
8Vuc/0iD50KIp0wpZTFappoPZz6dTWYdTwSj3D+AQwfgKwVRNxI7vmSUGounSxLihhxvu9PNjoG5
suSU/MMwXVMT4pxvCJAg3kUVaGxdRPKpWEmI/PXuBxcqxk6hizUmqjY3nOB+OqEtl1OntUo84Exf
6A8mH8BN1vkBNTCU3VKFO2/VRc4soUvg/loErNv5vhFdaOq09bPl7KTn1Kj9XOdQUAGgcF5GrA1d
sQqzyidoayD9EYyIZsnOAncBLh/4njzq0DdaQwPXSjWOQr/LZqrWiq+ms3flBqJRptfceyZhYSWo
pLrJ2GPxDpBr71fEnKlASnTTtSrXMc34uRL9R/ZabRHe0PZgOIvgRZSwqt/+3lpFlBqpq9XChoo3
waOHLR7ZTlAP8aEZbBf843WJOIxXACUQZVWCt6fHoaO4ssz/kAjzGxXnX4DGzWDgb6xtj/y/k90x
pl/PNp0Y8y8yl+4eRtuPYb8LH14LzGRobUX8xc0K3JNJroBC+CW2GzilhSPzSyimpOcQoA3Gpj7j
mXf2oxwBLTZ4wCAVUjHZ0AcZlVliHQ5ZlsrLgkOVFk1NNmy1H8hZEViurQSVxH4Z3HXS0OQbYGF8
CdWvnF//WoO27OgDiZnih/sxA/NnsHkcPiPKg8kQ21h/GUI+NjxGbggiYEXZCSCcBIv9JFXrHTSo
AE9/KTkkmYu+kKcauKPOZjt2A279SZRHnhQ+hwagEQkFe9vIct3/qoH96fnZcpBsKAhnxGuVChid
xNm/8VVqJIHUzhgasZICKY2Kggd9I3PgWuBYFpyrSe9iKBzUYA45+6whL9nOLSWKIxBiYs6CZfho
zAMxHsZtLvM+h0tt3StsUArUseahIa1y18A4GEqA6Hnb76EDzp/vqKnIIdEhdEPmDQqviHOXdIal
Sfsi5xQ8IHQN7O6msGEjdA2feS6oRzsHCWD1zZO3S1t3lclvlXrIt+VYdGq0oO6v2J89ASkSoPl+
Ufffidtvr+rmEB3+D8hJEzfMACND/XOg9tpZmFCMEiIUAjMLEDLy8qblnQWhMuBhEZFuYvhpUojT
8lPApzhbI43itPXz4Y9O1AgH10bMjXveyhKS5g57raIgTPoigCdZ/3UFzGiE+v9aU7yFlA0Z2307
Q7lcFfdXLZvpunzLI4XxhoEHPjV30eVix7+0U2TiJ0fYdCRxV3aE5H8pJh29vgdL/0+guLKHlQkF
HVCnryzHR4JMr45Zuz3DTdOP5XFmVnW1P7QPOdk3V+6J0mA1zFmbzaQrxU5tBC14zP9PChxeCDU+
vKWGcJaBRfPrAosz2mmUVfjA8eG32H6erl9FRSxv3rtAM5JSYSpaBGv+UFmiuz7/Vtp5Xn6TINEF
6r2rckM4o7qKq4sZSjNe4CrC73dRC7zSHs7g+8T3LF6ZKAe2Ic96FgdHD+SGFC7wjLpxH3BOZaj/
WmnAEYIlbcE9uWXrVBuqplOvb+LzsD5BbJ3w1rFCHwDaNyolIddizJeSezfKwr3IBmDZ8aqSAHp7
+LW0Elou9QFfCE1nCMQKYODAk/2ucwKJzhBtHdsrktdMbI0lvDUNhCmV8rxVeDjIXCnTVOTZp0Ce
T5q4yq+4T89wh4AC1+JCksyCtbvM5sO+9a7QZwybbRdYW++JiU9TS5CC1/crIDlQ7pDmQFoizQ7S
y8g7aRgSW2mqfuSaoq5mB9NE56oQfS2y8fcgc5VcledAjpt8bm837Is1rvqeDG0EM7c0NigUsG1N
gYM46IxCy81CcjKXzuZHbJi/EBwZv4cvUoryYJ86y+TXOyrK27RLq7xfChuvdwBwnxTRz/sRG7C0
br39VS0tCIpwOIYaaZz7eeOkXSj1hmysI1gf900XRerzMcnfvXe/XIj7pm4Q9eoo80PK+EeezCNl
g7rbDBqUZ/oWVFNkiVmT9jIA3QbvqblRK2nmrKKyvQ3F5l+g08Y4fzO/KZJKjxFSFdPv6+hY4DKY
2Troi0NprEZAYeX4fA2R0/D6IlX+DmUiv0Lg+P4VRw6osJps9syfEXZQd+qDQvlCHreS2naqi60y
+H/CLMglQWK0cNqDlQa/mbo9sduakkFxdHDXuBX3Mnmqd15KNQwoz99tcQtaVQe3Nv7u5JPb00zf
5NEbvSGfESg5aYwuJDuCnAUg2pWWy7H+naakk01auTa5wNyM7DoXQIwqkvCwVXnrXldWZw/RxbLj
wfew9qjIShPMa2D9VuvHKoMxnCXtiWpAwHCZOmh4iPDeT8slMUavz41/JvyiefM2EX9QQlwJSOS3
fVILG6QfkA75WTgmXkxRYZG2qYXMXzfxXQNuCxOw4sN8vZbE0dSyHP3OOhXKy7AQdHuCVgBWjue9
uVOv5aJB7nCz8zWWRlacWcTy8FHCd/KSW/GptmnfHXLKEaI2sn2rzaN7qSXvGyIVhV6bg6SBRpk/
PLb9e6QcyPebD2yp//O6+MN2T0CaKeJwyoUdjOQazNtJjtU/+Tfzs0vcVwyHeOxRDYaBMxjbmwvm
oKotFyJzMpP8vSeuq1U217XSKgCsj05+KmKNE9g9GgrL+/joJZ75eHGNfgDj1rVAtRjFu9llUqFS
SDQw8oNTtuYarAfDh9tPui+gHP6dcRMzZybNqJcoyMWkLL0ngDJeiSjShShLaBnivBNjdNZTTeX4
kaOKGoogFVRWwfwviUUmGpNSPOneF59AulK04un8+F8TFYPYkHhTe2yulD3yMVTKmbpVdGdyL3b0
ePNo7lIrmH1AaVBsoGpwbp4dDxguYEQ6JO3Im2DlViWuXXAMfa1jIvR6+iH4AJRIaYFG3wXjb1VC
bTCAVuRB5+PLItpY18+FjIhN6Qf18tZaN22p7kIRjgFMPnOax2drViL3TsqYwH6E0F5vmvcYEChO
K4RyUfG9BgKd7A/8X1bkjVqfsB8sUpaH+kQWPTnQRSBjOqAIiyf65ZSqvnSDD2YDQ5sV/bdpO4QQ
7phQX44plKcuYfgwqEO38qjBXwQtZMMsLt98Sb6ayJHvkiXmTRztsOZeKYjnR1NUxRK3boxciGgQ
K/qOVSmTdh4mFyifowjqJJkvUBLxW8tKewO+GEhQVyUj5XLm7tCactaKPKUwmlbf7eEMZOkgD9fE
zDGBIsSnzuWFfx8vqCRhqYWouw11Ud9IeqAx6ahzai0p/AR0VJSILfpQDK3KCk8l+5ebEvdPZLwh
nRfFKkhE840X2QAI4RTPNVqynKJjZxEUa1XTIIkqsRpZo0V2crADRhLGmiz1AUFgIBqm5/cna00W
Nfe7DlfxNjhMQzx6+XJkUJzVH6snRo/dDXhk4tsREA3zWuLllrgF4AUkzKVZHGshBuLfM97kqh6a
AVy2VrBPo0AoY1RNFlj3UFswhtf+NFF9QJUt6z2u5pb4lYv/7nGPb9pm9HiFEAEWtyygKNnP66rp
2pcY8xsgym1XzSCWKy8gui18lMgS2WAkBbas5dfmr225emYDsEbx11Cat2cmitjJIM/kVW6xUSSI
PQ4yXyIJNUpXuKtRiW+RsQAeSOYNzPj5KLmroP4eyRhLk8ZHGB7rbfeSl48SVZ2C+lj46nrBFA4s
jr76apUnRLfCWNeuMIHfnRQXTwHpYSemUg/KEBWRqvqUslb8Bde5WsjZX0w9oY3XYDeZLKgOCq73
AN9AqUqlfOgAqclmmCPAceTrxtslf1L6L3xyteTtf1lr2bSHFO4cswLIeOyFeVymqyH1uNzBwVl4
9AP9j7FGEwMSCEmRmhAcb1A5Lc5/JSaKIch0tcZQBF6Jep5xDaoTzS7p1eZS5OStI0FPgogB/ycd
vz2igVqCpskUKNPkDMeI6Xe9Mgixm+OTYAYVHumvHN2dVlvjycPIPDcUCq1hPs56aHEnZ3BQs78s
XWi2ICcYyqHqk90zgfY8vWL2/37AAop4tmA2HO9Lt+RLNWlMZsjs4aiZAb+fDk2JIF9KGlwyhg8I
qY/0c8dqrHXTXh4fz6mctF5v08tiIKqXRbDNkeCXki5HzWrInx7KCIxEZUuzDnfBsyK6/gqURb+b
DU8mNLeYnai1NKJgOD5QCJr3uarR/JPUAJT5XzVblNWCspywpJm7/WxTdYwqZNR/FOyGL9r+5FwY
JNdLUz95DVeLWasD9v4u1lliPStSnJOF+viE52lRiEGvHAxCfOBii2O9cV+yGuANOvmJSUcLqC1f
vM9WH2e//AjeMFSUCr6vLcDnQxzTk5dUbpjeWpO8X2ozDs+q84zS6XKv9dcrtZP5B9d16V1poK86
BMeTxISmiIWMwSiYhSLa5Ug0+68gi+WOfZlEPmf+Wk1Nt73klR+NXM6GLZwzMpwya0r6mDQo8/Ld
eGyxirBN+FIRjXDDPTuTRk/fpsesD3WGr4WLhHrVLZyfSAewu+OGPsnUNA3RaQRWZ72A1YgL+cS4
s+OkQcPWIOmzb4GUl8Yx/7Uw514MAdIovgbu9H8HlFUDJH0UJbv4AHqF3SZG/7S46vsCnULYRe9b
Fn3zbSd8Dl2G+1r1qEWTnRyu4IOVYWWjPuNcuorceneObJNuxRTVQXnEhhZEa6Am+NDYMA6u/dzL
EruTrI2DoDiOAp5kKoeZ03hIIgpYC+pyA++ZuEK6+DFqOpzRzfTMS5jd48dVNeRE9K1xlDOu20Id
KghGWHAdBWlClP82hlAWLVCALF5XDFwx4A7yZPpJ9dncoB5Y9K9xk+eMC1ao2qrzv3f8jv8aJcZt
or6Ybiw29wJ01osNBjVmIfMNll5EMN8ZvMBB1RLNvHI0UnadjG17hhMPpsoSBMG2VwbdZj8gv7U2
g9z6DDEV1bjW1clEszSTfMXOMs5RjMJV1ux25rLqRJcPQ/K2TMjdnA71kvrIqoKVY1wtD+pA1lWg
Y35Ob433GTBCfuq2QPCidmmedmvJRmtDy9DYDll89en5lk6oDugptVvF/fgFgw7mduIYHZO6f6qK
FlOXyiZfiV4citR9gzyhO5USgl5iiA1UkqwHUMevjSOonPg2pQvVFynOTMxhyl1jl/7paUclbJrR
lk++GrC84ECCLANWska6YEnSAKIGzEbpCIOvqTrgihjbvjJ+qeLaXDecH+kuy4G6hZYWmiMHgIQU
RvDBD9sxTYD8csYrTI66XiqkzbJx+tXYFBqruc1fwP7fdv+Ckq1YYaMa8dmKNHPSJyuHdwTerSWM
mx34/ZUqNznTXolM0AqFbXr4RdnX9u9QkUoFVcS9R8b2KJwDZxnRoCm2W23pndTDecJ9klhLHEWQ
GxhKF0c0tMKrAfJR97/1Vvueo/vo7ItM/TaTdSvA35yCcHcmsYvDnao7LH/NkB0VhPnPRTZIR0HE
CINRZ8ujVFLeDocwkRKSy29YgCb42gw5k6BVJziFvR5BY/oE/J1TiYipL3f1jsy7OGuyHGqRsN4G
bItudUObdoEvPk+o/GAyiddF1R8rJcnHuravFtYd0FPcDA/HD83uo09OJZVkXUZ6GB3MSEYH6np/
2dLay9VGk+7ajyCiG3i541hntESBlP8bG0IqCpK66WNgCrZQAedFfc2Zz6gf4JeYIosWOmlNfJyu
FPD0qa8+efSUbCdJBUkRzOOo0kHmtaLKOw4U0vLA0TdfZjaz+Y8XJYFiBQktrE3hNIZNChjkh33N
U9zn0hpc6wKuT/lu2heTzTiOQeGzATpPB0I+qn3mfZQVsHcpQGxFAJdx/gpAMW/Kg7dcDBZKAkzI
N6HmKSL0owffKboDqeV10BAMaC8s6h+qb9xUqSbbF2JnwTAEFkAgaS/l4TBqb39ontAIbmYkRK3b
xAAdCIMJ/i4H7U+IJw9WAzK+PdaLh7GE/N9mOXifXBHMy0Ez/MvaSGmRWL4gCmSRDRH8k+cveibB
3cRi8ycIQgWHYN5UWJLCMR8zWmZWOBdI0SaV6cGl5Qh9iWwlsCtwBCSORpAdFaDFUmEPNHfAlZV9
zzf/BC4pAFVTaDUK6y1fHRNTzNxx8cd2vhIvnmqEhztyXTJhZFyxjCZXCGq1Pk3+Bo7XEiR8NDnX
/H/OCxHy5eyEAskVCwFp0BX4fa2wdRQ9kUj3GPusEINq9n7qDBmzMYeXtSNxFk/lHJVl96LYxk0w
mvivC5dipQIw1VgB0UIdPAfS6/JaYd2VLeh6Zvha4gHD8XpbKHdc42lE2KZd8d0Z3bEcfK1HBV5c
Iri6vTafbutoiNzkIb9SYHxFvcs4kyiaXr3pM7hnrqr3+UvIKlf+k2uLrc9bpM6XJn+7NWyKvWVZ
dciqkshsvCiJA307vuDDVpPESca7BUiNsBTNwPsivSGie8JHS8367Uc5brhS0S5ny9Dr3+3VCxRX
q49OqhRm7zG2OKgubnK2uQOg1S49dkKuiWmYY/Wg7vSZfjNVP2Rxmne4iAfBMakMjlNB+6NO0bQn
wk1/usZEhLQD1fR/IjxE88Fmw0MbA7nNYUO9naI+NKzXWVQDPTkcrgVxyF56uexYQ/57za7OjwZh
mqyrjJ0zUpGTUB49XjjK6mgur4FQUBqrj7iH8d6Z4tKuG42g56MCQ3tUCZ9CKYfQdWVNPRv6kE+F
PLOVGb4BxFnJ0C4zuQDXHXWgpO9QNdQuyixjVaJgkP6tPG496SaB6aoK0n9QSiLDdSBm/GXEfUw2
ew3AUJGPTdfU02AaPnvd8aUe76BRJ7SkwntjVCMNJeR9LkpMcesO439loxTqfYgnn6xh6rSxdxQ9
flwkUJncrk/1jFZKCvb+laavNIgVN01IUGiNSvcuuzWU7v87DpeTaOjUq1x12xI1ZOXOeLZSoGWV
yhnbJ+QPXzIzCXqcPFw+3tC+UKvm42EtpvjpXPbYPH8MyMwcxkbPejmP1uZvKUUKIz33bSPwKtVo
RKqgmBnQOjPAtGWen0ZuWwARVaFrX4N2GmUy7Mc4nBcXRxJmqE/sw8BhnRv8Usf0PERXh5MWjfWb
CT78O7a0WJE1idGMCuxybnvoEwzVMXSBapxVJWFTrgJ71QrcvhbPIt1YP3nFKXrdHFx3GmIboUtW
W7zPVfy5AyIMFjcS3JQTnUguobE+QgRM43UCXzB0MQKd5u2XBI5K1V1wYVAOJ0AOtXMfFE6Ny+Rp
LJGiaGVnHeZfVVcpwcOSYF6yJiL02JSYH9RveCPwO1M+gx20rrBQLqLjJRIb/1HTUfIwcL5ntvFD
ZT7acyBNGaHDsMsQ34dwhfgpDT3m3apLRfa6coyAq5yWCzz9U2p9VP6iXq/7lC3Fox9GHS6ayQq3
ssJJ/61Jo8AnZm3M140F7DuM2Nletuv6V+jP64h3qERXvBfirSoM5egCj/ziWn31JXbzNxGmjRmI
0Lc+tDb0YGoHZtoJW+yvsD08WjMZLsNma/Q6W/x+KB9IsfRo0WIGJUHI4EAnOOdVWWD4/7UG/RB3
jKBcDAtihEdwO1i9kR/KlKw6MqglqTHnNfpjXl4BlVLUzy5O+Y6N4Ds22rAzaSyYi/x2Jll89EJw
NYzggXZ/c1HWlWLovvyoVqB/BLBQ6NiO0gkbJaQgm3g1cI5x7gECqUqphCAGOgwRy1Htji1mA2vZ
o97NSsfLbi2EqEU/bbEwCHpj/prT6AXdQpOAWZFg6JYv+3KiQZqMlVqy/KxcABOwXnb9qaZMQ79Z
77gDyH8j3Ac9qqG2CqdHNS2seWlA0TKdOaLXbPxObVLnZ5lwq53bg5/smMwSXlYKHc2iw5udJJ9a
9lzwzx7pzL2J4gM5D/JckMklJW6R+I5eOfYjvyM5yD2le63vAhMxY8/j2/NpFP6XRahs9VtA3FeZ
uFOa+517FPTHjsBg/FrzOmG8eL341j65Q23QdPdVtNTVHqAwutnU5M8VC4sDbat55981AUj7U+fF
w0sUOZcAzHcSwIUiAMy5r2hRM/tmx+7PMBtPIsxF9NE2LpEYoZ2Gonh9303d2P3HkhfUAd8pdSWd
hOx+H9c/nQhW4Eql4NFGbni/OmJ1hbvRJiu1tNpB5cvX8vDuSbc4YyqDs2YudyCucDnZkk2GadHb
KpQ0I8lZ/PGKlYcOGU72b83tcV9pWtPxeFc4od0giAQTTYazoLNz3qDy9pZq3CL7WyFRFKuAfKJN
sQj++3tlH/LXHrUk6INRE9TzID2JRS9GnHwoFjJ2BpuK+9UKitsXFy10xhKFupRyuWYQaQbPmHY6
AGw6D4birRGBS4Mg67Gt96vdtoTpb0Q3a5dTTd1ZlF6tW5388GGKfGNsBj0FtHgRkhKzPph9r6t3
qgJtE7qLtGGxEwTiHGEDi+8KV0T7SAi/ukOvMTHCGM1lsHXEUvTkp+jRBU8u05hCjo1TW7Y2mj7S
qFaG5LXOIe39hBfit4ABMz+qEYGfiGaFdgrDrojq0Vj3x08JUB0S5twWeMbw3YvqOZ0RRelyVD3+
e1dN9zRjkReNVzS2q7ipVZJy4NubgttfIN/Fg06udvnzJw8GtsHv7RzVbYZQr2jKTpiNiPckFgcg
qdqJSHkf52Lv8yni/w87OEez4S60m7tkzIVvwo7jxhlrDcxzVDW2bn/rGM7V+OJt41RsSSMNqKZq
+iXOx2JsjAdGTbcaxf2dBF5lwJmq2ZsTL/9KgIxSddDOAxkW2IAhFcePdKmKSxMNKDuy2MVDNRIZ
leVhtcDl5KDW6Khys7aqbUK/oH7LQQSEFI0bmt5GhO8XFExyvGDZv/ASUhv5QAPbstF4kfb+3A8E
TeEUwGHknUvM8YIALX1z4yoVO61FLva3gOtn5fyHM+DDPsz9w3GM89v+c57uPFiBdw4dLRbwWWeP
XkJZ1d09IQ8LvnUAOGR7YEdM6fWR7haBoSzb2tLAwfZuj8gtpsobv74IgvO/jFmUs+wJFyZIXxBM
/DJ910rgWuwC8tfVX1SX626dXcfD8LOsq0xeTo2JB/kROJWZFj+HczMKFjTTlDfZoLG9A44Wws1H
L8mEpAtmEMv1SjOuyafitOBXWnYeAei0kKhCkpMwkqBgmr7S6f6SGDa6hAciaJ8EGxhCA1UPQUyZ
YH+fTTj+QdoqYIrVT57lS1UC9aYfA/n4xF7gazBtOxePB8P4fjPX7D6cYlJ9JGHYYAATDiIDJFan
0e/SYh4hfICNbb03jqgAJzIUzf9jCdzsKsdTDUjZT+EBO0TnMdyN9FJR0pw7TgN3dcdU8xLzk5Hu
NGOThWZiP+QRddoHAAhB9S++fqI3qW+zE8KnYZNFjBt/szA1eFuFu53Ef5XqiKbtcRU2/Hwp6+5T
Wxu/XWJlu05EBZ+Auyu7yTVOufuDWrcLtfuCfs9xO19hTtD5ECgPvQOIi/Zc4Jn9nbdUBQTtSWs6
QaW79/edKUOGhd0oJb9sc1UTY0/qEgcRwPSkpZW6FVbfodDwNlaD/YUFEoJCG5Vogjf4PSSD51Oo
tmYycIFMVKafiRITI1yZM1RUN72TaZ7io9qMn5NlGeQwnQfQCy/4qhcVVOzLr21o8RdTkPE8iE6Z
SEuk82sEiG7HWYwF4G00X7/jRb79MLeZCeNsYo4wUH+O8IVsOdF3XhORPKuDySzL6MqYYf4iOp51
caGAMVcpWk5B4ttQfQ/s8ymFJAdpKdsxhnlzAC5MUrz5JEWoOS7WkWTWphrcfgWOnQkS/9nAteSk
O92C57UGYs6uWyB1PqI2mNJpYwf6cp0sR8s3KsEYV67Nuf/16mfuW+F/ogce2pNcXoRSU6jEtghh
znSqoAg3DMF9esWkD8VFPJA9yHRU4bM47ZZ9Fn73O6tYRD7JtQrYR5hRZL/K971h8oGmeOOOoIpW
poSIQ+qwgg4WBAwbUu9kkD3pw+4PtlLAytAvK2cM2CWhsL88VuGheFAm2rVbgnvXEsuYF6MPaBO4
mf28mQhw4wJHr4AwMTfriHhIR8UZZ+VvGjVt1jKVCG74JtQFOJCOaJcpjg6bYD1EEk19qZn3BWTI
Y4t/NgJExIPFYNpyvlkxrkkjAkkOKEgcPIgRwQoclqMVpnsyfopW8Q4Nk5uN+2KkkX3mePgaqSqD
YgevHyKXmo2EO/tw9vX32k7in+ITAfqCtLZgQ2WU9aF64Shmqzt7xa+5/rOn7itNJ7NE3b0EVGK3
/VP6xWQOBKRsx6cyDJw05dAFZrM/CuL9Fn0HSUoDvm6mZ0wdpPnzbiDQldMbYiV6nFC24oueiYty
cb8PTZqbhzIwLyjjpa+5tGCnTUUznILkklkWJcezHGXGTNNyDidDBhHqE/c2sxQ8gfTMxxq351y4
t7iY0u8TDcorfksBvYVUQMCe+gWju6QH64oQaQf2yX5+NUpBiYq5t+W6kVYYYCiz7n7H1bH6zPXj
TsIrEYsL0a1ZS4+GiodCTAK01Hej8UjEXMDfefX005zMb7PJBP8on5PFiYAoddJQDVPjKAh9Z6yb
LqsscOaNOnZnVKdiWVNh0lK+5gxzkwPXDfEm7/qFIL4o+K324xsXFcZZnuJH1xQ5B+JXxlbHxKDz
vgHTeJoKpstAWmjxDa9mUjwamtJrkCHqwAlA4gqmUopcO0+JA1dnlZXwK2Iud8MpV1cUFB8Pz2LQ
hfdzIsSAX5tRPCPOJIuwS14tIFkqH8uuTZ51pAX2KPoPYlh+C2hm+d7Pxm+eTwZovuw66HNNMdbN
RZDNuSGrJBPHkmTcNeNVrcRPm4UhAtAE0JHxnLGCHexFGbXmVK5CPCMvbTvdGA0LynNG2NE+VTPo
/UZ4r/sRElS0I1Ter3sHuUjJkJYNJ2uBIKEGOW27ju8YMdZkJ8WcUt+rXBwpiuSB+KJOrzblXXYt
J7v++w21+fxwv7qc3ON9srTOKFdu36oc7Wpiw0qdSfCJeW6PAc86YBSkbsJJ7keUkeZ8DvqhEfzF
Dqw3L2QqcBbbYL1YhI7gmwnCTKMGaeN7kgpH8gViSt54P1vRIOaZVzXO3vgx//RjBa1b8QNCYbH1
f1khgjUFQhirlygIBRduwLVeL5Isl6ymmSYc56JkaYzwO4bEYxBIib/BgRTv2fNqbR5/PaFgHnQN
ZB0Eajr98Vtp+Mmz0imGl2c/w4gT1ODGH1mBIQgE0Y+ldZG7yvBEl4kFGq0HbiHNIG5BwMBHdjgG
JlgSEIAtgfqZAlrpdOMBsMXb2zh34UBnk82TRM6ZHX4NQYThTrDecdTkcJ86NVbSrU1VtIgBuiYh
eG8yaK5iXx4epoakw0bTpD3wbI9+Dd1VaWlQt9B177wMn13f4G0KK8hFsesRbz7Rg7rxYpfwRy/j
WM/Y+c0qZ9EiDyDRSUR5n9BpKf+m3jAvMu03mqJNnpQKF0w3wJH/I1kYfNJYFbXKYx2b3O8jWc7/
Ez0hricNYG+Fz5mSlUeydsVIVYjOpk3PjdgHT02Q4BbHsVIR9S+qR8AM1SkGuGX9e1Aa/S3HPGU+
DiGY+zfzRFrPxLvo2CbeYztwn2oWyMGv7VLnX0wVrW9m6m4J8yhT86JZqT5c/7VLbbowLOobDsP8
Pm3+Qy+OqaeAja91xNlnOqHCD0AEU3a3uUbqTIxqh0K5w+pBk74Q63QHRXMoS7YHygFXdoSHUqOl
V7gtOUX1vhmloHvfHnTxwBJobuMR0NwUmJMYkAzQNh3er3UK5SdqFRoA7noH89dp309OVeFRFqxO
Mqx/TbGSa1seKVDa9fRiDqAVwdCXYZZjfm9IePC6nn2MAb5nhKxmWLRz5K4aHY3yFqoPNTSxhT3v
R1iyAjXAN1I0PGwVQj0olGVFJLVUOtQP/s3/jA7iYOkXeWorNik0y5oTypweeCqo7+eEmWMxIZlc
7zPAjAy/fGKh23iElPjk9PQMvTSIfJk0CB+ExXiNpzPZaavxlu1qQ+5Sh8Ltg5nsItArYrQGilv6
nF38BEgRvlfR3iPElSdemzKvbf4fuJAcbQIcgoCu/MITgqfQcNLOldGsvCanx3LORT43cjbS9BeY
ujeIBTsaIwyZRdz8FK29rAM5rCJOuoKr5lidEEAcx06SiMsmsoryB2XYjqxd8MseiWI3ER5oib49
AP5H4NKoKhoQK9edLqfmLc5ETLCvW0ph7Zq+V2WR+1URrKGnz4rg1eBBs+g2goANTZI4T2apljfW
ze8LbIQdJ41w6EoWCnV0G/Zw62oHjh2/obwjAXGJW0XMxrLiGArd4bDLHaRM76hL0BkMO5C3/eUH
5qa+KWlpYMwg1Jl7Harr5n8QwzbxWwA5vMwfxIRZNaApcCiF0euIHXmjqNZg7V0q9bGymD+sVYEp
lxRytwIn6M7KntTfEpNOSyZajI/99cJAsXh1QhI9ieeJM3UnXifxglrhEm0cXh1mVua3zFxTeHA0
6yLjTnUN3IridROLfKcMd1uH7xjliJSAe6vY4VhJ5WygzDRZxSx5INdxJ5a6gijD6xGhCBQgL4hU
kdUhRta43AXEwZWlt2Mvf2MRwz2NtIcFpfvjaOtGr+SSKVI1GTEcaNznL7WGbBNDnSVdPZf70ch2
r9RXi09NT5MXt3cnpSoFF8Y9rqyYdgXE5Tm5TfMVlZQz4asfi4tgP+ddsjGeBDcQrL5obGDlQMf8
Wcgj2BjpJBRYxqRnR6NpA6jR32Ljh+Yb/PtpveJJb5ZxFnUnonwoLZ9am5RokbVXuI5Pk3dJdW59
90aVBwfkwKVpQncfqjWSoa83zLZG3WTych0zKmc9mf3/GGEzQj6/MJDfBkKl+ESLqEgkuCuJDNAq
QVZgcYBb86iMPh9Z64yn/DfDZ2pwD9I58npRYyxllcH8oqVrKDql37++LkMBK3Ig8f79nLC2hbof
Cz7gzK0IzmArrQlSL3lqEy0s/WRfahcOUCBhy+Fh1hy692QvKR3D1icnC1cZjOwpyB6Q3qaHOHWF
sU7b8n/nEF8WABI8wqTOanF20oflIuvQx41yuQ+dgz+JbvnfHhTO/sOvv7fAiKwhSdzTr9fRfy2U
fYJg6LKw0ZRhiUsa1qkxTs5Jak2249iSbbQFMKi7iaEZpT2U0zD4evf7dfYYU78lNmafrWBzUZHX
gAJGtcuOUkgDvKkF7jyQPAdMHtHVSr3Wr9sd5LobyLtP2XWEiEoHKS5MEf6otlZg2hn7HeaP10BW
fNtLYqJNwF7b3RcoVv8j2OL6OI9kW7zFV5g6B1GJUJAwl4YJS3GyMkri5gNu9cdArD1714yrjl2F
WEbbrR0c3XHhIHNEaMBe9eq/+oY4+y3SfPjp8Ar7t242a4KJOP92H7E7hw6MHsMvBBEss8Cbolj2
tvaFr4fDxH503M2ntGn+De1YmMnwSWV0r10lccfsfHW/H78V5lQcUAUyeU0DjjP0sr5QPBolKkyD
JY+0nv6fxBGDRkqrMxUML+xiHZxO8x81kFbsE33f8YFcAe9FBt3uHGZbTVoH6EJuWW+/ctoHK69z
qssmYVmDUfplL4fBivsgH5g/sTxrnF5xrER1YTCr3NBMIZ29cReUnZhgyhFwiK1XeCxVd8LoS4gT
j9FyIYqe6jvCSg8yhIaDnAVOgPh2dDQsolDUFFe68oOUCbZHVMJy13I3g+iWTr/p316gaa3iEHlt
qywvfwfaBbc0qGhlsS6qFnulL+c414B6g9JmQ7jHLhy+roe1FJRuHsiAqA3EGkBxvGfRf9+spoy/
Qatvarc4GECkCQ+tMNX+blFPTCIrS2M2hcFOstBRBROHZYGnFgRiNjVoRMtWAhs0ZSA6S3wOyecW
nqKlnKm6WjvDaiuylN/SrHcoTj3O94tL3l/VzslyLp2KGxsjGYMTrvvyNinapI9bLOeBHfucDCLW
iVU3KWy8phGqP022uhQNTnY+/ZrV7/pQbnHttTRy6T4snBZmwNKRx0VRj+uBWyvgJUM9e/hGm6Wi
k4lsRwURC4Ozbtq9c/3XJ4ljdAHRp85woEXsVlq3Fn3Lgma/slA9nn789fpO4uYfE839upXRXksm
1EN1VFQzQ8OJde850AkMf2JOfsBX/haLUaqmtKocVq01SG5/B7sV+eDIiTNzle2N+lZZX7DM7aZu
0TGd/XYAvHm4AeW7E3oxp3Eap2uZrxIHaGimRbJffoWtS5lfcU1GXVr2rwtx7ulolu808jB3Ca7g
Sg3pjYS8UOKqBWvLmC1t0EWzlm6p6BfQJdhQW2HSiWzXosUIkRfJrnTf1lHwD6XlBvpmKBhqJabM
xfYP9p+i3RPZGgAEWKPrdQevQfqZD9OnZtvn/yS5gdATkVJAK9B3vCZ52RWpjbO6JD0d4zr8l3g2
RV/v2KruprnQnRFFT0ndf16phvfSyv3Kh1UioryUWFa3DfYk2Fh5SzztWPXw5KJGggG6BDN8HWtR
syHubjWADeySWe5BB7+wL3eOriRz/7RwZn6CUtAI/nK9jXH1OALfoJ8V8M2zIFAKIePEL26LQ3GD
3XwKJl0UnKvjyH+HbI3zi4wTUGoylK8K8La+7ocKAH9miIf5frSszqkX1CzeQW8eKFbCH/0pJZyq
JMbQaEphDFnvRGVWpixQmieNj3X8ED4xouplujYzbzX7zMo85iZAO9yD+CQtZZ/vbz0Pl7wE1jrU
r04Vi6NC6JGMVCkZ0wvHUhLfAk5hY/BdiYkItMnRVmTscI10GvkvEzG8UEPjHnBaQ1WInfrJ1Mwi
NUvfSqoXAGCKwPegXVpKcqSXJBNr239l/ZsJmYwLQ/v6jSIvltWjxTQ7D4k6PUIU0LC3snBXz+ve
njmmEC/VQsdAX8/UgA0G8Fykps055nCajcQRoJjZIjA+uiHw9ac4ofehkGoT/hvE2w9RdY/i33oq
crqolLL+UnYf3hK10q/oEavn851YIkc0VBplfxgstXNlBrCy/RYOpOMG48eD7DLqbO9do+BiQHpI
OtDdztb8svucZO18RASpM+cnWKL3ozsyKxgOam7hD38MDiqdmRi7knYQcS/Qiw0tjNgWFaeBJl5y
kDbM0T8i7zM15uTWHfJIn5ex/vKAykTJJhxWb3TQXvkp8do/JAYK8Fgv1AeKRSuGFC2ANr1WH7ei
AOTbw5kUEsdU50GSB8Uw+PwJpS5CXE2ONEwP2HrJpgmup9B07V10f0MCSTyaarBN63mXyZwq3A1z
U57NLR8IXep0J2eIh2Aujqmuq008ORbrRbfnpq6xT884y5tZSu6HQwSzVOpRqMJ/TQZvLK+PUUdQ
+B9CerHMXoPP6ls1xWM5L6mJAdG+y14RmtyPNJyagyeJjzmCy5QJlANe1yxQhf0Qwg8LWplHyV1T
UMFk+oLZJQFxUv9F8yeUlAq5RzAnYKxtk12k+nYHuj1d+f6kVWBDMKkE5+5GBUt1zhaVBPfmS8sE
6KXG0xXMmdG5Y0/5d9FGeap9XkUEfm/S3w3+9J7s2E95znyEdbSPfvTS8enY79UP4n7VeReJS6Mn
D1YUAtIsy/CRBzHIMSbfTzHiZqSQGN+iej6AeHjv44v5llEe8tQkLH1IKi9x/2EOEX2J1HNNLE9y
+7/TBO2f+0jFwx+FyhnVLrPnox0X5aQwPBRkvldI3Vq4VbPow7xLJiziMUJkQo595hyuHmJDb/et
40pwuM/ONvDcUA7L8mqjG3EU8IscXacP4njHK6mkTjMLHuNGiK+/K5thCWnpHnVYdt8oTVPHYGYw
IrRibpBVKnbR6s64C5ttWyUaPi9cZ+Plge2Hmy4WbwA1ppsqSmN5+sz309ffjINI4WDhBM2dfAtr
0o+/O4IhzUCDMOYChOBMQMAFREoj8kIa9uoVsrobLRpVLDuAUEa4afmRtpiX1/O0rVCT9GIrzCkg
oqn5VM9vz5j5F4i9HIn2hqf9hG54cMz1umqVpAkPc/bSCOMLigYwflJ9hzgpAXPmZCfjlBtJxCAS
PFcx9DJ2i8ck80r3g236Xq+Cm4gKz6peM875unXruaVG3i/EhoGbDHAVqA+Y7rSh1ZU1c7fOCxTf
PGrN4KTMGmen4a+lz8oeNn/lQxt6wK6xehNU9tk6aUZdVZ0t2zaNxe9g0beN5y//94Qkh/Gq2zCC
RypsGiMW1ZhkPDfiJSmwzz2zqQ1EmlN3QnmRrvRnf6yIHtSYBatN4Y2kYIR6hC7HJDtmak1Nefre
b4LhgimhtfmHnjhrRm3M0l/HU8k0MpbNhrP/UypXMUufsLUhhbaOja6MqLxpZ/klSqxsTiAsIBBz
/MNr4VowRbuhC5qpDcPhIRuOptS2ghQN+NIiojniWowtZB7kHxUX0ETWcOJedYiG2fJEOx4onjIj
FDHiz6LLoYTR6Bt9uL45GYZn6tRfFQEvhj0qRVVMi1SLY6nvSJCZV0CiTSyvfnEdbmQeFRbvmF4I
w0D5nCAAofPFP7ETf/1dsDX3uRk8N1FeklFe1m7gALkPVKq/UPHJFeaY5f6KRtznuauz0sfUZVLX
OcHnfmPoHkvEz5PQxRNM9V0VVjelC66XTPNfBLtejgeLmVKKlIzAQgo+87gB+tWhPORj40+TOP57
Lf4MG/v/a2dIq944zwr3fTlF+nqslVKG8oSFz79HwTlDZAL1HKYKCmPQa0h0MRh1T6t/IKaXUeFs
SaBJ1oJ4gMgbWcgEwNYMsbd463uWMLLoPCJeJyqKfNfzesgW5Al/SffJBVCuihtxCNigiqu7m9oy
PyODhS/qQm9iD8V+LLgXrWqcxeGoAxp2JOMEsickEX4fBRkcdQ3ZZnHDp+TTcOkBVXK8yTwYWLLW
HjP8YG2iQS0rqp2MQCuxhQGA707QB/KC/aorKUpqsNBEm4CHgTBVhI7TesxRjsCRHqaClYtAiRz1
PEg98NP6/x/xcRVNaR/Nrsb2oM3wFLnxW2su0rkL8lgf8/Z4pkAkLwuVgz5J9VpkLU0QWgt3EhR5
CmtavzxXLoGQaqDoqc3xOSYj/Ff+cirh7uNcqokAx8dFAuuCWxKtTsNRaH5+lT0UiB1T6XG4k8sh
zuCP1oPQ1cRNTE8MAKswiU0i6vXAXMesa6OOJpj4xBNPL7xCNuGsPszo/vwvE0KRtq/mPPVhMcEU
NAoYD+SH93E2axP5qagYb2Qpnb0k68P3YCVTdgzZBBOx6lEyGBQcHGCKCcRg6A9KRTkk70YFPCLp
d5BWdZxxNapT/mTGndFK+gysF4r0Eb7YdM5rJublw4MTUTQ4+f0rd03UeBaWdEeW+RrsDVJ5Eb3F
Tl4lKC121alOx4/fkb6Sqa8LCfHaqkpYA44wSUYA23pZKHZYwN0HSv2tb3r/usnd42mZVf2VcFxj
TYwQydX/B+xx2043hzDxT2b5kDJRezzc3Z7p2qpy1ChQTYY0LPTEjwfSo4QEBqjh1Dhq46V2oIw0
Y+L8tzq1dtwFRwc1W7QN/iPEGghCBddZ/JjtBhE6qM2jpHUazL1JiledVhrujEPERh+qRKrdHrO2
dkLRia9TFwEYfHxprbiIbzX5xOUqOw+Bb3r6ob99xwu50ugDf9SXERxjWmMKumc5OSe278vGkYuJ
Vb345pRMd3oo1klcIm9T9d4v4TN7fNkWLg243BuKWzu8TlPGdTUk97kOpd8xRlk7H6xEoQXjICZt
mZRDdg+dEzTgaGyxXB5zMlzhVY2kJU59LkPb/OlVde0GkltFnHzuC0urMK/Q5WLdA4kLOpN2hJcb
vtI9ManEaLAkn4DrOlyeLdE6/KDLx1DfRKTe5E44tnRo1F+ZSvovX7xbwGRRaWmm2ILcvMap3q12
9z6iectGQ0F8Y4pRtsXQyX7/DXOQ0mcbQX1GAU2Mhu/kYcIRPxneZCNPLHWRBS5fRR88Vg8j/o0w
aFl58IxVoZa5yqQLtH3JbhsorBD4m+UbUDjsiWEOMW+sdXdaVjRlauomPd61Zpjbpteq6wnamUyN
MuxpRGCGeOfFQCqd24zGDet+THpP9bwenuewUya73+4B5JzcdEhIvBJpG9l9SF2sMkjJBdkjtuYg
8JIOE5abw1ygq1wbArjksPC+4tBLw8w/DAQ10IYHLvDO6H8g6WbFIF8kk3HTHDP+HOfIovhZtZQ9
LztQTVhEXzPvclJ3mFK5SXNXqpO/u0RJRyn3BnG+NCNntCeqB0X1hYTIWSem0WoQNno2XZmFKK+F
wrXwQ+Ro2z3AJ5jCc3VQuJvChA2pZrk00+yY8XKgQx1DBJwtespHQgIRcHGwlJfc7kq1Bq/syUUR
xeBeNM6h7onyDAi4y75ERwnfrxbZICqIpUICHs66flk2KySd9sk5cBj6HMBdLf3xOZDfZsD2oYCv
hwmiAGhNuZEcMwOzeOOYWVuRC2ih0jUr9JaLKMQBhEFPlojQ4dT/mmoj0sFAUHOe452k1H2jHb3X
+GhnM4aQkCD+7cxi2s5D3WaKTDpgXH2OYlwL1zcQzSq7roQ2R3kAWs7THJuxeLfmnrIjUhPSKee5
Sh1IdZsHfPB4t5Bm9SG2SqCKUv2zy9uFXlo7/4+21iiwi10Om6osudQh36VTBoHiffU5QJYkz0sn
4ziFX8UjmUyO50HSLAAXdg5c2eHU7O8ELyGWIGbMF9/s66nlnveUfkaILTNXWL4ZXOeYwO3Wh1vY
YRYrIWrETjq0qdUPON/Vl4lFKL5p2GW47bcZXaqE4RgG/GpiGMvdWIi6n5h6CEmE6RKZB4Gp90jL
0CXqewrr+5Fa2HFJkMcwjp7IHhk5JTeJ1ICnZwXJJFElW83ssL/IVbBIg1pGvBJBo1m5sBH0pHjQ
r53PtEJdc4wh7JvWhMalWNW2TiHNJM8oCQd19GFDW1JyImcAWZdyw92WoHkdpHycJgXuMaCN/Oop
cOMOMNwmYUtRhM2nk4kXEOT4+01T1hFUfH5ELvAzENcS2661urgwHnwrSllDmSkPKSnMnBnMHHNr
fCfvmC0f0yc5mRcCsfyn1QOwizBTWibPXCAl/I38F1J2zKnCCgH6MMFvuygAkSaNaVvcdzqMX/Nc
aCZQMdR5V+vVIMgap7wDtQxCkhl2x3YO3CkLbusvsEOjKm7kM0PGqsHB8w+FhbukIJQArPK0v3nQ
PjItIqQUf9FpnlDgR2AqjdmyqfqsYPPS2DegXJCcFDtz+PtgxQ2mfa65KoNjwA/Iypj9DR8WxVqG
E0glZzwDwHViiuNDe9J0XBArwqiZ7fwRL4bB8CEzgwHIJ2kJukAbpXf8uL+Ey+xr/RrFLvpKz9cM
+65bO7RmgbRnC6VNYvBnZTTF93v/fxMK7xQ3fRHOrEiDThrfftinWK0inVdzr+aD+NJ6zdZIsF32
EjiD0Pn8JoCh+EtWEYNuUZiCDNRDj3Qty5U2ZBhKFwvhq9mBRQtPmcTCvhRKkZmjDpdSGx7IzDl1
G8CXvC1PGSNsq39neF+OisKVvP1ti5odAn3trIQK9Aqlm7o4i5uQXF2Oan8zj7M4xHQEa5bnU3Se
rr4GNYVhqAMYWtLlz0VOpy9QbopV1rwCwSYN0crRV7jf5O4mzNmLGuGE2tBBr9vx2PbZFbqSwDMG
UEFhilGLH827H0WDrxNKGup8O9PO/a3FqzikHNimlb/r8SR9jPpK3W/4ll4kO+qd4+3PXyYM34f2
qFUott8glmCk1iYvfb9aP+5GaVrbddnvI0LHAU+VBXLcEUHIjpiXDpASj9wixaoi2riPqV7++P15
ZW/DWP31JROT6NUUOWy4uTl1I5DGa9WgO89xm8+pHj4W8MipwJj+wUcJBt1Hr1yCKNLmEBNxx0Y1
npmSMr25suWPMlgD6jQuF23tIcKLecXEnR2UEKPG/Do30zJ+qPd3slJhPZF9AHFzmmUTutIpAMJC
uJ65BKX3RiJP49R8gHYA87Y6M9YPnyIvEUrVk7rlWqNw5dor0HPbeLr+cy9tq+qKIOE5t2WsiNDb
wIZgAvUJTRcXrDRVNiJ8ABdJS8Jgpc9mgqffmFW9u7jaq4LjXV/osom1muytWu2OUeDkn7etB4oj
ceguMFI3xpi1CrgPL5uSAXIVh2UJmV6GBjxyi6Foi6im0FoPFj+DIEbOjyGb66cePoJlvJAc+KVQ
sr2c0mABvguEcBhSaEMkVAgzjp2CtebyLrZ9AmOkGlIvSr/iHiO6yYwOfAIDu7vZ1Zr1CDP7uKT3
DGGbRBerFPRfigeZqZZalFevz/c7mxsQvEAeASFF077FtEmjyrzUv0ODaP8xLwOmcE+jHKmcnX1q
o6ivDsTipLHg9FTSZYX7dYJ4xQg4mrqFjAlIzZ2pstWUNdZmdOAlrWgAshwpO++iJttJa1idxkNq
CeygTUB2jeDWsowFHO7anRklpK726UOAFTv8c38rmC/GGwl1HnpOiZFN1/gdE/X6lOYUBs8EdXm2
C8QE5ZQ8CrD4HgcjkWmERIfwqTuwt6CxxO0DqIIwY32+W5lpeN+y7IEemEW77TMd+FbuKRqvzw99
pzxqgsGVsfFqoGPlwf7WJld3yzFZiBdKL0GBKmT322HQy/WIFHJkiGYY4wqmRUqgsgDIR75Fon7o
ZCSJjMSLUooLP+XcQK7ZMH/8kzqYhunM8WLt420dZ3P/azy87/SyU3BMrrdoa9QiPf97+ksmIaq4
Jja6oo5YFizHlJUrP92TP/wHTd+ESLgi0HQQW6l7SEdit47cJiHMqE/l+8PAupgkABAVvfHtlE6h
hWlzWGjCRAZoE+gVwrzSOSCEWvIP3uivsOVr1tTH6pDNZKQQA/VOEHVLptBVutdXUELvDjTZoPUQ
QfWeRSyDEwwqtwLUuyqK0S4CjgFeE8nlK0PjXI9CAuliTptSFM0r/0TP+ccpcd+wCdtXJE8zBC1X
K4OBRmE7RCdkx/vuFsKniPEt1XmUZEPzITz7SXmkUys2d7OBYiaIBWeT8lWsbr0fQcjsmhlrg+Ku
Q2ORlQwhZh6FY/ydXpzEslAisvDQNxGJPQDj2gJjZa5vLk7s7PJC3VbQ8NhaZnKCLqQjSw2Q2p2u
GtcINPs/BYUYmQkkPiKxMMddWcT97t3agpXyuAkkah7eypUfJ+etDTgh6UFFuVbiEaj1JgK9Y+BA
AH12ADrphPQol2xNvE+LFAKdk//5yZ9qiMXfG4uJzsFuFMY5FFlQMzB/6XRCViQKOqKVgWnDvTn1
M3zIPTIbrfzSZ+5PR3NSZ09PTeydJhjLGfhkCdT7NdrCkQiI8PZJtx2HuL3HiG2w1GVAM7SvgMIP
auGEInn6eWNUP6ytCe3DPf9ZF9a0j8YW5XIRrQfblcGYi9cd0HcI3zH/ksmj2E1w0W6j2RQQ0JPB
YwwLE12uYm2h0iKOj4ZZb64KUwoOH8H4R+AEvL1KoYQAlIe7UukZaRwWaK4h9f8pIihqk1Mfg+Bj
7jn2leK8BvEy7RDoh6wkBwuG5s5tf4Iq2WBen9gXBv63999z83gpBk/8TStNeCo6a3lu3QDqtSy3
7VtWmLIp7TksctxpUFFdACSSNBWPMraxvHmQt124DXhb51J5TmXpfgfg1vpe1IiyRZOPu77QzCr6
JEvuUJjeFncUcm7PseRt9nKxq0wh+nmP1jS8jCNap7Qxc7+MNoNGOhb7gctbVi9qm8HjzHyYTx0D
jkgKw447CdE0vTDy0g1iTmkhkj43vYdEEv5k0vURrPWJVSB1lvzi8jtysy2bEGxDU/Ux8c2h7Hfw
JzEo0prpRWLl+BGw8RJ4B0GMwdCH8umBX8feARz26Xd8vubdsLNYsVTLJRETZKMMcqkczUas5N7f
6Y1Hy/a5q+yhGRZJmTx9u0rHP6q5pA4F8acgOsvwwFAjjSMYOCVfwc5rTp3aKqA8AesE/t3djprF
W/WscOQFg4LxJwHRc39wLeJrJ2jm1YbUdNukWCxcuLM/RR1Jer8HhYFEl9CuSmIRUvJg9dK52dmw
W4qzaejSYgBMf4BAkw7Z8ihJdDiSC23ynUgbU7bcOSVjK0mji3+klXI4RDDb5s7hDPPHC6dqhOlF
SCkoCN5EhGGXKjjhVy/1i3DKfl3NK6q+i0Gq/havsbazH4lZ3Xek1Koq9pC1Dhe3H85BHH4KY8oP
tTJzYP5rt6OdtBINkAe+Le8SQ4hk3uBSY0qxa12Gwo8SFojEmKOc+Luek3+pamPC/8VdP/NrSSh7
p7gNnRtMtt62krWTHS8futRmiZNfEhN5+hT/zrZRGchuP1sXBsD8D9Is4bxHJB9VnVruFPZiwqec
hwIiqe08l3cBubvyYihTELtJTQ50vboFwYYXN/GuoqflkCxg6jho2jzqSt3lm2MMAHoTred8qWRu
iUKQbI0xSXVncXNGmxZx1PoAH00+AWJbiYk1ruh8Z+m6lCEgxnZCR+isxSouxFi4hp6YzM42NIxI
KFPZgYtoQcm1bzBuv3x90fxEbwNO491tX7QbbXk8++nIs9f5g/4UwuHos48Da3bhQuXp/DKHOqBz
coCpjjcx9AeX6ohwOTnLHLMDBS4rVqpz90kCi+83y1n3atifyFrspwkyFpyhC5+Z+1zO37Jjt1xR
DEJ3cbBvfNOYR9IoO5TWrgnSehAi/uz5eqxG5ZJ2smrqYfDKiMSaMfVh7aRi9d7Wf8pFKJUYstdq
Q20ejj9DYBkVJl52Ltr+UPToHre60Iywz2B8vsm6uTlUJhBFHEdjTkiT8zdkd8BDS856f5Q8KhIf
IBp9tUrLQwgynYAWGk35P/bLHmC8fLQmW5Uq+3UVB1zG7uicuY+ubeoYwVhMaUE3VXAeKStgWNCz
WjsPpXFkpVkfhlE2GWlPb7NNf2aIqeon1gDwHOnK8Z7w4jwtBZ2pX6zOmYJ1X30VT8vPo1wZxwbD
uPyTVN12a0hqq3Ez+tkRepJTxLeeqpkqRZnHwpihMYxrYC3sct3W9G/pzg90j2G0i5eqPqOXzQYq
jW+1wwVTK3JNL+4dvU9uNpqOU8Inw9ZX/cpDg/d1vwFV34ufXD9pOpVNIpo0X9PziHzttNrAYerZ
zI2+knaBq1kXHwTlgNcqhste9jTcwe7gFrjqKtSm7BVr8OX9ZAYvV8x2G/vHGgO7kSvOryKhlZZ5
Kdd1HhFitexCs9rgcbIb6JRIGZyJBIhLN6YZcLh9Tn1gLYJfkBX2BZfMgYWehY0lEQS0SCDAI7Ts
g4KIzf/UzLRmXU6mF3S/wQ5oimZPyIGDlrboNcVQYNs2AqLkK7dYr3xy0V4g8jR6hnVg+kOQpskF
CxQVLi7F4JCHLb4QLJbsmDzIjHNO//XyN2tyWVVpnFhkJWdkX73NFoqsCP/Ap8Wvs9EO8wB4Pfpb
Rw1seRYSCaC4WLTT79fkc+9KcUkstwJwCpEcOb7jIrHEk0w9Xs/7hwzMslkOTuuGANMK1Ah+ruHL
tSeicOsPvw50NkQRBP3WGbNzwjs81D63AdBEIqa37PyZ5NR08cArN2IggvyAcNSkrVrDJL3LBnW/
3u/9PzSWHe9IeKhGjYAom3FR0ti1gamqT0aqKg485H2xcFSPabCi4D2ubsjaOAryFQVTvw/YuSC8
OezH7IbKqhqJmpLa0XmKm3zpu8H83g2rITOTMPj4Od3Vo8Z/mFMFLH05mofwJdxqnqAPlzmakzLP
q7LAw6Fk6Ixixu9xn5uvm8rwKVb6LDrQYdS7hgEH/+0AWYcKL1xoIrdmHEgh15ZnBQUg6AZFUFPc
CkVfZ0iRnUkb7Tu2FtcS/ddPJygUxiu83iAyWY0fB6H6STKVU+YZu8LGedfvSYYOiqlumpPWa25P
YJhmRD/0VhLfExk+P3/CgH9Nk8kUB1Rs6yR3FNpcIrtrshSkbXpjtI/+v4Oq6ffP/T3JpthBbL+L
y+AS6yeSfwjN3NZ9JVciHagQZlKkWVHE5QxknuhZ9l/u4juk/KvcnP8y8327Rwd1mjjZYpT8RBi7
YGse/Tl98NpGDE2OSPjcFXPLjM2MVo0N9huuiMMPQ3w3EbGdDLXULo2HVe1IUK0AkxB8hZz9h1EP
vG5kW7/N+6onpGFZTLbZ2wzsPXLG8xkndkHOPCZp63+Tqrg/5uf2m/qIksQNEpqCbPWWhKn2vSvB
fbG5DwO0Cz6j7Rtxd1PvkVq/YOuQ0S2HFcddD1KaTW4DYCR7p9TFw64mKh+SplLQ5Ts/NjsV1s6T
DfaTJHoukwDYcTiq+7VrtiXjObwjmRGEEsXXm6ubbu4wozSlUO++pPav2koElXZC3Ug7w9IVYBf1
zNBT382KZO3soDPFppSLfrTO6z8EuzHQjCkMZu3hF3GpTqevC7cUhZYOCWGA+pjyQfaovpApnpWo
pgdFqrEIgKvZyoSszg6+Kj3wxdW/y/hKcpe02XrrjcTRlvEiwuPr34dglZ8uXkTMnbzgYXS7uZlO
J/PQFzp92arzaj71IDQi2hNVJMZ4APMaROUs3iqwj2J8IKFzEpXeYx366REz7Ep0uuXeHKdLXjU+
SAtM+ANOWN5AeCqHgxPduMK8XxYGAaxUPodGwUjWN8x0yXJcHgF2vTqfSg/sbY1M/mgrK275AuY7
FrGMfxO0pZX05Wr3aTqk3h2sGsXQi9P2yV2WaYEnCkRHyXrCn7u1rYAIzVP6edIkCZanZ0eT77as
tu1KSzx/Za8q8/2eIDTpv9UwTZoDAuTAoUfWMnGq694nG2YEdrLAWQdpyFp/0/OrSo3bVEMlhoTq
h3/xHg3yovjtrWDFtB0oWbvwOXD9fZvJLMoB+Pte8uxcWdyxz/qhi9MpDJgKIErK13NjwraNRGAr
96NXNXtc3XarEc2JYzuL/pAE2HN/lne3up39R4jEteB0NGfeFmroNRa5M/KK/YkQNokoo20oXnmM
1JWGX8JLHY2mQMDx1a0GSV11DgDRKXBeqimHmcztjUfXnGUSjedLwRzhpIZTAoH9VmH9EvpDGZZE
8cv0IPm03WuuXpklZmaZ4cSZUcUCZkTT+/D/XtJSIw8Y/uLshalizgxYV2SrHmUdGVFXMqpiY/oZ
qWA+2w7WP55kSy5J5TTa98GTXsav+B8yU55XbYK8e8y0wSx9ng59EZwoTxFUIK+vHtvnY+VrOP0+
anPuCTfncjjTZC2Kq6lNzBPrmPmsk/gOG4nKhMqqGNkPoHy41zvMGDoLL9q/f0GBC2k0a+HUzXT0
xsL/LbEVd7l84BXMNzA256DbLOZFboEdqItgLd0/Zhe0yMQxf1Iqjm7K8VVC6QICw++TtgTdk8ZA
saJPgdcJd/dadFhcdSiG4VcFUsTZgOu4bSsUz1zz3YhcFXPM9WEBowepoXgTtFUK5KotCDM0iZf5
J9JOSmyXC0NVXbhja3TYMz8JXOJr4hgp4RA9ezbEBbRBd0S5NIT3x6WQ4vGuBHqrexPxLn137anx
0D1QBmTyAEcn/n+OCBxAkhsOJc/UkxG8GFHWIHbpZJE3JYWXkAvgVaZtewN/cOP7NJtHTHX+rJFD
AeNKmFJ7YZA1WNZHI4Jm0ETXhm8vu6Y7jgTBXMEaHUU7ct5fc4qGcVDAw6oytXFC0hKq9Jh+fRFY
V677KGVfkngDz5ckcbKQuZNlHEnojjuGcQnFhq1H15C5Q3hoNgmxqqUfjNOpwllXc2uJklcU6/iE
ZjcuSppWaY4cZ7daMaqaPR2kryJPPJlM++QKdxL2a9UnBIRvasVQ0QDxYgQ24QVghTHWf4B91Cfy
cheGEeCzJbt5v56buDaGb2UwEnB7Yc73Mi3D3/EzpAxf/bChRJ4s73hLeLag9jU9G6mLDtzhm7Y2
xNdMsSsjUwNmcKYUiuoKSyY1GZlpl2cNMKqfDlUj+ugRH6BZuXyOhkqrxd68j+HbFLJRqKV+1Ivk
JOsgvy71H1jqjHDxtmnANBGJLQAivwTkVenJd6M31wua26LkXXfkzgJ4oqHGeH3rqG9ZAqcDaJ8s
IVbsnZFFn7YwU7H9ikMcK/R65TFiGZ5SirGVxCELMHHTpj6NeUVQnce3r95Pe7o8kT2NfBir74z6
O3oHx5y4H3d14SLe9grQlMoi4zxWHqlMTz/o1c+NTlEWVQKW/DrSqBK9DucVZTzmJlzh2+rntao7
WkaVXjyU98AhlFiz1fGVhd3gXKPlTDqCuM6VNglDoImTVUEMB+syiDsdHPnOVoW7mNMKneQzT0k4
n4oAT8OUKw1869f6K6c3A7CjFB2C3NeNVmMVxmYG1C9mWUQm2TmLCRRQ7pnseUggKusqu1hi8ky1
cJNNdIXjTxioUAxbuHjDQfabqHFXtXWDMSnDMIoeDnugJG0PtZkIdCxk52x8uGKmYAo0W8h+PzZM
3mw+Q9kq65uAjN5U6E/4W+5USthHXb/WnZaYLcoXoTH+TR7BCEaw+RwU+GGGUIMLNlz7UxBh4jo6
0/MZBQk0yWiKdOkIcQJI5uMB5Onu+X4CkeiJAYOfFBS0IG8EnyDnC5+oaGNapArY4vv+9Tki9TWu
MGGVRL2OJeWOyEIopTJfAuDI+Q47L0oTZNkuD716VW1eYyASnQR+KwqRm6ujRy/ibaEy8dNM+/TE
B++OQqHQYG1d+qVtZeIKD9h1c+l8eEyJHkWEbfAids3YFFsgLC4Okcfg9F8a+MbTm1t2u0qjsDLh
HRUQYe+2JXSmCTJGE4rO08QCFI278F+qhjLHqdf69bS/2t6hETSDs1eALI/oHCLxzjQXMtudBu6s
IW3sOqJuqwEWI+jT6mLaNWaQiN3q9xE+OyOEmWfQIqEsCZRPpeFipiwhbjD2etlf7cDAoAqAUZqo
nHbMkIYVZW6qzS3pyImN4JKWNUZ2c3+3bH03EgB47NNsg268rmXjgaADFVQHMMtlBcHz8eOvprPt
dF0Mytk0D1mYwXd3hCNEipUD3lmexf7KG2YEZCsVerfiSA3DZAApS+o+NPcvm9t0pXFV5qH/P+ZK
486Q3asY+58TZUzKDQBlaqm4zKT7cN584UapStWuCkxD1O01fM5oleA5IPHYwNGpMFFbGikOaLMz
x0mCQYewTaFgPkw2MkxWdTnydc6Ou5SH8URIKOki/YsXrGmKceq3GP87vQ6V3AQeajbqgks+jOsU
0pqJtve43sHDsMNi3QKvqN4cQxnyU9/mjc4BXNtNWtNjrwHIp5GFcIR6Kn68cOzXgyC9dMXRIDnt
ToAwit8oH9qJqO+ALyhZKhDKdbTYk9ic2KDPd3ClKLl3GW5GScfgFdXAVjczoU2weLwE5ofSkE6v
IiJ8EgWWP6YLg+gbyTUygKBlLFWsL8IvWtBrnlo6p6yKSA5iK4GGkBzfGww1Fwzjf5wo+fVLJxXO
lc36m+7sot1sDQvyKF1i3HuEHPqrWrZra2SOYIUUiAittfl+Vu9f80gZpkHA7fv1kvRQhNLQJnjI
/FSIr/v00aAacdhfAgGXrIaGWFb4Q0xvqcPfob/ZPbpsgxpFfBxR9oFU61AZiBK2TrZqTruGHiCj
61SC8pjF1R4e4D5JfcwOsTDBrAxuZHlApXs4VKb0kc5HBKZpIUJuHn7Hu5RsourJ79VTZLXQ/Ln5
+p0s29LVQGzeKsveosUpEUpQ3LbUv+LEecZ7zJNzrW6GVnyzAyHP1G/nZIsr9fVXqYeXtMAyvazR
w64QWjvJycfKxKZSeskHb9AZtK8sgCAK7yIfuaUS4BzNPblcd5wl7LLaD/N3Mx312s2+p4UQw1Pw
mqEIWik7Ga9USEaS8K95J6o4vTdabdsMNh4eOxIqI4EcHfFcgwn7tuqq7H5M1KkiVmnwvu25Ainc
Zqhep8S4paQUIKUgYpGgp5E2Qdtlb/IeETllEqQFzTxB6RHQ4Oup46ZNnLg3PP2uE750rz9f7drZ
4XFJb5IOjttQC0P8CnrPwflNaCi6cTeKQIR6Dii036RL/TSfBYC0McK3wiVN19YszCYWKflO79i5
qHC6l9nf5q4oRkEd+kSdQKEUiYh2IthHxuyBfxfQ/HJIjg54hcRDVEpxqdiTQrweAKTrKxL3ZFbQ
7Ud1EW6AOmEi/Fnn1/GbLW3orsdeWjLnDsHDgsl3WxfY9O4Lk/O1D3/vm1+r/bOFhk8Zzo+nyaSQ
YLQOAVL8okQh2xwQQqlq5461jUi2otgO7gpMD/DwmKcxb5XZHOzZjuGIO4IiCD3rKk62J2WJTsFM
qRUwPPzCSv8ThrQdP6TZOY79XCtZDlgsU8qvLnEzwNARkPwFiGa07xQVlhCSM92yqMuwjj1+XPgu
E67tLCdBUoG8FtOSCktOtXA51iGsflFz1FMd8IQVv1UkX/BlNQLAm/qPWm0lzTBGs3Qhp/VWMwrf
UnwAmdgvx0eHbcTUbRHWuuA5Ry1QU6D3R+T+rB09VoS+F78ChJ280NxE0NTVVi7RsuTnxk/eIwCw
ZKdMKJC7CvP7Gx4gE5S4GYCj2bA6TJ3g+sB6m1i5fupNUHT5hKWiFEWzfgh5xmibhXzlh8wWzleA
99UagjagGXyxSCBPKb1tOyrHggi7a5ivet+T/BTh8DeaBmf3aDYBdp4Di2sNE+630nzyS+8Wd3iC
XEwWi0ZSdfh8PotvnqNsu44o4EeKMNzTbmjYE5D9LeySZVHP4xj0ET7CL9b+5rY+GCsp2ETEKQ9f
Ndeg91uxIMljqWN2vLjp0JTNVIZHagoHB1jmUUNviI58qCqwidFKajjvANhkK/3KhYtyk/eVVGrp
HEhSgwMQziSnANGb+mjEesMLmjaKkjLfz8Kb8iTUdv1ScMbIyFOIwCY1E8Ybwc0k3aEfu8CjSGgl
IRRa6TsEuLiz+4bDcgPmxdJ5lOSKw5NIXWLEYhTURTlDwP992XsQzIkNuDUWk+xxxctknaAVcgwZ
PAc3Afx4Qk0ULhJXQNuugzd7iZtWbRTBeMbjNDcYtr4SwpCJ/zvPnru6iypr1rqWsj480p4cHzKO
MPQwsUWmLkElUSd9MCKDcWbfE4Hny1ZETts1kdXNVNNB0FGfNQH1Zj+Za2CV69SB7dYp7jEkFKmh
P7JoaYOwHz+kEsll0zSgmO0PK3FaJCQZi5ZnMduvGYSQcB6hXxNHnAtGqbGn8AJKC6Y2rTbcv7jl
pzC5hs3nfZcHO0gNww5AKtPnj6FePLlBxA0rTh7MXn/XvTQWATgWcUMLKNGWFIna3aiqOILa7RCJ
GEHWTcmw9B/B3aJGTu9GsR2GqQZOEctBFGEFKmgb+NjTLLE/voqoGK0ydcegq6sVDAxp3BgyMxNl
1PSLECWuq29H6mcJWJmE/o+5q0ARqnIlhLJT0VwMd0sNBCD3Bgbc8uVDBmqeczBfmTjx6Vi3Qt52
ERX8WEMDWnoRx9gG4JLJYAfb0zeLa9sL6PIstTzLxPFrwY60NLxetAt/mUbTPQ+Z7RVKoHrLGfcP
yY2xiZHRH82nBb6X6N373WNMJD27AeEjlcITd0htFA+DNahsH2DvVDUl7jMP04ZdhkFpOeB4J0bS
pnismw1tzfjC/+tIAEOq+E5ZDsaOB8y6yS0ptr767Bhw6uTu0Q8D6fpVLdKkv9Sx8tabnZ9CAwaj
8FO/zvXiE+AwUZXkaPYtki2svwSQ9J0EPBAbY8hc+uv8Gv30zjP2s5NtSmwILafTBHIHr5Vrzv3w
kCosNABb86brn86/I54f5ZuF5qc30Gia1rhYmthV8X1yEXqT02Ok/bP8TaOBDCJO6nRby2VGyshx
Tw4X5EQsSfEksTR7eiQmTrV0pr/keAzpNAX+T5n+iDGbCRaYrr/dCHDU2bKGb5WdNDdLgUTrJpdU
Nsw59y3ytxgQ7mrDxr/vjSWafFMaJrvFvxsiZ5+RP0FCTmoopN1FIbDM2Ok1ZtkFjthH8BQip8NE
9Z4OtQy0gmYGNB/9E79lhSFImsTasU5Lb78HDXXVnLaPpo97J7KkNK8HPzzXuMrCeNem/gP/jcfG
g96Rjm+Y5vkgQjUmdh9fyNAZhQSY7gR2Ih9OJioNrJZs4g5T2NABXdUquYNXO2wPEak9ACspPRhq
1CTkzDnSYTyPyPrsxsj3xCzjjeMP3RsHMuPbsSJ7IJfYdk9h5DLX8VCs9DGpoM1JYoWn0/W4y9FE
4UdOSE1d/teXvpMSO3ZWbiyOgnOQ2KaoxMm48C8a0ObTsGcUESSn08X1zPnSY35FGem2EIkr/SSk
0x4L+0Uxpro+rqdyJGn1wh5oixB/WvmXYVbTPi76l+ScRdy4dIOmfrhWC5RtmVW+4BEgs0w/L7gG
+9fX19rPPuyq2AONOmkZoti+ATJjZJuTibaTzFa4y//v+ailEZ7UZ6AGU2OiDcfOvHSCmSInOtoD
lJoI1iyP17JALP3gLhueRNxXg67E9QYDQ9Z2X2oCNjY6RToXAZ7cz9ef5s2aAC7lQn5Ck7IfuMPv
Q6WFkKXriwHTIn831aHvqadJh+ECY73fAcLs8qSbBtoa7NTrQavUezXsI/zgaJi1oeBH6FwfYrc9
8MRmbK08LHnUCNVf/+iL4mxgrRLRbXgmyi/0xFhzHTIxTnNosdLV246K070TaGovQweGAKt2KLNG
k0O9P9ubhSMe8EKKGv2LNqKrLxG/sflonTzgzmos3/TuiW8YDdMp7/iVt2kAAu9Uy339V0AgulSy
Mx5FpSO/A8UN1Z0T7VkwyMLK9iKcEXVMvGzMLrvupo3sztn0Z7TcrrVDUKgAm08mzw+Fubc04/wN
nzTm1ZbnYjTm8jndn3kPzQOuxhCQS4eZ+eqPhzZrac0LrdREyiUc+HxwxOaCdSO0P2huPza++fcM
Bf0F0NOR2C0dax3LjV7Da4x7AEjVpYNtSAiB+LQuuLmEdgZRymlmtzNC0ixvjc88xlgpB4UnbPQZ
iL+xyU1VHxRmTeVOZcNapEDXDmD8vw39o5KARI3toPQgSxhmiPpSWQen8lWsw7Q0Jro5cQVDd+/2
eaWcLLyQgT/cXA2Br/EO1JMBPfu1nZBTLwUEgaIO2GQXpMxq8i2W/Kh6jN9DffTEWoqWM/zo6/if
k2/uU91wmd0syGpdTkPBuide0LMBlQosSQ310q6oPmc19SePGekW8KBw3l5qv2ypdFMKIiXrDOaK
29XyjLlcz2KQWn1iBqK88bLX/iA07Ug7OMBH+VTB3hdO+4MPU7M4IgQB/XLNcKOP1N0CsH/6uQtX
sPOpkx3wW3UX+Rpjir9L6K5TIQuts+nnm9clK7OikU1gwWJ4LH6dKfgWKdWBAq5HEQsQgym4zl2x
j3XL1t1VqNivAneAr9Vw0hOgf2Lzab1qLIM9Zji0VHkDncf27bkRfd/Nz9e4il9GcUU+bHaQOI9s
2mcGzETrv4OG7nHqMEedcEoa3sjMvq2vfGiKnlpx7gJX9i3OaVZOLKBy0yvTW7pF+/YCYC9zwPxd
sQEmmQC2p0omTc1vMgiG/hWLlsX0VGvk6pUt9ejMBwzZ1F6Nnritpw67w8YfyGaasv8fnuvCT2r7
IElpl9IoXiehZFECWbsAmv5US76NRg+Hfeojlfk39jU9EfEsscPGNh5++R1vtK9nUrPDl0BPZGst
qr3q2hBc9K1WHl5CCkuL60DjVB/EdQZe6U5ctRE4kEg4bLmjoIh2xFcRGgSfm4zCNhkLHzRnuVPw
HO58/hFnxgb3iBekXetNg3LCFZTcdS3lQ9Q1M4kIpSGeyju+DqhZ5ntIAt5V9yWV0R7Q1KIKrMiE
E2nDwWlsKvS37loLkeSR1gwNHW+jYWBHxGBaC5dWYkPZay8bxlcUBDQ3a9N0eTNA7wedrU34apkb
YoGYIg7k40kTGl1E6UvdxQOynt/OJ1AoRNjXyiXgTNLPXgyJl+xIfTgp7vAXYfhVPypfTLAlbvbF
vBMArwQC7xrEmnldVT8qjvIVst8jSFvTGBrJ3CzMNFaWljhW21z+UuPDDe0v9wlblmq0bxTaytN9
DWAZepAXVkUDOux9/XV8Sjh1r2znbon/SvZ2wuNL3MDhKHVcQDg3f1DEy4l4Zx0uHpQETwRQO+Yd
nk9geKjeK3p4hBbvEqrMeIOkfLmqwKrfWjWFJSKMK0JDTWksskCIVmfmFmkqqZ5k5WitDqWtkRwQ
8Ptd0JgkuB/0lPxkCjkW5b9KGxqagTWxnn09qwXyd4bS8RH+o2hBkpmuzhqTdk9x4ubF7n3BpU8H
g9tabuE8Xpq1DobCGBkgw16IwbOUHBqkpdvOXR/HveKzvn0KgUq9KkUvcE1eC3J078rATC9jm0YN
FSfc5/4FGIP2Xml/mfraiMcBZlYslBX4gdLLh8BG/TPQjpdR0P52usz0oDB/aj3QlY6Uecy2Bu/8
NesI3iSnke0ZbkZ4Gk64728Y/HIcgpxbFR5je4AcKHEAxcNuvdU5ESMwzCEruY0EGssK7Z1c7Lc8
wIQvg4PwyfGk9mrhUIeIy/NfRI8N+dOCycIC4cfm+rVW644/Q8lwaCB4G2+hidOdiovhXIBThGm0
q3++jktKunDn00TmEjVItlsXDcVxGDyyuQzZec5HSdJM5PBxw9clFhucE7/Eb4wevKFmz9ZxydR4
5z7BTXdIk13tSVtxbCnR3of+xV0Rh+FeMElZRy1tKl+9yJVO7+5XO62y19E74c5tAvzmWetBxKTM
sf6uVppAih+jct0SYs85lM2tJqbIboYSS9KwmJXB3JB9CO8Hx52Z+LFOMCvHcJHZf6YPTHRNm3kQ
mQGG4jJyn55uWsa9CcM3YFwdO/0PS9g1wBtoU2sbZdblFkrOYBBRxNX9cWFR4kNwWJKVbLUKSVyO
jRrkeqhE3+43FatCM6hB1LkqiekxqsLpfmg1snUKXfhvqlSzS1YHc21zYKSfqA8Da2G51KhIaxjN
MgRvinIplyt1yODgD/ISJNP1KJU6Vm2+6PjCHCQ+W/NaRHUI1Hl4rfPs2t3HysXomdJ3d0X3VCep
vc2aqhQDHJWND8nlsFdTS7RKeaZUoDLs0RvYtVUU2M752cKDgnQtmEdo263WP2+KutZk4YOegYmY
M3XgWdXxRpnwY+dMfsT+yn1oSAc7Pf4zhkF9Mnl5rMY2Dg2fvANcw2ksDpwQpYCfwERNqr7hLnux
KKQU2EYmS9CUWt1mGlcmPkBx4e4sxaZiUMAq2Cea5IrRDjo0GWfFAR6L6D7umpsrt8AAHU1FH9wJ
2x7zKANiOHVtxya3lKD4yoKQe34Rt+0ELKtcrp0k62k158fXxPPHbqjrkg87FUScN8knXZjH4VxW
Q3UYSieBMXYB+Z7Dw00+byeaEdjK+9lS2/8sOm9/NPmee1frXSsI1F+IuvRXA4VJTFSE5J18jWXv
xUilxkjPZvfXRLph8+e6MSku/Y59Hr5ONRmusb3NKdOz6c8xG1JUrphlR5o4i1Hd9eY/rP6GeffK
KTNcBHkJ45rVtN/qNL7Z5jzaya7BMhIjbwh+wKhcPdjSZdQg55JuEuCMJjzsxlvIzRyqH3/d7Mdf
MonDRkRzLGBoY8Rcf8b7cfE8RP3A5ch9b9EB3Dh06TuBelrTCY0F2z35z+IsaO1fNZkU2csalaMN
VZ8OxBZnM+WLUbcn+fHUv4WlYy6wgU3TK9vaIFYpCYrysAPJiUcPkKcTt8iCj0H/EneTdu388UXo
BzT7aRV4sLw6+mYapYV3qR8V/VJvppBxM7/ifJfUC/6w2+tnttwxXBLpZ/5r30+mqDAJOciE4T5x
ffys5/2FE3HV/+ibr6Kq/lcwc8+n2s814LExNQWLE9CKr4+JmII8ZsFnhYIgjoNxXU/aLdmkzyVA
FBmMQ1hp3227ZHKI7MdU+BdV7poRPnjrxSkByvxCsjJeN4TFmNsPXklRk/elEwQQvVtaueou4HQB
NWX7ZRAnQC/o7OZ2lNqjmMaG9Qx+OiRt8sLYwW+BaQk5mOJ+JgGh5loN4O6z7ldkdwA6nvb6hXJ+
PlDrJPmORI2k7vwft1UZArLX1NIPTlq/D5/u8TkNnkimEqZNcawENrZLgHQwb7xbVoOHX9pyVnEs
FRqjdSz+yt7blZy41PSIKU1oH79abDlR9MDZJOPTut4Jq1VNvE2xE8xD8kZs6mLueI8MCjqg+LNy
DCsPHreU1eCNW3fg4mpDHtoaPUlCsnOWsPE0GtHltWTvl2lqudfuE6LgcZrKZx2rX6YlXhtv1Z14
PyxlUGb0RuY+cPRINKcV4GvVfS5B0XMPKuISNWYMrmlETNfieY1FBnBjHCBdLktUJAtorPy+BWj/
a5YYdRWZi8Jb3cXOmZ5LYRa14blk5yP40EkmnSx8aRSV6LIPGY3PUlNcvK+4C3F1HsRpaIIu5eNE
pnUf0dVm/MphsB7YXjIoDJ4AdJKrIoziX09QH6pmwbMrZZKm3aJLdOH8xeew5D/1q/hkAx6LmaBE
ogiSNuwOnWmVIUMRdr/3sPWkT4Gmfw/ELMfByGZeZqcPu1zJlhj4C0ArzNMTYPcDtRB/Ic9F/NDM
c12TjJdlnoAvBtY/sNMzZyQ3fqcMxuPKX07tlCx02zNzIqWHVTFGJTglH+f+ryZyjhjkWBPXwoni
C74ULm8YzdQlfHF4SFVpqAUBUfGGaqOuF5tMvYnxik4Ox4qrKrAsQ6z7VG7epop51dHb4ZnXO2FN
jXiGPBzXe/Co0eQtbB66I4GsEgn2UlqhDnBidv3CqJ63xTBg5Lx4tC/cvLIGs/tJ9ZNSerOC6sxn
KM/URgVkgY4PiVPMBILQSGx4Bd2EjjT4C5655khvdH6kdnrzQF/j6dVFC129kiikKO3sMtnHu7Bi
7UOiHOWd90zTS8HE4jauEfAuNaE4V15l6SIq8Up0EBj1RviPKpDnAWLyg4rM1050nH/95eXEAHWb
82V0oh6YeedtOF9piBemXYwhUAiUk6ManMXeKXDc2EDjANO8HZ6HJV6dOcvQjGIxk2+ph/ljnXZW
qTgoAMKKBgi56/4rdTdFQVTAa4WCn7OPoF1HA9gcwAW2qkwN/8nVRpNS/HzpRt8cm+orhw0dGMVq
zW7GMcGC8bz5ob/Egdz/n6kBO2TWczBjBT0K4utDFYTURRXm2osEs2rIbR1f8XWgxSJINjCRNxUq
gZsXvOSyXVCvK0b0Rrj4hv3MUArB6oj5hX4Yl/4ZJ1ymV/yFE7RkqRWomEmm2a18VYlzHMIJupKi
xyXfC4zWxh8dib648xHcqTCXnk+X43E/+sz7ur3GlAzwCzHsXyyAihjHnaS6M8R6VOZEzH/aGTtq
oJSmH9YjGxM/m+aDyiYIta80xeNvQq1I2uPW+gg4Hb6HkoSu7hMrfiUcXzbFFqCmpH3OYzpU0fuI
TL7ui+Uk3FTOg7cuGacCdZ8y6282Z+b2mDrIfq8cGilpMwImujdHLSb2AtgXhD4jxMfnDtRHkfiL
elahGSDCZHDhPYixL0oufWJ7GHmS1iMhtMSZV50jSVcdJ8dhLOcFF1adCL/lUjwFxJPiyfaNRcu4
w7Wxipn6ZLawVVKG8AVtZUqLIeE+5qQo8KiERV6dtzbQ0Yw4hmtbIjVmKRCDZbVyVl/nzdff9mZT
t82pPFdxd3ru9KqCnxXKhdYh2b/3jTkhtmYyahVSAxQEDDVq9ZTXhWvjzXmWgemQbuBl8t886lfX
lhBmWyBRmXTdq5bUkqhBNeHtlQZGKTT0vtr8H+GuFIhtCHJ38VDrqsImMdL/Y8dx6LdXnxEvtIgx
ziM+1BhUkhZBSzD/9qbwqfyDcleRmpoaYoOC4gyggdj73sp0fw4QUTKT4/wRMI/Ay2C37P52S6zF
BmjAFdf3fJys/BRdCyNAz7nB+SeMBtyRwOiz4zaATj/zMjXU92gn3KV+Y2Y1XWX3OIH7OS9HymzH
zZs18Cg+3CeEDTO0ikUd4IOWWmHEKRMmfK37fRZscbBVrZhs0O58DBb/EkqOOgzKfavuVQ0ygcha
cejm0nwsUOdEbVJ3kJGFsxrikQkhNno/mFb2R7xz57EjGeyrbx6nowKO9abbjpqg36Q9hY+KynUI
f8YJQ9qYcyDmhsSjeHrmy7PP1ty10fOcRN8TfAKAnYT/0zgnWVGUcq+TFcI080YSqWFjM5J38bxc
41OTVmoqvT7kgl73YrL/d7uDz/fnSIqj1uDiVlct189jRTl9d+F67vJquwgE/fPtVA6/UINnlWST
p9xdbfTij37yEFbnGI+Iq/huMhyHjCdDPpUmXtpHiXBzFxX5rrnaJuYevomD2aiYLVHItR/KIcsB
cu7k9yuS9y+pDaj4SW4qj8+uFqFRd0vr1cqCzvUMdUyiXolp/R8WE4WuqXx12bR/qqQplILQ+UjD
myGUeOxq4mRFtNcDqSh3iBAWZdug+HxVTeJvNeX0WSALTzvMGh6NGtVM1U0XlO3ARh4KzYeCsmmD
DtwXbba59Pt4hK/CBASh+3WtLBUjOB1du3HasPtH5fx4nmNr4prlp3yFnIjninRZzCuyyhBtJCVO
DU/1lI5iZRfIgpJYgvxsmwJWJkyB0t1OI+xOpDLDLG3CB19dJgAy3trNeGjXMOXOb2lFPxzCjHyX
CkqhzLO0P/V+qwjS24x5C3f27D5xM9StG/L0cNjMVG8RDzlkMNpqhABlW/EPfoSlpFihKmLqcdM7
VBlTDkkTyBhg6rJurT/liqGoChA4cS+EPtjnZ9XTq7FZjDTDmPHGLP4jw2AFx1bPb4e+lTsdtQeY
X09GNy84MYY8MOPK/Lli4k6rYlFlx6IsuxQLJuuMD+Ll9SAtj789OwrMbhn2SLnPpbaPCvoGniCO
+9kJPnvfkyfDBEF1uULOnML1eoZSNfMHoyTSSqXCWaArPwV484P9I1DU26+j479J35vgPoZD04AS
MBhTdB09BW/7cG5TKb5D3HYzYR7ZJvOJxhdCfETyjI1mChxR7s+0CYcOblJTDEORSMfoSm1tEzb7
IkdQbv+rS4lqwsZZlVEisq4gqvQF0vYYvf5EbK9Wm7tQz1I/apOQVmxrDqZIJkqMbpllwgkNUKEl
xTvyRoLdcSPvXZu3C6s1NUYsLSPfYcDa0UGKs4aNom+GeCvy5Xg3aZXbJ/LBbgRZgm9Ps1XlHF6K
btk6ZJxjJRlzKYmg5LVx3iwqJA2y5RP35emhP++OtiaD64go6G7Wy48/3szaybzUHPEzOWnvP5e7
MiuyYWLDcBki/8rkb7wMitgD3N0/tHGw0bGaxmtwSL9WdZxY5QgXnHaNiImRlWSZyaNeCxWHcR3L
l5SsNKANjvZDxa3G2HbVweUxdYPBAXeRmyteY7cYlwY6eVMLn/RCcmMD55aZwoB3arB+OYhIddV/
Z6oBerLBtf28WT21UeUi+HXSjqJo6xsCC2v69GE4AL/d8XwFLqshOC8cFMfXPAAJSlfp+gqZ5Aa6
++skBqBxy1bueiZtbbCj5/EVZ9WWs7IFmlhhXUOMTwwm7vBgFVE6b0CWcL0T/HvkDpJ7WTFshKMT
LTwhPaWqFjVaaooSN69NymCEbJodriBXXbrDS8jP/h+PpuExyadozdtt38gA6PifrVdUv6u8MFWE
1BkGXKfKvfwghrWnEp5ujnaKlDfYX7Liit8sUuMI9Js/PZzEduZBavgC+ouFqhIrGFvQZE8u9PDv
nWBcjhGGvTKLjx+1g4yUsNt3/VonkoJNsvb9zqtioWVrZii/3rg90zit5Z2Ngcc3MNlfyp9fXnxZ
gKlvg7g7M7lTAB5CFvxWAc1GCO22aNubcMs9rvHcTGEUGHJTw0Sc7NXnqyTnME/q6Bj1PYzeqCGS
v/IDLnEhPWUlJkIXYkJPLUuogh4duWarW9BfidOwyc9+S5i+oQ0y63ioYe8ccTu8X2iiQ/DSpln2
7E+SaG47uBEKVq/2pgCHrQ19EmKyivhHnr3z7s7OB320x3oRKoAclskRzAeMfjmYqkQfbSrRQ9YM
K4SB0B/LvuSPQpnXjfR1cV3bMZ9p9W+ttzd3XLfOBp1T12h4AkFkJODzuUGftLkvUJscEeSXLh1U
ECvGjYc6b0LlLTCl8NhQFgDJS7LGJMRdSnJ1xdWlWIszc3nb+/wAaEPahn0PYTHmMNvqj8uNiG8T
Ua9SxeSsdnm45WT7Bwd3wpEmWt1BkB+74Y5Rjg/PkzWVUKPGveYrIuM3TREfVgy9N9u/xbYErz8Z
jPH0I2SV2jYWPHI+BkEPTW8ajKZACem0g2NQE/N2+GOnxHCCx+32seoGQsr3+TCNacYR6PrGsSLS
sonKC49bQYa+D8nCEWIitW8Jl6gKKZCDmAcjuYo6TAtG37mEqOHdaqZb8vfJNW1lFvEADL9Lkjc9
L6Jg5dCFYL6ADJi3T2CTSlf1tWJVuLBpEDJrO+Lo8/u2e/PXbPHsJq72WedLDosRLs8vXE9m5Gzb
HqnM3+QVXUrQOs4GCEt50mEJU2xnd/VPXhpb3HJvN5lZYKUu+Rsx6QZRQzZaakNoLideD0kC5S4m
mR6XeqkxuIcJf+9X9ryvapWMh/F/TDmk6FS225LoGgT2sK1fp9S/OPUb9fNiJBZj2F3Ji7mTzoi6
H7bL8wMC/GQ5FGr9LLZDHUxzfQ3pBTd0wk+er4Gj3d91aA3h9kkv9fGgc3QcUgp6DRbfBtMg09oE
oACba31DWiGjFJoLb4m+JZxVXSrDyIn0Ob/qCQ5sR/fRh0dgs2qK5eXMHocCNMjuOSX+L9f/Cg8n
6OvJPtKvH/hajsZo8XRJXKuA6UhU9cLbqzvlejiKLaKuxADiziaD8vB7AO210+8DQMaXC00cnw7a
2rDTzj/uQgsRCgj746NuG8OrTaB2qXMBF2cEV7C4GZMG54iym6Nt3kiHiyWuru0V/BlPmR2QtbMQ
YYyxbX2hizrKsNy1g+nq4EmVK0Be7Tka/cASbb9TC/832UMaKe831gNBndEhi5wmgUUCNcA+xz03
ek64sRsWMcagVdbVqbzjj6/K4imAfWRnCdPqgHjTUDFOM3Nl/WpQGy7SB8YURE7bq7I4OgP/mLPK
IE2y58c9Fsi4V972XEdJK1fIUIVg5zf2966ldt5gd+mVmhrfJFhmfCAhDy4l1PV7FibNF1mSTrdp
tMFINOcRiZYw1QUXsB6eZoSfAi5UH7mvm98Lqp6tZN6qdTElpHhN1z4V97nNExe6PerMURG2I2AK
HEnU4eJ/XqjnqE0tY7WNY01D8Vr6lAVLsUG+pAHj+Iig+gJkAZ0E2j3+Bz+rU4YaKcQn9K/mwGVw
Rw/HGgKyUDeSM4kT10CYijNMiL9dHGgL2k1dwxTiuj8mgTv3YgqSU75IaqtYkw2yWDVYfnuqntXl
KvhVYDFOldjHQ7cucOBEhzbPTVZrdYTq6Nt6xQCd0OeQAZHsRS4of6bD4383f9xSapzXsKYMpjI4
jpHb0z4Enz2HAX7ADjrf6BgaRPwIG7VWBeRgW4djsxy0L/dWHU1oAdhpFy9URv/oATU+l27rJN3R
kXLQpZovNE0aWhp/zFTOfF9ShvmXE4BbqMfhRQOIaUDplHIODvrib+Ry94T9wB2jdVN5voa+sGwX
El2/HBJBo6hTdMtSL/9Jq9GhiCpgZnLP/N+ApJvbSt17RirZkMRfbyVeFHVFcM4p873JDSKELOai
vzGdIc4bnRnx7JH6SvcYWys83z8Sr3+f+LBkOEnEoOxSBbsAredjf9obipxtvIf0rhbk9H+vr+7r
EiGXAmACys2/7sS8/jmChi5s4e8NQmzAihs7FIVO0uKx78UxJKJZLhBLOX4wxdsYN1a7vJFIxVpK
sENGwaFRl51ArH4J4/jdELGNfNUF96o91ZrlP5jhcM/rKNf3h2kiCS8GM0GRrLIY0SqyI3FBJhdW
mzfmg201UUxDA8K6AEpdNKHiXBEYq3eQqqj5rioY+ti6fIlYDlcWmHsZ33BVlUwkCy+PXLltv0vR
M7yyNbZtZqvjixMM2AA8BWb12VGtdtW4hWMRXsuXDLtrI9PYSSx0yVLkmuH7dO8w10DEbxxVXKoR
cDZHYhOxrRokjSjFGx0UGCTQBVq8gqtvk0itgN0h0PUdnQt6HEhJROyTCw4xONm2/TOaXCfUoMJF
UdP/TMICNG4exXHRFkx+IT23eSHmNzeWM3Kt7+86GBa5opgEKxIxSoHp/weo8SbXrKp0w69fjcbA
xYRKyWk+ooElRrpAUZu2Tf6Fy8CsHE/j2l9IRo9EIjvh8wZuYSuYFvU58gSlRt2lTdb1ndG7RmYa
mRVJ1YGdFpT+s7bQrCpgZZATT3SMJ9Utuhgzq4Eo5ux7ma0bsC1tNIvgLsZ19rWi05CPgDuNvxzw
ETFjb9CEE6j247mph75Wkw9x1X/oUwtVmpF4kF1gm4niZ63l6vCZXUEU1vALqsGov/vrYUQG2US2
S4p75vDO5TBcLJnGarqpoBM59jCLqEwcsxVJMnRbws/yGPwpybXl7JgorKDCvr/ptRDeMnViq0TS
7hfqfnWuozVScJTaIhb8ytUz8TXbFpotFxD9OvT/TcECTvULZx7A5E+3I2Wzgx+C6uQ90/Y2gz7p
PYIeuhtPw+Dtv2XnMr7E2mKI3W6nE/7aO5ak8y4XANGAUSUNJF8Cxfy3kwgK36TqMGJFMoNtNN8v
J+ZdQbP3kbDqq8Eve6eESbLATmqFun5bDmRgJo+E45UBlyfO0UAWmKYhPevvCjR04TghET/DKDdd
mkZh+FyO/glionH/OR2xQ1aWAAJen+5XSmhY2q0oe3KtV3U7AfX6jKvorbjvmXdeG53arvSwARAC
OnOW0iFyTMC2h0XVivz3NhO/N8+bO/ox1kyVLOuQn1aRFJ/nV3SudDnlPve6Bs1eJPuokcBvtwJB
RNwcsMJlmDKCj/HckNfx0d8+bvZXv+oLXAweHaB2slLk7IlHsyC5WXG0COL6rFE6CNgg/EoUvEb9
KwfJ5tXfpu//foGzFuQPZ3n92mq7pUrKuo/+dgqcYJq3eFxRB9wiYJXKN0XTu+JM6KNQlXhVlcHw
tUQSHP0ZikgLDNvf+2MyqTy407PGZ4QialTeGl3iQOZUzVB0SPWBtLHUw7sRe89PTkFeJM/nvuod
XpdBShm7P7gc5tQIt9UC1RSVVQRLjp5GH50iz653pxywk9g181t3HlQPMiCfvMBUdMZV3GizB17J
pj3rL+nYsbK6CHCcRU2lMnHVVGb+WT441LpLuQpn6+WfPOfWCIC5oKYnOLJ6CPE08rWRkOJ76rvq
8H1MxyV2hVdGRldqOyM0oRLowlm6uoC2iLDpyDJOmArOnXnU1LRKhp6XLkBztWEIODmlb5RRz9q5
hYCjVJD89Wc1sHqVsIud5M08x3ceb51gwtn5q/zjaOxXJOyviLIPC7iCMABrRU/wZRHjjEOOeOma
0jPrjEmBvcckDBst9GGzn5Hen+oYdln1PB5v6kuaSoTpVixQ5RXIjzmK5Rnp+ZSwFiV9NV3VdJxm
TNEPxFuf/B/FVJWdPkFUwagIOcnx7h6sby62UWg1+QNACuvntysm8HDfIGcesbVrdD0GVyyiUlT9
qujTZd5fN3DX7hBtLJW5HdRkhkCElGuAjFTA32Rgqoq/l/HGUdU045nAasi9Je/Fpcj6LyFY7NB4
fzcy6QKMYzLrveFAa1CJoOrlSPrBvZ9Pzws22qAdbldzMIOgiDg1hFWJNBGFhdBMfyxuAc6CkGdo
QEZk6POFdfWEJUB18MNyBOIP7UuRQoXo4Yy8EL3z2BsgkaFB+3DbgNSKy2n4KOsM6x/4pgAVhpWm
N4nkwcEJFHwJRbjYaPvwBH2orP7dO2at54Rd+KyloCsVNHRAVdzoKUZXWilczwaz/yoQ4MqylNcA
h2ylavwqVlmuFczn9PoipoKjUvYkGiKPhxD9hDebG7oG56v6mz/ZZ7ALvJueV22K0G/jP3Xq6aM1
jJvQkkB2bfTkHf9XBqDiglb/sMIQ/1AyBo51o8LdDoUU5x9XtKQ/gQpcPy0LR+EPPqZX9hFtXsjQ
HNNdCogV39zxybmvpeXIPwqmYWEU+FBZYENSBw7Dg2cFdvyr8ZdLzwUMhYvBKDPoxiaa85lS9YMs
om42AMCGWcbV/JWzTm4FAhxgYbpfDS/naeru4+9kos9iF3osPtFszkhjLWOU6vf7Iz0Wj5adQRmf
Ddpkuindm8g53NCrNHfpEcuWvI6L0HAxNdycJ9FYgpkC7+1kDSGBvbJELyuFSvd31kNPpxdXC0Zf
8oGT1/3ChbnPj1LW84P0CsIz9lOsCH3thbWxEKoxJ67y0gceOXA1WsQKDwGi6tKwCY1bzSlqIwNW
enoWEABtqeVUQLI9O0hQrSk25ZZEPnEAt40Ab6GK8nIqIx4+YL++spybtEaePRUwIe2DcwU5g7kU
whdxfqR9NpSuFAC2KA7Smzfz1tdxLjFgefcQ4NHmHbp5h5PiGH1bHMj3LIMB1bNPE20oXcDKcKzw
wlSRDE8vDGaE6G38Keu86cZGLXBeT/y146/iG3MB9rKkGrXLFI1iVLTnh8oFmXFrEXSGIAKEAf8c
4xtR+PdDJqCiQ2jQ/azgikFlsCtZr9hzF/abUiCPqCg9BVCoFNWPmLDBGzQKcwPr9yYFLs8WC4Ar
AjIPmX5FfvfF7+vXg7VV4ysz2S1+Zxf9vXxh17Him7hKJW9LJWB3IkmMYHv++QbQdGKGWzjkCVcv
szpLgu8wa4CGc5LUkGl9tCdt2lv5tyi07YGzohyIoL+8vbZ2M1jBSPBHvNhJu+A41kv9MfQFdYVu
U615hug5yYk/zt0ZtqOoKvW4NzKjsnCWLev/yOTeZugBdohseCEceaoSvJQn3vWCFQ4yQ1vLxKWX
Z5ryG+BPeQUTo/4pc1iGSFc/vTlpGh72MYGjB/TjISulvo0QGMmx5RScXuMDWHVTaSyxsom3KSLH
vQwplW6DeVtoUcc9GDkZubmDaA/9tU1CSiKTc0smVpQWMNcEjxMml6rUS5V+0z7/V3EX+zVI6HP0
DStP9Snm2vfqUlP/rjkoYKcSB4cjjWicwfCG8ArK0oPBxUZu/dI0s+zNUTTVanS8SJNvdJOD2tdq
PYgmawbpkJN/KpQqp8sdM3nHq4mqpdsbaerp5ZjenuqEL0kctNGxpjL1AaGgD16nlDPXAVp4Vl5r
uf4KY7vVAQcBCrGDbw8iHD6gzND1a3rw5rWgE3qOMvr+mnjB4DisIajJLMVOXCr9T/OhO4pgbWSd
krW4BRm7oFpBdfEovFfbZCLQ4AvZUp0NEom+2gAQKI2nj0x+GBJDEbB7YkQY1LrIVxho083v/jTK
A8E5rPPidr85A+pYI8A3yUTvmLdXqVdxeRL1IGO+RjrufiyD3jy0dhzAe1b1nQBIBnzm7BCZ3ufd
gkzYpK91LYJizYjK+4eC5mMXPkYGdfbLyOGJeeSU0OBSyj8OncWnSUnyO5v/k9Bqkr5rwE5FUirr
tuXgECRsyE8Ibm3ZbsfqtwB/9mfMg9RVWe0xjXuWntznzBclOqtqTsbb62Qotd5jleLyhaibRowm
+RJDhDHzvLfDduw3kmxkaARZW33uQDX/nowwTvW8gTP6d52EnekSu5ZilzP9phRZQFeMASUzw6/o
fEY1OLdvpqGCiIRsMsFdJmYvNP89CJU0GRWrLWfSWBaxcxZhjcMW+EA8v7pI5CdPZ5uSgbgQ4qDs
TR0x4U/gpNwa2C024fPXulG5AwbGQs4RZgMg9Zt2yOUJkLfxcKHImP7CtSwwBUctQ/Ge++KoPc+8
jEGRtanRLAyzEvBUVRVArPfYECQymFlnM6EZUrtd4xFhYepWIqc4okGmOLHxOHCwMGpIjdP9E128
bWiCPvlxHYS5c2Z+eq4JC+YvbC2L+xHnL2bTOpaXnm/vPSdbkuYSD4JwDLgJ2e8FjdPlNnaqG4Pr
Gw+flRhstdCY2Pz4T0pV1Y5hGMFhYEPIBnayvjirESTftCbi/j85vbRBgSdGgV1v8Tjh+7YH0zDK
/TacdRPJcbomRtInhh5pOCK+gDxyNzCTTeGRYcgjzbqkMQuqdx6DY5nC8JHV7QvMulFV781ciwAT
807mfzUJfm5fDddPWZBSGl5rl77aho5VLzOEbIh7sOhlSQV7AZI6Cw/RVCvgGnkowpkQJnixkqfE
0qADKz7Al28f46ZgJBm/BPuidkVXuyP+A+Gcwqd2d0zQKEjXLsxY6EVxqEfRtHykBz0bF0yUetX/
OD+fMchSRChgrw7Z9uqsCv3ao5NF8i8Pmg3inwTI9GNmv3YCup4DFMBKwmCcX8w/XL7XtUR4lryh
HAhJWSae8T0LWmCqU3qwZWGWFJjQYz3XHd/LzWNtfznHp2/em0lfZlT8KFg613eFnZmdhMnO2ALD
FIeYeIeFqTRjUsplaE6RX4FEt0hLMgSJq6HUuDJfEknLsTno8pXAL2nXZQp3EbTl9XSzheNmfbQn
fN+DD8wGJyC+D68nZPoOYBt0PWV+lcmm7mUEMK+CuvXexaN++UV5l8vFKyp4np3AuHPMqjGkRJob
GoZPAWhuIj3gA+kDVcNGMTWXh2smyb7uMikSi6UGtOaZVmY5JUO074v1o2rwqhsmI6Ij0pzE0itd
KNEzdFptZXT/VVsJrEn0Qisxy+2zd4aSofhytbEMv3v6nXJRTf4yz7rW4uah0wPo7cEyVftU8y6p
Telv9Hff6YLru98rJXK14uCY1qJM6MU5TI3qMoNFdJf4MmRx1gDksZofw6L0N8qOeRInhr9AZury
oxyMfpEp0xt5MFiuk9Gn6OYM929DMfozoVYcSl3an4felu3nFyL2N44N6dnle+hcRnc4mIqRSyEm
AFOc46VcLziTHuuZELlov/90R/7qcQMCQAoynmLnK22dILg4Khznr0uRrVTEvxw69UTwO3QWWHHa
FPnsn1FW5o5ALPDO6UKB7unB0ZMoypLohuGIbZJAIZUD2FORc3CMGY5l4gFRiKEb6uu4F9armQ71
JsD2zWQW+TqbMmqZ9hIGaHsYisV0qrkDQXC7ZLYTDc8yJTj46cdo+Hr/kDhMAYZ9ophqBmVWou4K
UG/kd0UomV1/sorc+hkCWmyFaBUW3NGfedyCJQxA3/ZV4LVMKLxa5nzwAXGKJEOcmgvztDurY+hd
+4paS5YdZeRoxgX/botER957QVrvIXKyQGMTtS3KqhWxC645ox0FCiYFTDT1K/atAkP6nQ5IyEs9
pASaCfD3TzaFPDBFeIiRd3Jk4e5ivzMM7pwUmxEVWmq04jhI+6/DseM49VPKBrKtwtn1chmlVbRB
trh/9/NVxUYaGAjn3y+k0M2wiknxjRI+6MkteztwYetULaMq1y6IGxQ5HezPZzhwqRLpFl9zkVxV
h20prBjMYglWuoOrsSK7HH5CuSMbciIkNpTaCM4rOSyOzYzisdHQNJ/wyoPMAY2xfi8nJw4vV03k
jT1y+G9B9uN/x9nkOl5q2A0QQn7h+x9nuTM/FmD+2JWaw1t4bNfaC/V3+8MVDuv3Ahyiq78nbqDX
p2VrJZexr+JB9458D6EyEjQWZzB39dxJpD18DkuTyRIVgjH2EyXJpHt1hSb/mg8u1K1PSOAYJuls
vaqLSnoU15+robhU0uOAjZwKn+zAQ4wKP0C4gzx6HSQ8o2w2mSlPgfw0BghAjf0hON7sr6brS31J
oUTEW59Y0zYLGfJ27twROICW+zFeip5UQ9P3iM/+5tv9gn6v8qg+PvzJJUalJ68YW/CZIyvEKy8Q
JlpVQFyBZiF7I6TR8zy9kbJXKXBbNiF7RccPrlbWOnSTgxft8o+HV2J8ZGjx/InaHS+y6lkNSb5E
IO2DWW7EnTgfxDz1Jf7dmSW/epJR2f2RXj86GCMa/YcyQOQLOe1LCz8Px8xnJtQkVRI+cNF0zj0l
S52G2qKjW6WxeGREcfTvMUBr21AkZ4Ta007yCysE0kJC7m6RBJtEkD6QuO14T8x+K1qO8/LyKPtz
X+1uYpp/s5rwictM1/5lTZLTQcJ2VRYqojiK2bVEM6YTF7JzbzhWgRAynJhbyLifUV3yzVi93kQj
hCJB0dDue0vCRP5kQ4PNjDnVbCCOVphmpZo9FqNCJZsrF4IEPkSnl7w2EBtP3wj5TzBdeqixH+lJ
tcMrz7WUxwAOtfUybARZeYeENzKaGdfXKZi4eM6zOVuupQp2sr7MMG+TKz7tGKlNuXDVe6i+Xa6a
Jb2+37UKrjov/Ijezpu22uj9xe+9KSYjOblq20JAuQJQDm7KGkLwyPDCg36slO+A4ggFqyGfg9PZ
e8GwH+1LuyhLSbxXtDFgUKVHXZ6GPhBrvwCnOY6bx5oPuFFZsarFy0KwWHScXzC6P4+7d7tUUadk
i4eJ6Zb8PUF1oAd/s/OK/EKNEp9dLri2G6RcYJK0OwHr7OJAZAatCRnwyE6aMtNmoFpgueWQIIvF
Sw5wIsYjtP7v1EUaXixEF6bkC9U6TTX/9LOnxWkauDjkQz8eZ0zvwKRnsKCA4p8+6LVuQLLjqRoH
nMdLuszVt62Qek+bLdH6SruIx3/WJboBY4tBW693IhuLUlBa8oM9wl/mIVdN4Xs/lO9XO+eo2JsV
0+xECHW8zRIJptLR7wIoewdY4ENjTIacllrp9J0l8raImSnyxmmJRzNGvVHXcGqR0i7p2IRR6b+d
yqnm3PUyirDxqatuVN/LNKTTc5oorXD0SJFUos0UAG9dBBH5ODtES9Vp2UB+vytgloGUkTBravUo
CVTmsyKtevDbQ1dPwq9d0GPRALRTQ8YCJdq+GaXqRZpg7wYQos9jJ+5/eceEzzL2NUGSj+wteX1b
y0dcjKAo1EI+EJvVn4LnEeXO4XJjvTF0h4ECd4DuC4SMFDNa3a6N4d6xlhquBLcXQDdwng6DwtSs
BCco4iF1GQvFZYHyAtBHX4i7SbLhIdB6WmPOnSoVI4P88p2EpuKT0MKakFK4jO1Q7Ve4/6qssK7T
PfOVnjJihzAGVQlbXo1VH6YoW6fz+ylxRNa0AL1FgxNQyNIszqDPi0889wGo78RIDjZBw/u4e4gP
wFQqyu8HzIhMSj0L61q81yY2eZVKPbGrypzpDjoAg+S+5S35/rl2eL3CRQVVwbquGaMEDZbxMZlM
L+y/m94u60xlNwFc+lPk9qT4yhAz42J/3/OcVnSi2EvKuMTlU/QJWdwistIk2p7m7g2dsCDIXdG7
gN3vnZveDEppFqNMh6ldoBFnTCDKwmpGj76kA0B1uR1ueisFLlYT3pnUaMNoGvHI8vYUlzEnPpt2
emt2ujEJs7DNpQ4cejWToLxhoaj81u7Fe1P7TXkI9Q4C3dZSnBmYA/W7NFdG9M7Kztr4GTLiWVTm
hG4m009uj4oOELIW8++Q3aLkQjaXM4QWwbDqQ0bzK4oSEoGZcnxrBmv+maP+xX1t5YyKS5LybQGv
BqXBhX+jGy0QWJiLFqZnlTN3Y8E+lJP+jAg3EblQIWXn/UqZFDIiGO5YVd72RLTyoVx66HyYCVSv
Vk5sVcBLulqoNsigVJvN13saUc75Lxv/tuYzBHlyjsX2w1KcEgDjz640YuogXnysPWDJ/ZbpzCr3
MSPtcFBac+vXafX6xA4njrFr7xNph/M6tmEIbaZTbUgNL/ox61SlffECZdom/XLvX/86mwyySQbV
umVY2mBHuz/jh12E+xzSzORh3/+JcClZXlwx2zOf/jHbEDfoDfJZ9dseD2XTmlqnsBdP6d7wfD9L
yM3+NT2ji3VMHbH3PCoqYGThWC+jhODpMLnlnxsZCovqtK8QqumD0p5tzS1m9ABpTpWQHwSQBxpz
uoX585IIgWNToR8eyQuGaNV80VTPtqUWaRIbV6tvCtf5iy4KepCxQPNtldY795/7M8LpYnR4izMo
3Uy3VVKx1nVmWUUuxMY7+JTpkRty/NgJa/jnQuURLB8h3zT7WQOwM3WgBt0yOWBWS5ooI7R/jYDG
aHAtgT8SCdZdWWgquGi3rcXdGwM1CW4L6esNFnxed408EWpbPmnAz+tr3XNBFXpgxSCDK3Nwwqsn
8LoYhDJsIiAOaUGbHhNMAqRM3tQkZmBDCl3PomkUfYv6h0iWxZvqk6Gk8IRWhAnw0Z1vEBgMiZ9K
XdMqzJC/paK3sfBWKHD7aKUbK/u7k2OPENLT8gBK6qCm3Twmr1NeiDV9a9IYL0hoDGIsZa0Y5a96
7unqzovCaVTPLLKdmiJlGajyxXfvPTtFeV7/rbOPAqQ6eFAnEREzmcPnIeXkr7XLE+NXZv5c2w7i
JiJcS8sO0/JvhrJpL/F4T8/6wGz3qy9KwI8MwYkfFUaA7m+TPCMWP644NirjWKZ+ZIgRhZjpTQVa
bIxrkLQWq8XalVR3CalNpAI710JsXlpHUQHtIaURHW6O8DwRkSImYUV4cjs6cM44jeQ2S6XXsWXP
vfFBm90t2kxDlf6x+x8AuSzppLXCljsknH6uYBhpHepl/bVAGO2tTcy74amAh5nFgwWw63cZnj6t
r1e5i8k0APgbsaM5WqJMvx3ErMSp8zcyjZ7K1DOqxXTRihJRsRQjjox0hrmFwBS+loHfAOPlqLni
cP6ZEPj4Tr2d3VU6yeMebDxRrvm71iqh2qmyxBEgGEO0L/qE0BRhw206zlsbuwHKahHYw2VRCQO3
kzoiMb4mRg/0qiYiBh7vlP2D0jwXG6nLFcRF1ZG3VBq8pqtTxbI220z9+xhGHzCy2vrAa879m6Lm
DLi1XH6QXtNcgsgWT+Tl91U4hizQWLnsB5t97+nkmltAEysmok1SV90nn7QQI7xNBC8JCfkwcTDn
QsPZEsKJ1O7Q3YNIYJPgy2GEIZBTcsxtcseLzMKT0E5XhK9n201jin611SxaI9VxD1BaGAsrh1AL
90HhiQnfNzqrNO5RmpXL+AIDik/cQZyA4zPIo3ImNsX5Mw5fKcRyxcmYWMrh34lVrtPgfSsgXKBO
uYJ2VSoJvtEkAycSt3SQxbdcJz87huFVdsSAH+lDMxflJQudPuCfB7QMoSAH7pNsxUWMLfmkxEQy
jUTDdL6MvNxmVP/LDn+KRDUMnOgA7WaN6grh9UGldsJ0p/u+XDO83V9PHQNtZ7YPmaVwVSM7wU0H
VxYwhZC9w8pfRQcMumuFxQx0hYSVpExIY2unvchW6lgE/TQ92NQJN2bmMpUdMRkyw5wc/e/KOulE
zlnQ9DbYtf9zqLrWafNi6AO7tVmkfMKf4GjXY2BSKYVpQjcscdqw1EYqjfoFnpAr4TKfIJXnX3xS
CxmCjJoJ74XH9gj3GITT5btgpN1UbW9mG+kZHyF4OQ3buvuDMCoPyY7Mn/aZP0BYl+mTnRREL1pq
TCVJLY633Ulvx+wETKVlgv0aEP1AkvJ1WIMytlNpgj4n7+gL0zgfuGpqLFhbNDrTq1Q0xtJKE7Lr
mGdYQRdg+4EU1P1vNvlZiqh2i9U+MdQyQHRqBvw17tc8YtPeRwXQEAVmMIg+GnxyoPFQjCv7Q/jJ
Zwgung/14tlYIfj/i+yYOsZ5pLjftRvK0s+DR91m3+WUbojb3Mt7sdYSXoA7IenmEZsRc9R9iK0n
oaWO9k058shLuq9eUzZJ2qlaba/5FybhF8/lqELKRGUTx1yPC826v0fRYquSHtOpgnGmTKU/LCuH
vXpjVSycWE5LNEceGs1aF2lkcZMq5TWpc3MsSWJeTY2KxLv3N9zRw5i+9gS1m9DGpl09itfylWrK
LALQIsJlzuPtqfzQpekPttB91fGI8SVCfomTsicBBxsfMfOv1wtYfFrbeTN3su4GmA8L+UTEmY/h
jH+TrhZPalQcoKUTQCzXgVBXWeNy+E3jQ1jY+V6DFi9UVX/JAv0BjANGe05OKJ+NCWadhoXRmDfo
l18ZQfo6+dYwArJs9e9pJDJPWyEOkUmh5QDGIiJq6DqAalRtNLnAYoWnJM3acIXPogm7xEABHVTF
vZ8UBoPTsSnJ9b6dxiBNzcf1VC6EwwkqI5C+fERdcNNo74HUVOOnWx6bE4Whw3o2yfcCDhlvJf/R
b79iULVQPLpjew3BQ2FJe5mY8h60rjNIJ2pQ1YpP3vvoJvQAqZC/trQjuAoG9YTsLivpT+T8nuVj
SjDHXNaPLYyA6d9we+AACH8m6KwD0+V7a0JD1/7eV1CynjgJzxqipeOmLylkG5Hkontg1+mUAPxK
PP5q9pjXIhBV599PVxJ2tsIV8E+IWuTVGMvh3dhe8xdKqmy61ANfYrjkQ5qMHDffOjkQNccofS5h
bNdub2VY5Cek0TaPs5RUhUovOmNPgIElu3ixnxLe5PtDIN5foCNKkT1ouGnuMcb/gVyfaxcQqNPc
D3PZIv6eCoMfuYcJPV0fJPTdyJ9KnA39DZF4/a4dVI74egnuP7xrn3OUJ1UmBorpQVXLkusI4yoB
U+5CZBtxqcYx/431s0RmYhdtONZXj7G7xeNqy/4L5j3yCBY+ujBR8Fqu0wyDKfZU/+JM2M5bQMY+
pALqEOR/inHZfTHX+NXix5VRoZQ//F/Fn48FGwxZNX9bwFpy8OuRjJq9+lt532X3X5vF4JMHKTbZ
CQ14kxEd+3pfJjXArJNmGAnKBD2ddRqxOW6VQ30xYwtzn1CWmt2GYVNOMac43ithOal8QQbTzDmB
ajUPg5MCMfP4ypIEPComtjqRnYYU8GD0XCexbSbOxqJE0bGGblZXro0fU9kNFuVv/NJ1ontM09ap
lmbUdqjsNno8eKBk2aJqhwAZW9rXNrQxKy4473TVKPJlRjBxgk3IhIWwrXCo7V5sV3jL7CZ/gC/0
guNx7Nl6+USdCf9PyqvnEr50krow2Dnt43R9JnaqppDXzoAyuUB7WJ5NKgNdUEDmQmrY/9v+SLiE
jIgspMtCZhUhv5Xi6Ri4nDopQj0NJN9INf/zpM3U/+tTdvZfQjC2MCV3OgFSG30avFwqevcVec5r
rzxkew3OiYAdzdyn3rY6Rz90qCaJVTX+7j7BxDPx8aC4qU/OQn5fXAwregdOK6rdydxPICO95tgO
uhi3c4lLCf4jbiHv+ZR6vHOZ5cTlBGemSaFwbz4BE7VDkrr6zvSs+CwPZQOAldnkMrNT+/xX0jiZ
mM37KSMCOsp6oHvaW+NErE5528RBGGLnVrLFvCToGz4B8WpWNkg21dqzozRDJeV97gqZmltxFdng
HluDYGq46SuKC9Y0bDSghefB4ZdP+a5CGrc2rT6iZ8Kr81KR2aJw3quY71YjP2XEXo84KyXHWQ8u
eQ7AScuU47A07mcdgha7HoAGTYYcL3Kc1Te1igFO8OEpYqv8I3cX8kvPAkXBzHiYIH0sw2EXWY8O
7lWW3SzMJzf65JpE9PxptviyaYKjyqR+bWdkjGcQEanswIccvjtCCkGBlt3SK9yteT4MgRuYa5cd
AE/psQ1JnlV1hIcOpkRpEFwruxCCIGdgN1Sh2Mpu7UdqjXZ7/IOEP1J0O8YgM1OafzwOuOrhwWoT
4BnprVtVGFtJa7qmzT733SnRYv969xMG1pHY8DphMzT0JyKpWhGBlSvyXUAkTe3xvjsv9zRyT1jZ
QF2wmV49N/bk9Ww+3MLF5f7bK5Sv8BRmi9t98wSd00O9IsGdpnSNeJcvZy4/0RFFPSFDhoJOnUZA
HXTXxi9URJ0sepw6fcpHqYvlnCZdjwrwPuY8DjA4R5HDEkwqxuJqBi+hPZbWWBtwAR8D5R/Jtw0A
xjzQGo3HQ1VZFnwOMwfAiij1A3VnSaamv9hr5iKLm3BKBJkSuhKrebvUTJQ8Q0L73V4qIWDRJnfl
GdhSuY3FbyQTLI7iI8lSbpn8lMvef1YCeCR/8f5HvRsM2YhtoetEpZi2aB1cOfQTm/FZoe7QoszO
kG2LqxoaKxYZP1LNZKeiE5M9Ha381V+ilKHDNMkEXynbj7r7eGXIrrF80x4y4WYoaWN8h9Zt4oE5
z0XD38XUxQtAYR1prlvN+w+vZRT5g9eAxduUv/8xskBM3wZZe4OuHIpKkMc9TAzbUbkavy+N1/q8
TV03z43JRmCUa3yjQN31U/7OsuPH24ezp4l/TZPEeOBGXQ/2LUx6yNLZzcTOyPUecL+4UVk+2deg
tqzIROfFVBvc01C+AEVd82u4vU2XtbVKF14Nmv9I0aWj1C9ceN73O2hJhcim59DuDL3zjlmU0Nh0
rAF7qsccvs5zklzaX+j7xvYoQWrjPVO3uIBjjQA0IKqkk6/ZNU0rhr3LbQXGxX7deQc+22LA8P2y
oo+sjiKxR5BRflicZxi8xjS7nMLZE58nwIrFp2vSvMryuC/AV1WZhiaTDcQk0vqFWPPY2G/ewgx0
GpgqMHzlw9AKaqttSP/rPNzHnS7AfFAXKYF2/P9Q37nX/K6tV5dq7pR/UAGLvyBKz6xqmJ1p5ADC
Du/9UyRArxQNa+oFvGLwrvOaugKcccb4YsZFtxc6yPA+CBHnodCxw/LfKHwq5Cq26kSalBDVmGJc
bIsA+LLHZb1toVVMJ6wgZ6gr5AEpOLG8n3KHUEtdiJ0XnyVG+JSQkFMF2MGUKDwKg+gu0N8tNpyI
tlhY6pX/hR/x3sHzASe3Wm8eNBaiRzjiPcI/3NYVULE2U8MHaJQArELeCQzZAU83LOXb9+VcHGFu
5jJHwnpaqVKjZRB791K3vuj43IdxzsvIalhDwUhOEGaEFtVCcj+5hsib9/4rhnm0HkRGFxpRQaKI
UluvlgIZqMLa0k/dw+AFoD/Bo5Xuqk6SEaODq+qEaawAxo1oJPqwQeq9eTqDmL1D8b3X2nnjnRNk
NpLdhY8PEY27q8ekx5aI84J3evQPKkM3arXmuEnpAw+6yO2jUyaJSSs6okMM68lNPUXZdR+x7WoI
HuPt4F5lKWotBY3L5DZ1s3CDTBoTmoXZa1uYFVgeT2vZST2uie+vhm16QVVDWiB9y5sQDKor5v7j
j3YWoim9VlpeDEBX6yj0uuW0Y5OGfUZM+TDdJHhjOntMkD5h5e1149Nj9yY2SzdKjIqqGdi0D/2K
ysUYOlXvo7/XO3a4vIWRMPAlqhLwkjf1+I2ObyA/qg/NY6LxhfvweKXuhD9WgdvzZxO3WWuJ3792
xOK09jLUg3NulHCoAHqbCSU1QH6m1frd+8eE5NsRdlTcFy0rJ0U6x74aFDmtzklJ/JkLmb3uegU9
90saeGMm/JyNBDfH4s+ACw0HUer+vxfII0m6ZaurALzCLXI9KRS9AJFejf5+IGth3X6209f+VjEz
xSKA+4zZMSQC4Gqgk8yBjz+KmWDazysVZjHJEUJJbm81ydK8qb8lsD9a5rriJAI9Ltb57BwNNiwD
amd3EAnuw+7qSxdZnbq6jCHSPTllulxq4F/UbZ012bPwwnFsej5P8weXPe18n8pafubuE31ha9FY
yZQGmSsZAAV6wfQnWAN6p3q01ew4+Y0F/DIs+aqY3ZbS3JYf126h09ZLfvkEIxHOMLgUEwLF+AKa
IXNjPq0FylVNU9XOilky+6Q0WdXaufeaH8SJqd8HZzYL2SzHCki/4Ph0pmKHj9NpjIvtDN+Fa1i5
qt59U4bzwWk2onx9qLTRWtkIf6xARvL1s0T5ukY21JvrUFSC5YfYatcq6R5bxBhYv8bl+VBBvuNK
GMVC14T9kB25vw0gT8jI3iOo2VWhwf91baa2OONLqRNMWRar4zEHh5NW6rrqvS4eykBh/hZ5ldr0
QD63Y3YecDpNKkuJnU2QvfKXzxcoEKppb0MNM2eB+TiXavDJ02rS05l49YZMzgFLRor5Wnib6qai
yQdPN4qVctELCwHnyaQDAIlu+XDPP6sv1sFutiatTjnc2lwdmf0Pl6fx5gjdbPTaf3hkKyJQe4Lf
zTkmTY/0vwiPbwapYGD8H8SIu29qGasF4EBAjrY/QiM8pdXwH0VWkpEA1/yfUGb3Cb4x5uV7EIAh
A8FplZHk5PNsTzb3e3cFAXDNX6zKDtllA5mZiY46qDCMvc4fGZ3Jdxkv5TauLi6BE3CJpjA/ogMc
y0hUXicZ6Pa23qPx5cfyjehWB2ozVx6ZeAOGUMB4Pt14MDc2FXrTAdL/+T61zXJsU4X7uSIkv9YQ
NYrmiLAlZg3ndNMcq+7znnoW3vybi4GSNVlO5aUtY58sMfDZxj6lYFvHEOs4pJjni2zwVv9rFc3Z
emR4pBU6pia/qrpY2rREMjKh/b4xqtlYA99NEZJkBWaXPAdaVIznZUg1c0SSdS0T+SRVDo0CkrU5
/AWTbmJ6b/CHVeQ9zJysk61un86gS6mFv8wSfv6I8mCZhDI1FvCeeW80j1PvXqCHYVI8Njxi6cvd
UQmfEQTbuXOFsLGp8IGBc/6Yo9chCQYHEfqJdgQbuK2/4wPyByzXuCLFPdLYK+RnNLUfm/AXL7jh
NUhzoJEOMmOD05Yi6szLr5DB7aZ4qb1pbetfK1Y5SFXQSygJcgm2awVy+V9djbPgu+hbtIlUZu6D
81tPDFjsI3AiwMcWbCsvGTZKe4W2Y8zJGXd54NlGyK8fQT8PfxqJ/WYOdVKH1gEuL6dbCXl/CJW+
djZeXSf41PU9I9zsq45R3b40dnqO3RRIZVgb7E/psi3wmp3xAhwh+CizUk63wuCPEuAiPuG8NbgD
VZzy3ZCNQHTDKFq4S1gqjV8NtAH6wm5IgOVv6jv3GJ+drUYdJVYHycCIW0gZ7Q9tZ9jfwKDrlh7f
q1m+Vkf+ARNEwtRj48gV4HGPn8qB5VVmDrWdyJeNvocMAeqI7RqeAty4eb9517u2qovx+pzVLgf9
aDFNTbT9X9uALJEB7O3enz6S4PWkHrTKHcRieDBRweZfjwc4lQ4LEYShL+JUqlwzLCnhYbGXIaWR
VZ3lPW3y/fDT4sYH/wIB594wZQx+RfmGEAefOn+YlH+lbFJt10+E/y9vZVi5oCuYRejgk/JOrjP/
pNls4pC4/vzsjgbRJl45XkKH4BJPzQkdR2ys9bF1g528VjfQkeBkPx6DC8xaAzWoz4zdXlbjX5hG
2q20MOI0uKLCF1klKc4DFx2BrokhrWuGN51OcpIz2IfkIUxA4Hat/DxiXf8aCcqmqELvZCZwxyLl
6e1queBfbYKFxbruEDApfPoMC+1yJRekmOWpm9P6uftP8Bqqxn21In2nEoIxPhfWbbiedT71m/26
GOWHElYzVm1dyIz7uiX7cR8NhJ/CPfRzyB/Oa8lMJl4NSarTGYqKy/eiS5RpkeCz5gzDj+1Pi3X9
nr7SOoM4cBwT6H+NyZ/hWMLqTDUmuySUKaZtrlGmTZoKSfUphmAvDjc7PPwVBL63S4jXvKPZDett
h/RsETDlKgzG80jrbODCX2yu+0KHXAXnnkse+ZT7KFTThkEE5OgVg8tuWNPvhAX8MHYlFWpb3UIx
14ojnd5L0BAzrBVhm6XaHPPbDAhybhn8I6vsw1QOMMxL7Iqn/onSCy7OLm3SVWKSRHgCosenVATF
wd/Wd3J7Gc/yLC8gOD6xDDnEzprOqL0xH23vhOjck46AwxSqITE5jhqxYroTINC/TWtbeOPV2mjX
uPnByDYbeuwaBxx8+wGzt0X1yZFoCAL2bcTVH1yNbK5xTA6+6qebG5M4hkuk3uAMKgIKbxbOa6rE
q4f5Ei6zm2nYQtMi9dgY/Ylt3AQ361DnncVr6zU5MRSA40zIFyXQ2T51kr1+76u7uzQ8wd7Z7KoY
Xeas7MaB+zyuinXu1ZA3AqnXR6YMkddIImkgCF3p2BJH1CGRFxH3Sxz6fgKzcRuYiKZXM/44aDcD
FpHFpLpbaR35ud4B2xBPANg84S+fj4UHSfP2nC66sDWMEmkXzjr+pWPRcs5ZeQs2UvcfN5qxW27f
pVo+3ILLN1KeQo8pvpD+7m8cvJ1GPegob+lqLQ+AbdPZhqnG+vXv3Vl1LJ2DPbqrsZBFf7biF2Gj
c6rmaUxaDGQ511Z1+Sb8jjmydsMl53kQ/8uIQKknEKRgoQGBQgMCee2KJWefnp6t8u5po1TzaFnt
hEEgaKHL9ilkcUq72lTXI1cf9M8/OM/04WDtcSpoeADO9HDd3RAiEzDtu7utkTvrFt74mh6j824D
C1S1KS8FsM4RCCXe+5nxZgssCd3/lgV9steubd12UyvMJjJLtDIPu2ytA4LBCkTM8TuNIMR6lyC3
5GRxObmq6wf5u32pIMFX9jwxP8qpQVCwPKUChpPEKVfcPZeIAOyyV4776KzQRv7sXnqloWV3/64r
Xcuw9+otHMt/ab/VAmqS+jyHfY+DCxzwffQTZtH+amC8PmESUeOjtbbzW/oFgt/8Wun7E2P38e0p
DmkynVVfmPmsG+Oze7y6K4kRzWVlzBvYIZQQPfRJpr4dgJ9v11vdRewSwTmByz08UFfDl6ZZxIHI
Bdwd27IDaraOCgDnwt4z4CEKMqgZr+kS1eDJrPBPfIdNUDFJa18PSUcFzLgVIxTdhr2tjDLsmf9n
hgb5mZUUyAH+Rox1RwMhWO9M7LuN3b74D5pibNYk820tfNaOuWYB3T/Fe/1ej6lWYBAYuzm9O8gj
hQcv6kF4lCW30EDU3HJa0lyH1W5Ksa2n25K6aCc0gMInqgBUTQYh1wZsMqF7tE45DdrM8F90xn/y
p4Gp/MyCjSNJlu/e1n3z7Z+/SazID/B0rE0vynpOs7U0oXa+mCATgJOUWtIhYZ6vamCMMG2q6EWV
eBiJ5UclqHOEjjvf9+ILNvYutxaNWuac58vZWLYPya8W+fruKKLUnLmCpGJaBzsb3PIg/j5lxuH1
2i+Hl8lhv6KpHsiJ7bKa2D4iy2bkUFHpZqYmOH+xhnFSoDUvT69OFmVMjAr5lFekYu+T/FKff2PR
FJaf9L3payDLgNz5RFzOqVcKHl0zsDrsQo2llzD0ZxzsUGCKyQNYSDMxcScSsJ8Ec44UbDK/zNtb
A7GnMA2X81owjh0qzrC0j1L+zyxKgbFEIVZJLjkkqsVJ+9BiXjwGxtVGE4X3rF7u63H5PMwdC3Hg
4BdvFmfWXTQbQggv7etfxLPJXSk1kxOkCx/FhfZLBMfAyE2SM+RpMGaYXQqQFFDT5Yix+7YzT3Kg
u5Z+rVMxKIL0EJvP9HmHVL8zOOv+ki55r9NlKQn5H6Pjh27MoBu3H5kfvhS+CFSwmprUW7BahU1D
G4vOXIscKYbEzH/2wt22Jy02svv/I7HsNslo8vb3mot7745s+2wLfTOZ0+QjPwU5ilZkAC8Y2gmo
4QwAYPgjBDUY/9WgfaHlrkLpTw+V2LowBupefDpvx+RHn8h4B1mX+wKfJXma/zTN69AgolR9Swak
obYOXTSqzgSqFW47IIY6SlWWTLANSpSskLr9Gd3/a6f7eEhal14c+kzGFynUfhbvtByL+uzOKVDF
08QnS3uFrhUbfH3k/l7Py00Mli7KeVz8/j+uG8r4Hx/nX8vpeL6MhmL94Um1WfSvtMxQ+VA/HNZm
FB71VAcnWmCB3O7jUUlad/9hJ+ksLYhpi067+A8nf/WCW2uvzCuhUruh9YareM5v1tMu3VW6j5Mq
1Ax7BcrkpW0HYMlxeUxEgvGVmyvxKlcPlyW6NsiLZqnfXhHPy2nZ2RnZ6o8RG+ERQwLtwZPHsspc
CqxgQxqxT+byxxH+ucib1QHqkh0+IacjMLnV/PJTMH4ApPx7fSPkcL9F+4V3eTubdE+DydENO0B2
Tq4s/r/MmWIajCsV/Fu6hlyMyQjAVBRQzTQI9fKt3W3xAFiq+N/J/zxKzH/NHD6QgutKYiSqDMKc
K4yjZQOcvHT5x9iAVa+3w31C8vHYkb45pnkVz/tF2KFy62DXxEQX6TF1uHdyAKRNG49i8s98r+ph
pvwrBZahyKpGMcI52sheQxtmmq4+MJVmAf/0Nxk5c0wllUbhyGpKWQT2KvlIcRusAK4nitCAqD9i
i3TCjvfm40+x9P/ddfzcNx1sK1g11B+rxZhxBoH6A3fhv6KLbpMj9b1wxyit0kiEzxhqWDuDX+WN
yAPIjtSTxPuQNTHWDSet5QhHes+Db6Ue3mlyDMmuWQxzD9FGqJqYWVpHpuridZQMRQ/r/BpzFsVL
/SMb7h5ARjMNxJxDRn1PQSIvLimCOKF1EttzIKejM19rqkw3r1l3LIimXOOf+WNGcxpXzk9h5jJM
bR+hG5Lt016qkbe7uh4u0+dNwB4qGzTstufvQ808gSx3j2sM7po79Uc/FqtY5NW8/F6eeX7pPuNi
NNxoXzQcswxGXvSjTRTyQ+YzxG+ST3/oq31wy01YGJsTGGHfpiR4e7e1RCkksptsEq/9wk4K8KVx
R+FM0MhD5QKMKHC1WV6y0NS4sHR0J+6jFdbXpCNEVhxnXf8Fhe1qV5EaS0fIne5+5bESWtdIo3tz
pPPgk8+JMSH9TpBBEvQnf/z5ooo/OK6QPx2IhIg2oXeWPexuPYUGdk/1A3Dbk09WxPArvYNP/Riv
Jn4BHCR4ll++5x8UKEdq4eX9xRv2BZyYKr/iYImwM67TxgOqulXxpbOUSuPexUuexBtB9ghEhye1
DU5AUiAfLrPYoovSja357XsBC4T8UqtWtHzwAmoObrAN5eUjDG1CFrfv5qvJLhy1TMPdVYJNFk8+
gD4Imb5lh3QNpGH6yOvNtBKXdd5DJSpjHkngs10i58uodXjgYIZjq5NWkW4qFBRjFB3sFcuCfIj+
5pAKfXDOFQ2R6PYWyFsjrmyqZsTHeHAbwKvZsjSY/dG2Uv+uvxj9bk/IpTs3Eou8TymuvUDbA4pt
bo2BRocRTg3sN+JcpaELAZfHRUNYulREEe+u8IaCIRoDiz3LkcxU8OUU7yziM80qtXfZQAzhpGd9
HRX6EXwp1nmNfLF3bZw3881dhuTO+bgpc+QMTP6lz9PvhHY/P55xmSmEHoRWdKO/NLAnTcHvCyPf
Nv7c1pXntCunk+60fCcFWrx5uW39eOVpyxMb8Jcv+oO6CcX5wd18KJkJqG0n9QGCOx1G3tmtXwH2
KcMi5L04BgX/26jJufNTEKhGNUwnFxI6JRNaDVjF/3CJQhIBjK2pUP7x90cReSrxrHX6hQ3DNAYa
7Htg9JrOnkp4v24zLu6fY9H6Ra7uFF0+G66K14wxP0A6wmRr3Rt+2B7oXaNrXPi1og5hg8ipNFSV
CKFxeiUFBvYoDxNjkSeyqGFjwSpv+gsnvjYcVnYsCwYHfR3OvXSTXxsMGVfBXDsST5dtciHeLL+n
6IB3IXhnSh5+9ISO33FDnGyuzxECM3b/NZOrpQKsC0ZOZz2eWoqtS0Ih1CeXPTW3Jw2P6qlXZbXR
30qrOBuKjos6f6/F9GKQ8H78R8tznTBYoUV3sbjIJZdS/K293rZl9ZuzyEIXT0ncX6FXki4/rciU
5iIGaeAYZQV4OsUEPbri/an4mYNXx4AyVoec7fIhAUhj86vdYIcU1F6fgR+yGg/VLmeQXRvNk2tL
ITFJOJt6vMS5gGZWtYqAfe7quAlJe8Asg4ucLemHjrrFa4fC501iFMJgMue6/HwCtK3Z35i4C3X8
+FpgUwM1/yH1tx1dBDSODrDiotq0IsyrKkuZ4nJipbLrfOyYp+koYcAFQV/9kHB8IZNij9GxxgnU
d0ZmKLXTvdM7dM4CTjdTKmw38lk4QxoavRUhWyJnD/MyLRMngj28nMaO6UphIz63iQo7OakmpTkw
EwH8O4wyrPM722gzBIq8MWw+TjyVmVAtxf+C1Cua0YbM5+rUJp8UcwY253s5UBby65c3gZhaI+Oq
4XLy9rS/eZ6bIL/OCBA60DnaAJunEyuw44+/aIJkEXwBGusGmbMWkXO8vxcm26xXWwErhB6d/KTl
SwzRkqQ8ozK7dZmpi4zTlA1nD93HkDiCd/1qM0BERWFinchtMISyK3kL4EL9qqY6AKbhwRT+TpUP
O4xXreeg3oQ4GK6pT3fLr+zEHg4hNINz2HSn+aQf6spoYHV/epsMpbKobMZsdJUrS0nHruQB7Dy4
XBzro9qjDEQdEmfT8PbDGjneilDl4zm2m67QpPmNrvPZ9xupNY0U2iwDvN4OoeaV7jFnKuVYkjFZ
lPfubr23sZal2iizXsU/YPcCoZ6BAwk53ccyLthJpmwjp2/1A8nWZzKaBf4vUvV1R7hGymGbTHTG
gJ9ypv+0HCfeIE5YmNC/7me0PNVueAsgsShdLJiMhQqDpfdxfB1OrrUcXATPc5VCkHr5fW/En5j/
xkxDTsTHDsZH4LowXsV/D02ZUMc3F8erTRKDDzSZYeJyC8znr5uSEMwbpvM+sYKNLykpSPPVU4XD
j+PKDKJIVtH+iXJJJdhoyi+6nofxC7faMW3bMv4X5J6lYRm5MFbMEz7cQz+86zKyi0LHO/1oiciv
oupyb6HC/OsITbMAz+9E7YOqgjo7SJDs2p0N4gdJ9hllgBtI6hjskSgv7ro6sD0h7J+GQFDl1EqJ
FeCQTxlBcrY5QO7C3w7UYNIjDk+ghExlzxRregPC6f3PSd1wuQqBtsyabkhNN0ls2lNfgzDsYzSW
EjE5tRZYKWWMAQZ6PnDjp1u4k8p9wcbNSquYkBDY2lGlH/WeagKBTOQlXSXvu+wuMO/ZpdIrYI5s
Ow8RJZSHgx/O5PLyeYCfzlfkax5Qh5AtxiHC7GmLC43oVA10VyAu8jWdTBcCxWaqjcm47pDf3yu6
gWTz2sicIPFxL5S4qISAb0iyu44iWrtOV/paCecGltvx0zaly/QgxImdjK7UTU1NNq0A0EMAFc8p
AN6R7cDX57wg958S19BjpwjzMAotZ3NCz6sMHriG/cqaHfnO8ZiPqhmUA/d8Ck4KD5fd/eTmzRjH
nCOLDc7xrmwTDIAcyBb4NpjvdIq5pwzBMu9UvPyjc4nh6Lp2ncuUdpAk0HEs+2cGw0OmGyXxmDJE
+J/Y0atXiwsKAEtwRbDV7OgmSC8QrNZ3QpURs9NszUDZjB9eeEYexgOZHTF8piNIaYVw7yUzSjod
4x4UlCSdRTwOmF5GhnBz/94lgiD6FAhVk2ksj8RbVakOIoDeglk6jPAMzxCckYgj+ZKGKDjG2Qfp
MgXRG6iaDlZxjvgYcr9ys90epbuGaKv4x/yd+z6hh4ByMi+FLYhB+uiTsUcie2LgXRBJk0sPKaOr
FJD5wtAQAxfypPnTrmkbi9se6eLv+4FHzfTWSaGuioirsGSAbyj4MqIZpn636GB8eix+BGK2GHD8
z9K7thO2O7kZDA+r4koBdhIO9jegDe7zycdpWXzJURbpznky19GLdOdyhQPfsqYaVtJ/n4Yrm2kg
CpIBdtKIiP5SlQ1P45yxAWcrPmofvMRsxlxCubHx+jFKaZYQSMHx+8+PvkeYOJWcfyYlRjAVJUgU
XZCIOgtRS+hF2p1pjlDWTbjgdRUY3tYUJjC27iwxwBNDh8fRAS51/bGqYj7/6I5C2DAaYs7mQiLV
W6rDKTVgfAn7yD5USdwUn7N1TSey4bN5W6HXezMCvWyEpTxrSTW6iiFfH1s354PYer+R1S2W9jMX
oT+PJu6gbbythOqShkXlYNvzEfZRPxX3NadyvLfCKyVHB7GNnP/bbP6+8XxCX1SoSLwev5I2rgCi
ZruQ/EsSvNiYMIZq8gAKP5NDcFS+cP7xgxAxf24hf0GzKqIrL7HQkPLbYKFDKSICDn8iiDk3vXKn
01NNafrRu2p5G9Ga+f7R1yAdrt+JSk8Qqo93qFsEGgRIwqwPDMh24vL9v2PZJ7BLIhs5/lsZ53+H
Er9fBNimm7kjkavc2q7s+8FR5N/R3ZlXkiOeEiNd2Tr8yHS/gXFupIbsAEacPsGCRdTaTMzWb7yh
H5dIbNmXU/aiIXCJlehivfCDLi1zzg6plfQqCbglQw7ovTnv+QIGRxEmJN4iiA7g5rzqUKdeahgA
grOE358Eq1T3J7smObTTV8V0VWlyjoQMNIiWbN4R2O08lQJRhmN7vF06wtrGsX8oXXIvWG+YmI34
WGuA295C1oXLwxAW4HJLzVZHcsvItecbzVw+xEioggxBAyUPyRgy5hb4Fk+9GCCim9f7EBmIoHmo
xxmguLLf1bXEeYlqva4skIx0yImegxlJStehwzG8t4VJ294fExC2dnQIQQVky5NYdl1OcDmh2rft
BfFo/sZTAGAlrmMuVeHdpu7CM1EekKfOyMu2jYm0gizKkMHiUv94VCskhXUtqFWRbLotNIhgC7wN
G1cvBrSi9h0ShMhm1BefsPBHTmvOL3L8rh3uwBeksyz8Yfw840J1soUlSM99CPai5Pu9ajO8E+rw
McjmjZYsbI7POpJVvVXFmcGoPLO+2D9PCt0onIHUINIVkKqflEt6qxYt+WgCnlhAJjzV0b+qwN2f
aGVhkEwxzGAw04oLK4YsZDbNwD9nBKZzeryw/RRyKhgwiDUWDoUCToboUWyC+OXfOkNmEQpVW9Va
bu19MkXj/BF90R14q16DyzjJyIpsEdUiypZcwPzh6faU2rbIpRUyiwAQ9wG3nBsk5YVbd879Ot8P
NiUeN5YUhLvQnC+cUQr+VqVY2yDazq8i/IXS4eHU+uxi90iE247lLy324WFOFdc0OYtQoTdfEByf
FriYh99nYcMpz2ciH1nENdtwqFthmMTA2tzTkd2DKVGkIgwMxigDQI4Gv4MjegRYdOaZ4KY4fBoU
Nq2OPUsctc73qMk1sge072ypnw5RfGCDfhBuPiSqAd1Ux/nuvxH4b+n+1DsYFqZ+NSGDWeX9myMN
gy4cemdJ3zoK6usFHn++N9R1dqdjZTmxqxAgVLQrSu2YiV0ya8q6OdKXvOxd0Q+nWqjO5PBStjJp
tTU7sDQPmLit+rTKIBUZwSr2X34aoP0FxdULqCfM3chPYveryx6XFB/cq0s44Zdzd6l9JImVUic9
BiM2QoCvvlWqKzUj5qmCr9YJ7sc46PIyLEO46Osaz7TsrlOCqa8F+nkW5Rv/KaeEg45S76C4foWr
IcxBvTKixREKL57xP5NvhauwRm1z3Uc/KzNGAYAratDLFiMXg1/3tyGU6Ch4XudCouIYvwJ+RK9l
fw4LFYVLUlsjVpvcVVU3JPGGIVSwX8kkM26SduSd++/QSJPe6478i0BEI6+RKGSRGb8GC68gxFwc
S3rVRQVvMRdmUNtM/a5E52rUdIff8GE6Ma7O/LijX/lMnMOx1tYaNZvdEHfPuEnTdVMp+kc2C5r8
Xb2cHAA7/pJugeRWj/0l9PX6lO3660EmG1Z/UpRt5euRVdRA6jxIondIRSzV2ld0+fJuGzegAVRp
xKeSo2R3W4SAdrX+rXQNalCve8d1bAJBqSDAmpeEjwaSAITG9nKDF1W5szROnE4MsUKyXUmHtVji
/jMXC//yqUL2EZl4VLlDoiTKi8cdNQfomTTLbDPkMkKEJtrdkc3Nw5KHfbI0x8vDt2ovsRdXl2ST
AS4/lBCxtXSDoYpcGXwvIFOP3qbGaf909O8XX25HjZt7BjB8yS9rbmtZANQAPB+8YhiSGc9TZlgW
jKYK3hBYOPy1Q3hm8suxVSHoG5ZGu6IhsXVz7wqf6oq7d0LkD/YPjmJwbhHp88f0yPoGCAW0/L/G
dSJqICMkkLpnnxOkTHihLSQbY8UmigsghTefFqYWyVDGfsdtm8k2r6BrMNKZ8DFyuGNovoC8taoj
0hgU1+dKXmppKiWwFF5rsBAyAapmRSGNCNAjDsj3th/zMxxi3zXGpjbIDS8COvIi3LBv+AkRt8+S
Xxhu+aM+9U52IlGLs+Ervz0cRGJ/r8fV9wH+Ht+sIAFOi1XfMT345pc/2rr22MlejRb7c5bTcMLh
U023rhSQ3GLs2ocJ43Oi7IQO3nvl99eVcJR5aMRo+/jo8YQ3wR2HQu/jWOyldeZ6dc+FqDiQuSgg
7nmcs+9zXgjF8y842oBjnXNXHZ8qYYaE2lDUQy1P0j3OeIG6waB30ii211sYixp2tgl4HSPn/CYL
YtcVAP+8EFgQ9zqbyazlmGQ5XcGgkuMorGUD5UKwgaf4MSGRamwQYefDmmmqKUScRdyXhZM0jcgq
siJvXYK68S1InPTZhvoDJck4MJ9vvOKl++fTVH34+tqr0YpgXkHX3ZZdWzNL2rSUCRLbdIgtF5HY
Dd+s1+I+8trlM7AxGVKF48aRLPTRwJ9o/EQvIj26yWho4vLhr5Gm5Cg/BLyUhcOoK8u755ooaLJc
mnrElh7PFbg2HnQ5Ao0r03py6iZRIx6ZBC7cZQq00rxQcDB1j1BzBBgERm8QA+wqTPC5Pd7VQ0f8
dTUubtELa+Ir5UuHu6SSBxNsBgYbByu1nnEbA5cAzpgzPivFJ83RjS2I5SYRoG/VrxKYXrMlADeh
lRDwMxqG7+93yKFIP/EiVwvYfHwf7XV4k2BfKWGKCVPPsb2WxbCtItlB8AXtk9WOJLWSn0Kcffrt
JoFQQ7XsnO9NJim6VPMPz23XlfTWomQbld/Sizb6PEvqGKxy8HNcMG0C3d0fMcs2XmsUjfOB/dkc
7jo+eQITac6lAEZ1cywl2P7iDUuMBMvEK02QQ2Gk5NXoz+pzECqVj2Q61GIpr/oq1ii3KjdYujS0
SC8DnclDkEkdFMYTyUt2KzXOzR+1c2m6ImgXiPE7thStVMjv2jv82Oql1xz5Gj/dROE3GpCJ6hv8
TUL3zClf99CrVPATHwBkxGyLKJ0aAGVJGjjhVlZsZzmGRx+fIZJOoHj328OePHk0x91rJ/cKaOHP
9bbckBSgvcdqYmDfjskihEonvf9csK0zPEyu14gB2PlHUg0jpc1qMxdKPWlXJxT+Qs7D3Ofsny8T
TDhn6o0xsYd2jTfiUgMu1I/4N5EEljBIXTkTiXei2b3GB1JhnojWJ5pz+d5ir3Ww3LjoM0vb18+L
ecf0EM4a3C0FYSG834AHJEJtolvBn3lEFjaoEZskDl5kuP1wphTz0gkz9T2f66Li9NpseYY52cPP
IPGUrMprOPJn0sgt96siz1RTNj5QiXFa7c1BN/DirBsDU+BIzZCqHNaASyK5OHTQB4Nw6xK3j46b
vRChr4FxSCUH9DyT5SAPWYUWLahk9XoHS4Yss2cyU6E3rjqg0r2Uy1WT5x+4PNKqnbuuehRZBL0O
EOrU+XbYKxUAbVQz3GqDUimOKZ+KLCSJcv1HCle7wmYTgZtVxBk1v/SKlY+r0tEbYlyDFIyzEX/n
Nd1GXmDkVwsix1XYbTiR1OwmJHcvJefSRApcoCmRKhmxBXkt/G9yNh5pwqvSmJnr2R0+Fd1KxA8I
3IxOnsPNF8u0oSHwBuQJrQChajqVdKKShz0Q8zvLg0MNf/7O7wvcKgnOvfFjiJXuRn0Vm0y5RCmH
YdpVBQxgJ2zbMuye5PnXMDmHN7kRQRABr3qUiZGsvmhaqoSKrwHwTU8QeByFsuZGz+zZbCNDwe7Z
Km1LeFB/bl12NOD7hpSaAOrrQ2+2+KgL0sgchr8zDYGaMXMIdEOcRGZ34C4qLpey+EXLdmaoNy80
YmXQOHjJQuJy+TjCcbS95DCvQH7Sq7I70sJmpAl0CbTARU8451mk/GGi4x3Xjjf0OPbaGoVks+/x
3BydvIBI3JnG13HE2ewcwWh4W2zkEJLeczJz5iibrugFjSUQHEw4Ec/kQO7ScMNvxIADJ8aHmsh6
bjN4z5I9NM3tDgK6fX3mmdRcmPGu/r6O/ZDef6/Sy1kHwtxXtrXLPZKUPsDjAYmZiYvTDTw1du5J
SZc43SZaGwwNUD212AR2sz5butwHrWMapB/38rNIxOfLlhlNANKmuEku5kO9pnobt3mcYtHBXfLu
HfwxFbh41vMC1JdK6rsEcxerKtzWSQQbUQt1W/aIGfcvBBWz2UYD88m8CRYV0I8UBQZWrG2p0N7V
DfVzrrn6k/wzuMVc2Uc2ojbhDIepOqTcKpkuhx6JBI6eFk+x8KZRgFjBYtXbqnPQclvEP7nhg6uY
/g9KZjOU/MJy+OwZtQRF0y4Yo6UtElba21EMVOh+6fBamM8lwsQmaC3y7IvH2XBuJCJmQ1BkOoYm
M+bcpqpzCgbZZg913eqFAwvu6/h5pAa5NP3Rjehhs7gGABonuG9IrTfr7RadMbD7ZSDvbuL2IbhG
21DOKDc1xXM3KXZH3vZ9X3lAxnKPcaA4uvP3o0f88N0LEhDZTTFa5ZwZ3DXLwwoF8QHY2SRu3Ytg
M2zhrixJkduc0Xpw39I0Tx7Q96Brie2y4iW7qDqnUCvOjnXhBXIjaIkkNchr8nmN8iG7HQIv00EN
Kt/b+HESRpoQoERD0qd0rpkpRo4bp+MmcMbkiZPirErm47loJ11WS+thoSqYWBMLV/f2K7m/8Bif
7Idyb4ycI5F7J77UFvhx6N3+tFtCF86ORY27K5FoIPpYcBjDHMJnA/rHCScmpuGNy8VFfKEYwVjV
JdSGQGrqk8hI5QzQKnDNqCAWG7UO/G720A8T6Wy7lSKLHyg/lxJfFEH3YaTjviyhWjPw4Ktltkem
R1Nv3Jrdv+1dh/uLpuPNS9IY033IjNriijeMVYp0QMeXZidunzuAZBm/3i+Mir5gHyjTOQFt/Gxm
LwbIw+h8OmUuh2ucP4uOhAWnwwjjDbkyWJQbG7Wp7sILYHQl9e/2L2pCbdrXWtLKNCmn6vaXTtoq
y8bcukyqO75hacpYCKkfsG1cyaaUd76CkI4qTO50XQJ3QqK7nRn21vST3hHIrv7RwPbhyEWma9Pr
3Cfx/ek+Yzzy89WG3poQWn4tl3llh/FmhPag+w2zh116PnF2rjOt8ZWas5H1YAb3LcLDXmUcRL0f
l0RFnQzWG6QnOn08T+XtuRvRfRQ93udXqBGs1n766UtPd+j7kK5GeEFucbhwhRYoE4F7mplNPzv5
7jL1dA2Z7zksTkuhVqliJufLAc1KpvJw73SuE26uE475xsC1jvIMmiTtR5Bc8gkclagtkVx3GpfY
nx11CiF6aFRUCo1AfKT4S/2gknPPpjdGuqzjfv4dfGgowiqbEPOKGqxyFlETtPT1TVM8VIY7yG7G
PNHAdKxxq0FrkT690yAKh7vhoh4x0BxYAjivaiwZLG97Z7Y4yQtMo9fGSRulQ2KCG316uT6ssrbZ
eEteMRs45LrYerQqMO8MYt+mTzYXqojndM33N86LlJSZOxFm/F++pI4mI5US6FW3MZWTErnQ90K6
MesvWgGRZIO+jcCT2FDkgw6jUShI/uwGx/JGHNnJoeb4KpdeBHJlG4Gbpq/g516ZI7ZJ9ZWrOzP1
j6Qy+A2NWyH/PfQJ4J+j6ro03FAPSvyS8FwkyLh8YTxo+kDBcbkHxs3D4mcYO+CHPnZ60BNt4tlr
Jiszm5Z0P1ZhlTrmU+r12/GuzWc98b/QaSiJgjaXNtcd0EuPYny6om1sVGdBTTs9bwA06weKnQuR
DhGRfDsjecjESidsWyJn4DPcRxSJJ04OJx7kIbxc56ebtRYKFtap23AljUNMCDZOEsuZZHZQpd/t
Yx2B6kyZpneqpCVBcz9uM6Rdp8j8MiorIOUCSqc1VwLGd0GmHmjcxnQJogypkr6KQxHzQYvLo6gf
F0ZOezZNJ0aYeS0DKIq2O7uL/3hb0zR8yk3EWkVbU+q2jWLr5sytV/Z69A3wy5DxrGFxKj7y/620
ZepXr+nlrhKsoy5mZ4akZwMmv4ucvOweVa0oD7Vjt09Y5OQoikf/0o8Ul7qg1aetSoQrguajx99D
aFCuvD01QqtUse0IqyS684c2eRXDbPBT6wUICzycJw6pEWX6f9Ad9y3t/hiRZviNxDNRZ4u3/sOJ
GKq470lypyRFWXAtKIDWDOzoQlXfXF8aBOGKap9S7MVUvWYf/+DPq0FOJAiNCYlHHOd3ncb05lW+
tYqzby/zT/238XOI5WHEcL/YpvlNsq7mLn1N5Bpp/3aq5FB1VIU7uC+45A07mfvmHyii6l2bwMQ3
lDczDlpaZ1v261OtgSPMTwyJNtVBRXfSeHRnP3hRDT5aGc1Q7uvOHkMpW7sLyaTCPKF+wXVa+321
YanTH/1Ae5aSd4K//GpsXDIniPi5BM3VsXqeoIR8P0F15Eb3YOpzWkpJOK8RRGbTh5AbJGHwPAzs
E40+QR01r3GRaPlRg1MGjAOdMfX2GwXFw/xn3LGtvR5v8pIkxn5cIlDfApytjy9LazfFtMS/ddwL
9q0M2REgbe1OijZzCIFXfdGOcWIeyFn9oQiI/Gg4t3Ph9NvTYh0PitNk/AQT30Pva8BiUuqYXpSd
eXz8hEsUAlv15MUj9MLm1lEbjYxrRWsMn3+81ZOVUBeG9bjKTOb1/z7kKH89aOF6X1c+FBABctjY
YmA2rn37cbrNE0xTnrwmEId2D5U7YIqtlzDuWPQzehb+otLM/R7T1lSn3JJrWAmo1ouBe5lxJ9d6
ClD3v9HGj50++Q2wZpueM7SxkODrYAR88lnwvOo+BfqMwsIMgBNl8ncE72qE4cMT7gXfpKObVgjW
MhshOqCyRk52CoDnODyFt99TaHUgN1Y/EaIqA6lrSRKX4BY8IB9gjUbJ3Y2MVJYENJ8RWHT6Dia1
KBgZkjuwgSwO2AkYq4lYMS6PY5B174viy+BFa9yERIYXLnLytCMar30YR3sfyCoL5mM12g8XB3fY
5fbP4CgsxNX5WmUUH+0qNO+kJlY/mZ4TKKRfI2yXTuZC/UoiRgGwW7UkPRB+AOSLahKdWIGYL2s+
kto97BVYg/KIJ+wjCWUUrqPPYXTxNjY3zMHpdihelCyxVyN0kw2tt2GKpdFviO8ZTHIuVG/NjX2N
RtShhMFNkGCZAA1hWMFxvPlUWq9eIAn0zSWt7LOoRDACgrRPyWebrsFibeQfzw90d7dR1Hs80rgS
KvuG9LJjLqofthTj1aNvYluKBmmANR1oBzCzguNu/YtoPifJ5ywcb29mNFuHj+tZL7cVwQnfBLKl
bHOgznQBjbh9/5zC1wn66zjVjL6svX+kTUq/OIt7DkV59HQXe6OOsIzcUkYQ9G+m1cS5dU8GfmxQ
nleCoCbrCZcjF1X17T2iZA3ZesdOkktIanFKleShF6tItoLwAQ07kDSUuwiECU6JcxyALwK6Fmp3
UOQm95tAxltclTQytyr7/Rt0+DVIeytMcJQbAgwzgVP1tZ929rRd8jZgCLJicP0V56rZaqPOipiH
wz9MCCu3ekEH80uKrZhVzV41fLSux9r2KlK9nw2n+3wtEP/3lo/qACGlvObCh6KdzqHBt2PMRnFA
igrhEO4LNODMEFDqCTHtIvUFllsL5pMdwY6Im7ky37hHGJJzk/GuiY2PokqkwGSIKGZz/1qDHetg
u36kef9nx4uyMFUjAnXvMiRZOsGEoaw1xxvAqluq1SOeCBEDwHb/qI9U8l5i2kAK23vnPWmH3+lB
Ri+CD1yfOcqgcCTIkRzCVRALFLOTbKJcfFKt9Gu93YvHDlzM75NMS5t3q8bHbLZWqyVg9FJ1ORum
6sXza+dI/8Wd28nC5T9/Erj8Dq9qHAFw9X40YDba2PIJXEBDq8xt7bkrEja5d86257e5Z2uO+yN2
G+KGBIUtxVgl5a6q6XK2Mek1E9ev/Zl+9i6AAiF+OrIHIuEzDIgPr75AWV/AXk0xEnNyW7fpuUY2
nqH0mBun7AUXHmlFQoGMchIhIhAEV/bb6DRww//C+dkZRDdCNB4gNlPmOh5Otsiq2MBsU4DWWRC8
5ZQ4ub13LLFEIGCx0I2pF90/GWBXYkD6RUA9wu9jqFgBIn69Oa1KGEe34jEJxnJU4F53ihM7Ds4G
3vFEfnT0eqIt7IPJOV8t6s+I1guMgsRepJRtTRWxxmsLggl8nzMTMKxoWWXV7L1GUJ5WNiklseBI
Y6+HgBjPQ1xXzswIbxdYYOPxDY0SkORiGOmZb82rCGECGfNhD20kZp2Glj5WiM57TIJCkZOdgJmJ
lYfEgnqaDwVQGU4Aj/1GEB4YLoeWzmMu4J/aOGbkJXVqaPKelfM2EHRiR8UlBYxBEH8zTS67vRA5
mZLCDRKbHHnDuJnom8mEoGcaebA52lTCBR5L7tRHzIR86RmHMeMVrGgE82/Xd/NndvN84nkcnYrO
e+eEEe6NVzftHgs2/Q6+gD3nBANhOTlapUgHWcGEbp+SPpljPADYCZ9Eaf6UH0q0EUb22B+zXM8B
49OM1qI/elcyseOmLUebIUwvQxMKFI5wdek0yvj9ibI54s6x9oKWsx6WvRhuYqtdmuil4cSJnIJu
5niRzKlgoFf3KWvr1Zb4H/0RV8HCM3Kalvd8/6HZdikFSx3LRGW7+4OabcmK6wTFPeoJxpw2ohk2
KckuJ1kA3KAHBPWh9rnchSBRimLN/OTZRJ4dUtMBib9arPJq1KKK5uNiN0MnruvsjLqwcuNlrqwq
zDY5+TXvR3fwU8KN0XahuHt7rcfUu6q7Fj78bq0RP7Pl5RZNooEBm+aIBwrktFWwg/7AiuclO0Wq
djmgOUITuKfIQMsolFOZRn3IMNGpEMwCwJnqeo+fqtWdpYfYCW1X+d6IXekByYrCsEjoFZP114lV
XUsdNoHNqkcjTCYPRCjEbtF0XvtzMJzvBxLUbojZH9yhB4VDc/tBqOU+ldv0AmeAkka1peJFj4ek
AERU/3NrXtBOHgv3Sy1yiDZFSRaLHsHqi4DKRuHu09oZWMD4gZCQmMi5/DJxgmfroShymx7JLLmL
xVPFnCB4sieFi8IEodjLKNzVFIgMRdkHd1NzhUOzzQjfe490vULCaLSz5cIp3A5a+tUF7lMb5pOf
ISQ/qqJgVxR6K88qUFvM6C0d4pTRg1RxdeiZQ+vBE6M18wQjFh5DC3QomAKH2W+d4kGls353HB1b
0G4hB6jVV8pR2Ub0JIT8PiBcPaNKlrZhMJkYMGLIB2XgmKs3zpeNhZ3KpKW6D8VE2/dutwrzeH4Q
Zm550zDV0GljAiVCka2oR+izVvOGUt/WTGFLLJYJguLI9kF4xgVehgf9HD26TTUvVkJ2o4zO3Sha
+yosyvYOFzWHrJ+EQsb0m4lV2A0H2JeQhjaZQaCLrwdQ4+AoVLvGN1Dg2JO6VUmE0Q1eYH0cJMgy
QOXJydM5ptoXltvNmYxPQbJRO96os3MZYrvAdI7nDCJ9vS0JMhIu7oF2LF0ZfOsfbpoipgS/voPq
cDNYlK53IQIs2MmSfFA88OpFD89u/5bSc+ROk2KMaXd05875wPeIyCvTIzT1rkvPD/zpxLitxLw1
oUNND5riwJfKRgPYxM2Wx2PCBMDHEpBbtvh5lfWvePXUmqH5y74VqOayIkfM32JVWHA9Ht0cpcsR
JiIRpXaN7zreKK2ILWYLCtrL+s01EhQC5YAKknH2/wWZZP5zpfUjBzRChKlFhr+GH9RtBSlDsfvu
1M5vJy+ftJrd1nFjutwWS9lKNq6olJ3SSZYvoaHWFEmvnoIHLO3nfSMUoYD29zS10l+czrVzqcRc
tqqAs5VGyElhw1zHGJMEugCOwufYl4N/o43NuyoEIP69NAC4MknTPKRVhSwIhDSkRPRh9gTQxHnf
3YwPYw0bNbstdwuGoDm43jcXBcEUMgpPL6PJObqQPpD2kx6TsVVzCOUBfLzKzbJLWzqcLRejsmPR
cpyPyvThinA9YTSpRdqNx9UyxytGQ3p78GgjRMH/T4NoNS8UQCD1jM4Ej+gURm2oHhFZVgUf5Wm/
gyka1iFPGMNWvUPyqQq9g28heqtqIbuuyHNrTcwQNmEQPg8sUZDWgVvkBS1ugr2UAGZ9l4jwnZYz
+F+efvaztrp8jrZ8gdCtvWaMlUIVGGPztcPeYdTaGOqT9JirjwpR2nmqdDwGSV+Rx+kgk4bwpbT1
uiIR1WCh5je5gqKhn2loX81yy+BjyE4LF/+G1PCOjFOZszkszcILM1NidXLGpv6bCEnYzkYJEaE0
6urT7OokM2G/gB/g+Zv9hn3RUtl1joPpD2OfA1LpheD6h3m2b8OPn9/qgeC3AmWVjloREIObLuv0
ENte9OYBTMJopNWjigooTOHjUGgFWkcI77sFBk9yDWJ17ZKdaAouPP5ccXGXoLNwrTOi/Ye1zE9k
QtVA5A45iCvCNCrxtlM0ygigyzK5g4pGtm9LYvTfch3NLfqTWCLHLDJrxowH7eVFRf5AAZv455j2
8a0nveonWKFVsGVpR8bZccyXXCN8W7zFnhIIzwRBdmdkcQBAJ9ccLpr41aAuB16LY5dL+Y/UEr4m
tADsCcvgZZJGYfO2dYsc5LfIo5qgbl2qW8sztS00mMZP1KMmVwFda91Paz8v39vQpN0NzQBAgR6j
Xj402wVQhJi675Xvv7YEPQ2FfJgLrVImJvnGMHp/D/O5wA0tciyykQim06QtF4sZMbj9iFzR7hDM
cSmr27F382CSe4iyzJiub/n+pbKzbjCW+kwVYR3Xy4+NAGKGpoAUBAkLNjlbsch+dqfKDl5l4xZT
stvJfHBGTP1qom93zXU2AW2ZvsUeBkCmMNPFuOo+EpgpzDRLXAehO3QYB0CB3Mkq33zDsDzh9kiX
V4tYjz9uqssuRJGTeYkXgco9+CrTJSuQpygbrsCPla2wgvjVnBUdEp8n2eZrxOXi/ZdJ94ami6i/
/aVo7jq/d0Nm9Q6I6Mr0e+ZKmCOb++N8u2JtD1xKFOxe1D8b/+mzzEOxPThrJLgtjcM6JtY72yAT
wzZnlBwT05jXvS9ca1qJ+2vdw6D+0hxPnQFmYQ3rGRMORo2+aszptb5D4yIpJGtqJ0MDet3fHDNe
Z1cxru+FcV4R5nzK27Zt9b4Yzil4phG9xVnI0RaUWseUV5fhWWbetLBjbMhWxIL7EF0Qn85fyIJw
xxDWv9iYnMA/cEmMq+EniMoXSfPpUM0tFziFa9H5JPTZfQ+E47zcGiIk+zh2vyclpxmU/kqI2weE
NpkojEXV2fOZMQkLWFOW3QdTVsv3yO223wXQKBp/FzSR2R3z65zYavo3Satguh2T25dVUZAVc14H
s7CpQwO17Eyk8FxuvPN32QsnVdgaUWMvKALZcFyuWTjq83GrZkuySQZtl8GI9GPrThDq4zpYqLeL
ZdBIGibtbpBZzQM3BnbJMU77iBPeCdyGXZynu2RaGe6TSYebeauczqCrCAPvM3u6sB2INEJmc4P4
pNwQ6xtk10sLwVW6PY/FVv/8jwg7fSRcgWYyrevdIrJV+MgYGvFWLaf0QkqpKgNBVc2t3sMzotIo
HhlzeW49h4U50F5IAi2ZUpWQr+Z/WdlZEzgRb4uY2S4o2fUig+6uZgMMwE/dq5QDr3/85MIm80/6
56XY0IS9c4fW45XQsKoATFed8aynnBiZxQG+sdj9dS1d0XFppDILHwn3yKWi2elR+MhFdJvaO3Kx
fDcQ55i1WdhrEXw6Ae6E9RJnW95Ihnqu/wDB4F0qKv/cTajcVYTgTLh9IrAdDv9Bq0frKWCooqwx
Li2KIC44+lSfHUh//T3L0Ahc3n+jOtxzzCp7rcWnIp3q+hxkVQoKC9RlbgEUAxql7kihmIAVcgol
AGZNOB29dxTtpUKiFQ2J6j1N2h241xf7Bo/hihmOR2Dn+hadGCeWFq/efcakKycKu1mhhcJ6ZUCD
ayXj2tzMAjxhiMmznJ6nDfGffkCG7xlzIDsAsnIKxhW6YQCctttL8e52QgImjS2k0dO7ONaSE5KA
2FFq+JatRWbiv32Uz+In/bNWqc+CVVy19m66Gcjnon/wuXf9PCHWuaKqVHr9rpECfh+eQtOnnjo7
cTj4WpCPW/bTCchi+GHko88CCpwdl6jipuiyYBQnDbsxr9VSOom0TJFvJdlhtsNUq+54ftVP23qK
MfYnAT2N3ancKxySNctVK+t+w9Zw2upm1QhePIUvGa3VasrmNzkPI7e+3NqiKmLCIYeZv9MTsMxM
DwIXVU0PW0D5f653gWQMdCDWl9xuTQTdxBiQECm2hvEr3tfSIMMJrI3P6fQeUANJUhNoBqATtXW9
6m9Vq92XDKYzTKn3CAZOiP++vRCj0vu0uV/HbUOj1QdC+Uhpz6QvhoDXMdPWzO8e8YNwuNFwFknv
QvhyBp1alR/IQlc2/tXPs+fx7BQPZNuM4oX+Pgu4oCQwaDt6xlxmrjd8q18WmeQJcOkLpMa0tnDb
MfgcegelrogtCydDjtaNuU1zpyKIKQGiZvu2uNTCC+YGLh9+mI0zv9YeC1eXswCEXMj8AjEQiAf+
B1cwUcmEyKKwz2Kg7izPAKtgZnYg28amjvuUPPQCJSAA3Ho1OdR4FtHmpot01PYunw4jm8kJ/k0t
Dz6+qCzslygGzEU9td87r07EhB7i5rylP8F/ln89VJCPqO1FfplLz965k0l9nPbTSj9GLjyFvl8F
W31+nnyWg+KW8EdjvWEjioqmIenGkpqxTe90k6Vg6aYm5emmyWHlejpI8fmFfltRVqm6btaO25zB
2SGY0wCZk7C69fxb2Znip6D+NTGat4V8u+F4yWXE4RwyQkkHLmQ9mBWCZHnhWiMK3XeT8OGIAU1H
sTbVA42/tDvkP7ohvsDuhGQcxpYMS1VAp2ylXn0K7u9VhHL+uXVtM8GQDu+0VFZmEISw7F+NDkIz
4Ujx0f+9E0G85oSLNeCMqWrHXVHUvST5PjFm/k3CRDc17shfZao12wl6MyHH+htkEN67dXQ/PrdJ
dOauiMTD7Wsi5VzbBggerSuNhG+0TPm7xXeEOfz7VjvklNPX+bVEpulAHTN6Kdzml5AyJefFuVMW
Fw+D99wkZlGz0GwlKqWc5p2aZstE6hyJGu3ZQhq0mS+m+4540fl8W6njRK0AOHL8iHH9bmw1oNW/
sntbYLwZPYvaFplJ64Lk9Y4/qOnBBY0yzYhrOLZ3gQUmUm6L3jNhRNmROahuAjG+0Dn61lXWFAY2
//+mLe+NTX12mYuR7eRkGFUGNIb/koLxpOQjsvn6yU1lfK+6HOhNszvAoldWVer1RrOTqTgk+WLz
NseRSlM/DRpBYn8grJrZ8d960u4d4vR+PUWxbr2wdBgikUZkD28tpDa0r1B9bm3VxB839xr+PMLD
9HxrH14HNnqVjXln4J3pkQ1hw6Pfx9NlT3slalCt6nLfRUQl183r/1hnmbYXvdDEILJv0aSkyNkb
lalSeTADwb0wYGCdu8/FUmxFpgIKlY5c3DnH/fVuTaYTsm0p+MkkcvOibkI444BbZSdrJnUA/WWG
tphTKjRvkrjnFSqbXeZBs1rX9GFhYx2p/GnGCjJmqZ/MT8k29Z904T85LV9BZUtZyGX8UqR2AFR/
5d4ni/sB93Hr7aDgUX7Uo2B30zRyl59RS29MUWMooBoULEcTE+UAy46qI1oe6/Pf6Fe9BHw7IYmY
40c702y4KX5UJSsdDckXzNLd05ynysQ+ZCtq81Ynk9VxYPQExZN0AZZXWp121sirP41qBwybMZev
qQABMHjaDRoSux8bgWQTR3Gf0VYW+SZPIW1qwPfXr/+Z+hliSj8V3XZmrn5+zHOEV0GGlQJOSPST
HFLeI6Zr+1k4UaWLO04yK0Ts/6xGCaxHo+DfAE2vxiDLnnSaLkgrzfxhYWemoNaH8iWOkyy+oy5a
y1UBy9Y8a84nbE3KzMyr6HjXyrRWczKPBZzJ9EuZzk6UyOCLiTWy31QthNrhwh6BRmFq7hdnmLiY
jb++W6oJOS3M1540wDR1ZpyF2UlD2zG21AtjXYmAX+eAOF6GYqfWElfOObmSs8JVOtUGACztqTXg
l6GqchcVkZ1B9FZ+S9Uo/7bMjfy8L+6HDdt61rCy3Lkutxs3YoavrAOL/V2nd12J6DmKW+7oJawo
ddiR7et4ZuQI8nIAeemK66mocECTRW1tP1ebDrOO9MpfsqUGP/o39TknY6szGdrZxIywBESpqPFH
Wre69i2EIpYY0SM8RV2NY4u6tyt9ZOG2hhaLcfa/JsLRHpqC8wjPl0Zou8x96yzNVX5/qPPooFH9
B2vayGnaqN5FnFGiTHrh3hyaRj+H7eYigpvOb5aeLAYu/JSRTZ0sLUqj7eUnLvNbSSFHxArOC1M3
bCJZZK4NKlHnNwh6cS0gKfl5DHmBeC3rbPcsgBC3qCUex0wHZifrNWQB8HWI1fmKmDL2APEq+uKe
m2WnhBae3FVYzRPjnWmPT1gRPNsM0KpKT323IKn52ldiMPsT6g+ktwBLXWQQAlGuNrAEuksU0CcH
tZcpP0nZeaPWl4ldLG7NZhI/EdVCQJI3JDM+/16z1pnZMDt8+XRdyzJwLaHq0g/LitKrmEeqTq7B
fQvvy2Wf0FQxH+I87ANlGMbteVL3R4l/Zj1M3nbe/xW/7mxbUtES2Cd/5JtUl6PhONO41lOXD9vn
k+3R7xaEqVFyC1QX/2S/JL/VIJKF9uSIn3LAPXamteP8X6xZ/96cMZUfHYOmXrvJgH5ex7JNyqDR
PHR6t4dYKoGxCvga7UnwwBb41v/55ockxjnD4TXKUr+wx6fVzFSRVPJNB1H9maKGoPGT1LNKMxRh
dHOznr0xlUBfLR7imn1TK1/vuepIK0yBPUWwFexy6+sFE4bAXUryhXDYGykM8cIVJ82v7qiP+snN
VX30B9RWz4Thk/7QXpMLiuUnXc0yqGl+Fpq4t3Ca9tFV9pGBGT1KS+XJTqSMrCj4Xs0C0tbYLrf9
Hl17QFQ/Kjv22x8wq7ymr5t3ggMlESNRtLR6sn4xNw2lNvLM1YrojpAAl245ptxCBukkPL6YBvP2
qQtxqFyYV1M440ilsErF+fymM+G2kKgVGz9fEwCPhBju3iO60LDjxuNq4Jer3OgotJ4MUdIMulth
UT8RSkJbaV1ZdEFTz0fOFfGXbw3kHM0H+krpr1/kkGzIz5+FaxYpBXH5wFGg1Xrd9w+6Y6+qRwlf
fK2yv3BpQL3HAI6UBwjVy/MfnU5CWccTm06p59z5axgt1DH29nwKs01KP7FoPbNIWUr/v3Ce/j34
zvWNLXjurcX/B9PeqNc0WLR/0OLzcyEqipj4V6leWq1wjN/8GK2DOKOdUOUrrlgHZu7ZKh6iWJRK
kFKXRzBN13aWCr1MpLwyNEllQUxiKPY63VLfHciuZ0pLgabbcNy/W1yeUa5JffE4JERH0oiVgl7D
K67d8coHCE7zreBMOGmNS+5kEiqqjWcKkGikqavB4Ou/5YmoDDowOAf5LYmtlmdhYc/VC5p2f4F/
1pgGTkRV0yfOtb+jrGviWzRtW9viXHWE9meTPZci9wfbhYBGcbdDWjaLMo/7BgCSju6f1N67fUBs
TGE7X+CiI3Di9r4x4SPZLVLXXafuQ/1AxLIz0NyR2Y/hDSRyCZnqMU0BgcRGow/h84so+PZ2xC30
Am5ZxyvucRtOfMyv+7D2CZPoGR/tdtgMljSs/vAlpZTuq+idU/xBpBvMGLV/2sZ8Iz6dDfF4HOHa
9y+siyhyZlQtBGPjUcVeuK152DleEHVLAD74tAJmELRbSQyDMsyfYjbM1N6ip2RPF/ssY8e5WnnU
30d84YOE8vvGeXgn6HPN/g1fJQQeBFUhsUQuVKM1puOqGU9I1Bf0E54VcrM/4Qq2N3BwwKDoAu2W
Gm05E2hxpeeIVhaPh1FjTmH709VIKL4RQV3yprXKFKQUdDNL2mmTdQvHKQZG/kUedYa66S8fZ4HB
z+H4u2gpT8RCKwpSCDdsbrWyFYxu+9oFZY4feOXBNW+/N9/0xiq97Zm4SiyQbda1RlZUCVybK/Wd
ZiuvubaZlwARh7WzfSq1vcXxP/f0R4tALkui4aVJpQ9SBuIWDJYPMUG/mTEUYo8noc2miNJR/knF
sg9dscj3gEdg9QFWhqvKQPDgcJ4kFz2DolhZwwo9tYQKg7S/c5u3H72hOfDw7SXPzxRCQo+seOa5
YEg7yNVZN1sX4PSEe1ITxoqiP1JehQPTrWsqS0OX1IktR+ktUhwhAIzGA98yuo0NxtiuR/YPwqMt
Xs4YrxdlklN1XtyxUJ4CaYpohHr2rEf1FsWhcDD8vmcUQneNZJPJNFisrtpoZ2Vmya/JuJYu3kwU
To7L71nHoEIVCVkY0qirbdoOu/nCiidE730lbZI4cUPeIvupAKIv/hStKFdEnjV+a4xMubcIPqGV
xqZLwL0oWE7AZWy+zNDhbWdoUa7biOgCpuf5Jht8fWumJHZSLdHk9q8pzDa6sESh+xUgE/7N+jDW
IaE5xNt8ftUzx56nIJSf5xS7RqzOKCDL2VbBTwGMYSUBTO9anOW9Lh3FGAm4c+hB0lzh/nxUNM54
T28VGDFNklhHKy2MicIDJ4W4LzR/nL6Ea2B7nvATQxuHV1yFb0KOcS1CocwgOf5QdbGyRnMw+4Z9
UaRLvEoLhyrgy1E5aCi8f4EluRCCSTPjPozJrjrABYUWV6saOsu4Eoqs9w4o8CvTdnZGeBBVnEmj
4BtwHkWsMDY8z8EFMaFEzccIZ3MXF8jYk+p0I7neQYOjnxF2P7AWgfHTWjGlPDedMKVhJLDEAv4m
W3vZm2lkUU0OnCnwEvFZVz0L6XL5W89UTuiFgXANXowXO4cWnHUCV0B6Ijz2bwh1OnPWDtnMAhnJ
m9O4v1b4HtOyG9hoq78/qCDS3lb52iti7OyR7qlWTob1pj8Gt10QMPGcnDUzRnmn81qqma3QnecA
deXz9yyOylrwYtKa93cmyMuQKTVK7Nvup+CHFPapSepb2EbvwJmdk5tx4E4XYTAuTpwETk6egew/
FgTgc+kAeE3KWsvMqoYXx9yW6i8j+Xz9+Cl0rUHLa1Yy+QTUffG4tsc5dwDASSb4tVo9gpmXFH//
gv/2xnWbwtsLUN7nGmF5z81JHprDXaOujabJTqXPXwzo7wbJL5VeuBu7yoEwraTq113zRxd4y+Az
lPThImbLq3cAj9rU7zGQDAkED1scXS7lPX12vjkQd34vCTbSnmxzBXAU69IoOWUz0iKtYgMBcBCv
h2PYholGch31uzqlbFR+pqLAo4HFTqt0cbvsa7CrJjLyOwIN1rlQxcXjfBKuWPYUipSv39owwtpW
WLrUEeRtOHiBnuJvZGFFX5KxlLbmftj17/1+F9ewZvzcoBRKsOGJfpO26EZv4pcEdFSmdvJfLwBX
z0plNbLkg0EYWArb1gFabsc4AM5va6ax/9sKWgH7roiX/IHi1KO+RWpZvQNx8gViqVVgk5LDnwW4
3MUUIrwETqY3ehbEpqwNCdz4sPaFU90LxnoqIsnpM6idhoSHCxEYqsYn3YKIwlMc/8h4ez9CSBGc
34JjfAXUV7AD32P67WOV/noKpk7b0QO9STl3AGDku8xgZJuEOoYCAO6b/Gaze6g60GgriNyweEa+
BpT1E/8LhnUVTkFJmqEQeHhzDpvm5O6pC3GA6Mi9hkVu5bNcqf8rJE8qCcftHvCkaOLFwibPLtSo
66dFB3g1u+PB5I2f4XRFxONexqTrI8mkubMr+TGyfbj0/caLeWBjYrFu4zYARjpqpW49tVCGXfxn
bs7x+v5vEQewsb3TcsVuggvuMPW15TaLtok08RH0QiBAUckJvOfpGhClRzeohdOSh5Fbd+D2VNgr
Q59Nm2RsyQJoD+kLnCpGX9X+5/zNfLX49xk3ukJ2xtworjqANhUgl4fzg6Xm7Rkc5Qm2Oouc8MYc
bU+zkj4uW9ozmsHfKfA/HKhDISOAKKO9KxZDNep+c2rd7KnYqX5QRfzzIkdY5Y9GDU/0P3z40v6X
HJVOkX1Oi9MhV4B5vs0Tm99AVjDwGICpUQTTx3erIww1EBzNU+XigPcrMdLICwsbKhpzGS7ceQkY
ql8dxxKE3E8YhBrKo4HfApFHfP2947gWAlRhygtGvVKKBigfrwJGT0PYk4pLjOOti2nii6RaDdO1
ujdv1/mZ1buo3UG3SAbrZSWADPsgrWMNWFH8RSrBErg3w17WOIew61AAQYhkFFgnMHovSCbHQHKw
PurNUdTly65gkadb7xtHgkRa0iY8YtdGxDd5S8hfGtMLnxcMnlnPk9+9EVAHZWzvFFv6NI3HeO8v
Pg4VbKlV2vsmgJfM/+g1o7nysawhIOHZGUZH2aViv3dYA5wieCFkhZ3wuIssB0Jhxz+4GmhrN9tw
Lcub0dfC5ZAOIXRJoLhe//yV40Gz7Oj7dxTlDWXh7r2LbAXJuxRS83HuyPdsNHBvyiolQVsOkpA4
503APxJfct3OTVw6dLhhk+8+Kk+QBkWO59SBYYS1WFT8jl8r0z5jsMWaOfE2jCOwDYmQ18IuC6ML
AFKVl4RlU4wCf1YMp2TM6HoFT4xN3MiAWw5eqYBxmHRmx89YGg8qOgB9lzCCkbQdm/FZGSM1Tglf
RmRhNuejnitUPexI1gvBOHUBdEIFL+RzFxR9K6pgrVFyhRiYy1Khd+J91jOM4ueDmB1faaZ6cmFT
GseK5oabv7ESPY9/4MJ8HnvGklae+2tCgu2pt5WLCbqNykx7a90TxUijb6hVFXlFLT8eAxhpjeFb
EB29h8vwqAgcM0Xn76TIK8ytK4jZsJqt+RvakQNq8eslmiguSEwmgPLM2didjgHGX74h1xXIV3b1
7vwilQHf4z/EI0/ZoEs7Jdn4T+02SxL9TIwdowbBKcFzy510y2meucVtkTSiXrk6SmPsF21DqURQ
JkllwR03O2Cj/8k+88siiuV4G2VpetFAHCeh0TBXMdrxiM/bMVs7bjKe/1mJGXeINUn1XJbmInhv
0NVr/4hpkwHKpJ+9vrcEVhjmwuSUJtGDfSHxoFlzI8In/OliiYi5tMKWpHezWZSfCFu+lI/7SmJM
qsWKTMhFKw25AoFDHZ86kQIY34gdWuXQoaBsE4XfTaNW1rO/45eo7HQ3QeVB7cGpUoF7cFbASvzw
ZbPrZ9tOZWrmpoDPteiKGVjcqc9o858fv27HMRhldT2sXOoM3HMTfCMom5xAz5Tlc5VJ1QEvq0pd
SGsd7Z8e+0ZCmmYI4/iNYd8QA5FMUGYRw98aMz6jIBK2WFw88+2QrXZzDbJ3gaOXaZYzkjW7LJDu
BXIS7Gy8SI+lfItqNj71vkxzNQGYYVe8/idXRG8kBt5RqhmntVtxKvEJqNp+M3Sw6bvUhA+gwEVq
9K0MCTUwCfl2C3FELUF/BOyFaGzYuA9hWfcEqD+7YIWGuJULCpoVJFbd44A5kXaamGg9PDTHQN+f
yZS1FG6gNbtUCNjPsTEOZpa4n6gQiB3loF1Qc4GqisYlvMOgM9LRj+8YGlffAPMwk9ROk6AewRCk
o/as82Q0dOWi6qZD+/A0RbClU41eSxMRiCtCQQEBkKEcMuwok4UP6+IdB/IsFl+5C0EpJ8HB0vgp
Sp8iTgMa5JFyfKtIuCIUPi7nHzRsgsYYClU1JUDlU6tJqNDk/9MlODIZ+lwJK128AmoHItx+51lG
wvfoL6+th5cBottHHox3DJuojifqZFxx7rdJmnKts+DvoIMhLsBqSzwFlQMc6HEdXgLm5aKsiruz
IPrhWRWwhusAGuE/UKpnqqEs8ZUVmIvepcbS6VtiJIoEWo1NvDDH6YeTmC8UWyT/dNYgxxslCgJw
Kw6f1cbe8WDMYGQMPYPaxr4iUhu3s1kiUr05FrZrmDBq8T3IpFDvghmNOnJrFAZv4BGlg33MTsgB
6h43+hM6b1wPC/Lk9wQ/m4hogspqN3ivPZOL8HzxI72br8SDYB8FinsKNFxAlbdq65TjoWiuhL1s
pAEeu5qCQVgjMnvLOFkfWiMe0SjvaQgHo7o9l5GEZe0VzmhU/ufVNXW8ALLzyDSWEBM/ARyW741P
25BAffjRLvq2zIr8Tzkxy1bHstW+Dzy/nBcbr4XWAoYNY2ZfJYYLi2mt0asEY+hbb4N9SEYXm7cX
D/F3a/drh8xHAM57r7wDT9bMt1UCuDHKPE/RxYEli4mBHAbBZGVup8rm/LfkQZLml/HEN+1LG552
GmU9P97TEvQjaPSctva0+7GrCbulZ7OxeXSKRVwkG+nHbxKXi0QS6bztLRjB44ypwW45R5ReUDFS
kGN6VjBPDNdPs3g2Nsf+ey7Lo/q7ls178KliADmrzrhJufyH/hgYmr6Ruf1XyGTQOUCkg5h/YCBz
Sc/pb1taDXyWOhdQvbORWmO3vTcvvesyjuW7SfhmR2Rztk7VXEGqTlD1pZ4x34KrFgi6G+Qtan4N
q3VQXdz7dbXLHjGiMxtE2OVnOXX/XKgyAzZyAloIyQ/PJe90iXiqm7C3vTRAZP3QofdPNap4rox7
zTz+LTjPVVuKeuNpMmQpUeiNAo0AMw4jFLgUjMBY9bbOLED0hmc9z4EHRMR5x4lFg1NeHXBRJLti
Mf1CiFuXKqCtXUpW0JYTPU2bk2CP7vx4Fs8nure3UnGs1oT/JHiaVQT+lK2GVqHVjDop+8bvLFQc
8iKYUo4zqsqaYcC86YmwVzt5gVFHadscr6ifi31dyCNYULWn7lKAZDuMa/b3SqUBR4PSC0l0H0ta
mgF90KrFS2F9kQehUbZ87mACKQYZYa/AY1nHpkeZ6FI4CW/C60F66lIZ9UU/ZyxSjz6hf6n8I4o7
ydmWn0IEid3YreSt3We+SXhIBo1iBWRfd3kuCrve4WOw2FY4GBUTblGV57dznjyD1t57EGUkvWtB
HkkXNm4nGMxkCBpZmbnGfrqx4sadppEWXNl6z6+wml05j7MiRqssYR+thBoML7L7TrpgHoH5+cTE
X3I3HCikgG117PJ7hwkwyvQKRxRMEavuKwzoErsUWRqW0lhGDrgeEBLpIJ/O6reFksNIOHbManpZ
67PwGLlxO4arGUUc80/KjAF/fcWPz4b3+XNPJBN3B26QxKVh2+sRkORDnyrzw6co3U/blLzVdo1c
iaDhmWntVBmlC0/FC5F/VlfH4lp6ylbwRp/pvYFQqc36M/uCngqhlGVlGETSwDLvohL22vUn+X4e
hFn+ODq8UtPd6T+H3IjE3x5Uj0iVe4NDrB+iVeAIQ4e3KUbWKcySeKZStPG87rBlSzeSAKvK7UFd
zgS56islj4bqeA/wpi9vjLbyhg1tOlIre1/YbiSouZ2TAqZcOlzLNUxOmwK5cgvlL2I1qVV1H3LK
5/KJzrfyJgOHqYRihDFWvB46gS44sXgvv1OCzZByB6pI2wVVq7mSqre+bs9xmexp1Iq5a/XyJjxE
IW3LCASbJ3llGUFgOShWk7GBcLQ/FlNlIa+AOoWM0xkrm1SzVmRRVU380pB36hyJLbG2J6s4IpGF
kQzbKzublio9XhTWfLk9PdGn31OOAgrsMyFChXOPJlNQ5HCfIDZSGealuhjCZFJSkYEfIRG1sobV
JqH3YldtiL08/ATJV5TZodqhDuBBItLb2TtR319sYjdIWfIXrvFhjqFJh2hVWhXdLHsbxyasLDwt
VDZcwtplYppbI8Qsbg4nuQ0Z+uaAguaFbQixpk8d4jgr2c1sIMdy1fBgU6A3Aok1rvnPET40f9mY
LfcN/x5ubZdG5qmBVduSqM80kOqvTdSIUIW6jSY+Gfbq9xUdOO6ztx1SQna91Hhv9dFDWwRjhD90
fBIbkj5JTTT9Sgl1Ua7w4kKYwx3yIvdRtTfmrDXcd2KrJy58J/iKMDquOkwupD0AidkrnAZSr9ls
E6oVOIHqa1jLI9HM9scXs1uiTSUi6U0f/4zdGC3ZuluIQenXeJUWHs+DDE1/UVzRryMDPkLeq+Rr
bscSazvlUidzVpGfIVO0dx93LumfHw7msAAUZbkwi58rtamVg6sy7kyqB2AInl1rvmeQlOf4B0El
lM0NsvNlGpGzFuINdM3mtHZ4ISVf9mPIg1vzp9QvUbg/zwMqcyI4Xx5ofawO2T/8b7ibMYEX2sre
75rDNmDRAVug3/tpCwkDN4dUx3+eeW2t2bTPETOc0SnLfLeeoM/3/tDoBnQiXMHEN4IwFpyPaX8C
7wHBPjko5Di5Ie9nk/PEnfQwwcC/YB1FtzvT9W1cGxXRmNf2J38fuxpsiID6F1mmBRQssHw/ns0V
9ZB61XNUxPCm5FUw2zY2LEL4ZXWyxyqq9GZ5uMIPawfUKfqZWi8tt3h/rMI/JSy0OH8CAXRz05Su
o6DEPxF4HPASXauCQETuSzzpEO5R9JlWLx1p9wXUUtIx4f06+NuqEqEvYfx8pHcwpN9c92qp86fU
ztuC/hBXVIBs8XGyilxI1M+IA/3wwSB3Vy1PWEwObLDDJwe1UdAz2+g/J9jxfPocmQK9dSlfK/Oi
rY6+LPUMaSxR6eJytR6y9eyn1DX5rxQo5orQ0mUhABJt/n+hp8Ms7F/P3n9XK7l35JAjhrwYgest
PtViSmzl8RHWtlZx6lnph1+eLSZ9cFymAdDW+myPo/QZSYOheeCYb4rFfQYoC1bqsols7Plu1jeG
vcv0gClfxKXZugK06JMY43P4WLKvbLEW8Oj8fG0ekV7U5ESwR7FMa0ylrFDb8N9NEEh8jlpVmaPn
uXnEUCWWCt4+2sZPv34PubKmWYFhaa6IWmhLeanCD/DcSzNzTrmOpn3t09XOdzg50zLgD88Sgm9O
CuH49gGSs+zg//6/v0VNvJyLqWp3yiablfA2EhctgX3iLxgvK/9tMKaXxPdvijaXkxviuV0E58Wy
rVk9iLl2qyKog/RHkH86q20tpploeHG9M5u2og8QFXJKwUHje11tV7jai4F44x6/RhsjbtwlSwy0
uZzSzMUMMmUaeMI1pLpQLARSLv2qyGHdUOcckKWbergTEAXAj7KT5Rd/62YDjWTvfdSPY9AxpKF1
z+WiWlRkOr8w/Cn+u70opEdYC3o0yw6s4fguvFLeUldWDX59c9dnApYo5Y4EXo7UbbSNKzzpwp0I
qIDr0D8WQoqkcfRdM5vTvebOT54v83HaDavQC4sAwfGqnOXIvZRNlMhmr6BzSYHWFXX5H+ig85A7
QuR4fvqowv+kWJISBvT5v2MXhc656TGtukVqIryKnzJTV9908HL6vSVXMs7kb1Ixug7KtY9XCP3b
KQHwBs6rFkIvXRRAzScQFBgWqpkJB9UwLFPXj8NSHwQceJLAAkE0GUGpOUat3Xrp5EUBA0+rPhF1
p4d85DoajloeVFQ7uhnklcmTyx1pc4+QBIIi98Y9D9s9wn6bd+JyJllXbfYzhlQ4i9vwp036MKgZ
ZXnzV02P2HS0vAPJfOdlf2hlX2+CI1QY8WsAzlevFCGiWnQNnvK6lT5+iv0MLGYcVsiWQtNrRT4z
cyhQ605R1WSQwCeoYf2wGUjDcc4WrS1olHAHe5vK0fdFelgZKLxylmKLQ/jUzFYF71NuzqtPZN8j
Ygx7UVSTrROvV+f26t1N2LURIf1NlsLOTYK6FptFwA0hVw4oQrqVdYpFWnXxqVhgg5nTqqz/6yst
Zf6TOMiWjNaMlBXNsXL/KVILBThxV+k+japyDN+uGayWtSIWgLzraEJ7xMFE/TEDotdSKGzr/abU
CvWM6M3bxe0jpu7n2bthSVxRCEqDqg6jPyRlzOBGqZxJfpxhzqWN1F5PZzF8wocJLL6FznMNRaiR
fK6CKLdeDSJDJMwQ22sG4FMr8bTxlGPrYbyyoJninazF2o1EtBhvT0sXR/Yvk/f5MvUVVIpji5vq
Z2c9Fr7cvCdJIOGwPaHDxHwH+7WKJ5jS9HfBaWtQL8bfkPzFjb1J1vEpltSQBSlAU36RS4LvhycJ
0CCKFX4yALwJycrZmfeUl/qNJ7AmG2CPZATapk5/MoG8u3MFh6K5WZC8m+x1iM2b5lRdmNaEXJhx
a5nQ0I5ZaLixERCh7o4awvbRifwcnOGzEKBPcVN3puPpnCmt2kH8ISel0zAUy+kLzKqlpfICmceI
2tgIfAsHdhSYCrQydJCJMz1YJ50IU4M9HstU+JcanXjnSdKOu1CHIp+5t6rAVndMl6MNo2qpdqaG
v1Hs8PUmWm9fzk5rvXrBGv8O6jtWwdiMPdNF89sGe68QOyRbdz3Tf/2/TtHff3wfBC/TRsLMg+i0
gUiaMNeQrOhtRx02rE3hZL6CYRp2dqRVL7tgmlapgWfkPLvZGGdxM4aEuAWZ7kWJbLtuthuNGI2+
ApU3m0y2jj9YJzpqRZd9CxrLNLvJlx5Q/hcgQ4XBK2TvuZKfcj81EzbipZekEY/OTqyx8fjS/QYT
uBqoIf2ZQOBlsAn5rOn9lESwLaZaCco3aQ96PyWynnFhECbtnOZ2SHZg8Dmty1m+u1XkX/wfdpXx
Jyk+10Q2GNxQtItLph+Z3eg7T7MoIZfOzf9Vro/qaReZNv4RvAqNCXRGeTZ3kV+AnPi0yx02csY9
TDzapusAjL783H1ZgkWhFl0XUMqLwlDoqol/MMya/1rMzu5i8lFCUVmCJtEvgLRoERV+kIS7xiAU
xyf8vFNVhRItbJ6SwErgqi9wUWRLFyECI2GbhtQZXJJhI6miiRCExfWF+D1cui0EBarYFjpvYpFm
XJ231nqERXIpHiBZeWU+TlrlQ2z1oqtTy1ugiHhbTfI8CFjEr/eXOCT9n+yUvH2UbULHeoIwpTba
l04wrJUL2cmkmwPkD22/pmUmUWGJcXv0FAT42Mz7+f84msSIoQlF70e1ubz7tG8OKtL0rae77+pU
YsfwFRsKbMLiCt4uzILZWbe03itpHv+lgQqREThGK69bHqeFPhJR5Ka/YeqCTb2Lec2DKhjN0Jn2
No/WHcqShF93nrgt1sR7yabSEtqjc9dH4GFJXM6fgT2Dqnlr5zRalAxzgNDIPhrCt+rE3S6OYKoV
0KKi/tjAk3lqYhDU2xvbNCU4om06ssuQHjgtYO2UOEnF+mBzc1GCNu646jS423k76mJzpteM6qvA
0fwZ03MSC8p9nGtvJLASVdJOxD4QOov03Dkp+g8Mk3LkrKCNW+OlmyznwXdPyyvIai2mgTLIrefX
HrBZaKk8fw3vn7rVZ+QW0h4yAOWli3QeKZUEEzqMhKPetNabIM0Lvd8wmI7wzV3qCqWSwYOpOLtf
WyuhKXa1n+GXJECLtPkIB3fFzAvjS2qQ1PJGOngPI4RsGhsMOyxlk64ck78cLsUuJ6pW9nozun8C
a+lxkdDHUDcUR+Q+jUNuU4Ky8J8XFPeYIQSJcYiu7dlTQebPRxixtda0BbKJz8NL4x6fvsryr6//
th6Jt7FANvmNQbdIwS6hzoOyZtSClp4d2mZFfgnQOja1qvmoVNjv6ZlzYVlKv86F2oWGVagW1RgI
lf7i9nXJlkPkkQKS7EmhqI+d/roOHRTCjbB4b4y4rZUdi9JSi+2FwEfmKlZJJD4GliENhvVkWMkx
xIIZKrACutcTZ6REFMjuwEQWlQOlbKRPMZE1A9d9OWKHI8jS7e66oTbX6Y8nkVze5tJ/5Lh8ZDx9
qhNt6HjQbP+fa4rYtGhWqp5/bVVTBKFmrTsb/xFZNLrOPMBs24gu6vd7bwGw7llsi/2LrJ5IqTOz
BW8anEd/je+rdflPgWx5lx4QaftOzM0OCPoXlqLygEBT1cpzmUySXt+4ykT2eD+ImT1tJe2idj/6
zlsI7MWQNG9DVzfT2FvTR/J8Ha8B3dulGg3Cq5p2S2R5J4bWLx1IIUDMdvH11Sv6TnVf0I0KKRQs
XOZKH1cuNZRuEmNeU7LKMbo7LIy4ckCyXlwNfZaV5txKkbLfLGhsI2uDwLObRfoFV0IPEKWkUOEa
ME11ZfpXEjxTZfR8tvx0OeuKB/hA09/+BAcB19bvTlbaOqvi+UCDZ2Co6ji7pRt+pjhFycHvdzaT
dcJY3t+waxWAV/2rcTgGFwIcJx7x1efTgBgcWScQMxTBBINQDFU/yTuyy/MoFeu9bOihNJz+Luyg
j/axe5CnYMjjohpxRruhN0tEA7RB/NNsjhJt/wVTq9xTjM9mnl+5TNuxo/262+INFDnC7hBWjXsA
XVC59z4yo88TIZbdkuXkqteKr/F3tS9d79r6PlapEPaDYlRHG3taapGC8zVH9Uvv19xEOogWsjG5
w7ybaTGHLmOeFwAWBieVfx7nfkqMYPo9sJ0ZusLtqFCSYIx5emeUuIVxxn174ifldIJVOOvoX1OZ
0wPr29S8o5hii0F11+MHdV1T9PYM0Do8OIFUmZfEpZa9EdIII/sbw7YAPxmSra6BLbp/21L4rYl+
L8k4TE5xonNKEOx+X8k9QsrlHSqzxWAjAkVDZjKcW0StyFAMoeCFAm3RHXWJJXnDqKzctr0tcJjs
+oLu59CsaTEQHAc9TdiMhWRZP2pEAW8XIgl+DSevUUJAzGT63sTEXw3JJFtfPBA4KliP6XFapMWv
7tfICa3rIW5ziSOE9TbfQihd9yDGXMPsmNaIKgFeIpJeTgyY6B8uRUdI8lfXD3vyWFUd++FUpcYc
a+t+82ylmkq+S6WcOSAGSdBKcaMPlFXoLQuljS5UZj7i2QiqP93QP8cTVmt1DlxTvEhIX6wrr/it
H/fsLtfuPZjXEwvT0xSDfnV+LVe57IUZnWTxKRJl37sOEQIsFcB3ovaEk4Xx2wN7A2shZYqOC3jN
zEZjZ+nneMBB2BUdC06HNo9HHFanwjRxx5jqW0VW2bnCDHTv8kJfa26dykXDwuQHMhkWkyVxfkXv
rHti/5Dwe5P/EpyVknd9M0Km9kCTiOgqTN9e0Wj4UQhodjpA1G9A4HH87075yyri/4dubAIjAx9S
0xsz+PZr+vNusyid8zHRGQSL3Bq4PmIMsJY3y7dscEytfoLuPNnZ9GlAz5IS8v5dd+CY6uKkeOPT
0EXsm8nAVA8q9JzEzIPR3eYu3afJmgNKi3qBmj6IMTO3CjugbHBzbmpUuWkuX3wUmfjOVadWcmI4
uNprN1VTM1RPGsFDto77juDbs07vrYZiPbjwINqPctxhnZztyK0elYS8Qv3xbkQiBajWRwa/dQsp
to17Z3/mRfvPqpoRLsNgTkJvRgkScm7zz0Aqqcayfftiw+Nouta4iljqeDlYurF8OJtylAd86bKg
Mr5QkpG0ZlcvE7h0YMRGoN+M/wBOJSVBLZvnVLPdB1DMI1xwePgpVdCvruqzVJLqylDU11xK2TRc
GyzyrDiz18W9WcxShEyLLLGlxYNCOXyG9hKHJgKbC7VTLOwT3DXUNgLQ9jCVz4nHNfOe8jkQpbCT
1Ok38dwZNSpnDnj7N2CCBwrdzXPMNGMJj9xJEgxi8cn8gUGrqngMn2DoXBXRIm6vIkFHIKdoRjDu
qHskA/6XGHW13S5I17Uzv9O73AzvYnLXbf++ILEge3+TBykvHqYwjtpxxxtkHBlDhWJTLOKDV/un
/VCO7gxshbfAUFpS22Xmh4s6V4RDciHzkBi+bbK2LJqyKn9MRSGvVroff/jw44uzB5YZ3O0AfXty
JO7saG+0x2uI9S+7g3A+hm6JGTesoBrZ0nYeXkqMxM8W66TKFdE6jvX/Uz0ce7NKtRXZ81dQCzjb
QMlAxbT/HbENqJzy+UaqAfN0vvkhbYd+JFbrqsHNrUowDeb1ZMRDddOyNtRwKaSy/9V53XTfKkuV
AVTPdnfYYl/AvEc4NkwQVI2vVyVEuUwy7hIxdr4zpr+iBevpimNEyaEkP82Mk44L9nLdNVSbQzMF
ASv74ovxqOAW6EHHdhXRZucXgevEwTqqljhhqpjzizFPsjwShAu/5L4ZKHuM8bgGGlK9C8Co+mHA
RQa+VniSL+MG+t+7IT5AtiUf12TNmE5+//re2MYNNXttMNFf0JReCWDM2uWS3qVpmGBqZztrNxiu
U0v8IoQV0GtKu+RizH4NsEDWoUgYIzVVvfCPshmsfBaUWkbM1AdvBEFdJqXV5GB4eMPIzjyFvKyp
asCzw+EhdIbMKyo4JBFfMiULJQGW8P+BSKDcPx9DoJNzzM1S/qQ05jQguaI4eDUmiUT2nR6hsktx
jkDdaY8HcOzWr8LPXtXoMgJKjYZdt22YzPgpnRuYBus8aQYgCbwqgkKmtW5cZHbYnv1lyXW1vm2/
44M9bgCZuAuiCiVFLfRMz0FpSKM4UMAf4MaiyWZRqjfZIa+wyw56hRArXotopKAsBpnO29/YgJJm
J3tu/u59hdpxIeVtdxMa6hVG02aeVOYkCNMYjg/9h1YnSdfRZhi2zDHsLed6Ya46fUFrGGYdD1VE
kpii4Bjb80SxDCv9qC62dhuTUjdtcPvR/p+RPR1NHI7Ok9eEZVq3D2v+uht9xDjyfhMaHaN3mRa7
mRvVX/XiWmXy/95mkg8Zeqt2W+6+lr1lbadgcq4sMXgkenS2raWw47b/K4VCFr+1OXLoks22co99
2hgtzPk6NTCUTV4d2BVx02jPzaflLoPTt8q+2/3y+bWr44V62TaWiHB+o9tMyqKY6ysVc8pmU1q/
aKwVltCWdPoX8objWxtHoGZauzHx57RNnDe5ONXH/o3RkKUFGE2FyYbcne2D5og2YyK/KzPDkw0X
sSnCcTfIO9atYyYQv8EPBF5K3nU3h9mack1/V3uaRfVtw7LIR13Ippe5eAy+qiYWPcr4xAphB9S5
iLL+PhkskCOAFQH0BbTtAiNQStGxSf4cxxngMNpGTU9FL4D3D5wkYsPmYw4NkzvGQgNtwmDRCyBZ
YsmRQP3+JykjJr9g3asDC0O5GtMChS2bphojz7dIbmVTMoCG+9l0U2qqED1AvF2r4vqBHFaHcULe
x/I+8YWONnCLtttuRKF/mM63x7NBHoHWm7rsB/laWvF8QkB4TuhgvG6myDd7c/bSXgcFpqFAuTgq
KL1LBRWsLYjJnZLTe63EPxLarkSwuMsxlBn/yj8nu7ny60QaZaiCJinCDDMyWxEkTRR+5F7T0N1q
+QghSlZ2kZXTP4zSUyIbTlupb+r78Mf3eRK2UXVKY3rvPLdpImBCbnhfzZls3j/fIMPu61V4+nc2
VE1pEvI07vZgEC3oVFZ12Bw8WyPXYXO+RhzBsRjpHsutsVbvKr+3CtE5et0sIPHzR3R/ZzdgEJLu
w2pAPW4azmLCVESPYcbkTMZKm/m10PhXTyF7Z82KypfezvSoIJFjiJ/9mEZhUzz9ioAxztMzL1t2
RzRjiXgLleyDVJsamC/aQCmLM0tr3c1b7s9s+WPcjymiBE8Z7jV8K9q+5e+hDGdyEAJU6BsXNi6x
QTiBs4HAZgxJaV/YV2tzhI//OPJG7/nkmxOlM/z3KOF3apNc8fHGYGNHDeJ9iMz0fGKi2hAQJLCY
FWdl2wvFMOFtLcyX5DwFiYmM1nqpeN5WX0gDoP+2gYdX4NNB6VVjkVM2lTvV4e23Z0GDYd18x4rM
C8VU0Cu8RsW/pctP2iREuNccHqGruSpOImHB5zIs+eY/KfOM5/h6R/J7rmuUGqZJL/+GrlgsQ8Y6
0rCPXQJUy5bR1FJIw2zi9W/ap0M1ikvl46XPGe79oXS25G9/oHwa7ZYWiy6Lm+CBA4lBx4n9Mfa6
Ec3Bpf1kEFdKCK+4LtREwYTOk2ItDQPOdQGaMHNXQZulvnGp4HK7XQg8TVsNC/t+HxLzUg0EwnHy
Jq6SK5vL8e9GdyB56+3O54kc30ZFsZb8rmKjUMiJchM8u65eqsSLPdJn3fMWxnqB/8kvmAIiPcN8
cxx4Fv4LMP/w+HDpG88y4+kgkvDrM2DLicyX6iVJVN2n9XLC/AgtK99pVGGpewYItOXjzpqQ/72M
JqDLlUYH5vJxp3oIHQvTate/X8UUaBeJyc0vIJM5/ng3pxsOCLa93CLCSp1xcKjp1q/AGYBw1lp1
KhU68tpP7+uxs9fnlFibM+cSIhuvYIynlZJVDvXfCM6hwugj6r30ZIudvgiBaRha4LZgkMvweLNJ
7q7PSxMlpi321jnTgLAZOqoC3iQsV09CIr75ossFTN7dTjAhQq0FWoxDYjUg/4GHWJG8u6jMjE6O
jiZrSbJ9qZ6TQ+HO3W1+gSwQl8955YjDOXA/XO66e6m7U19H8wVMjZsKnxE8ZdGAjd5oIpb4aBu9
GVPC0gxyk7aMY3aqGW/gvSyZPWu8zQ5QSHG9mOxblrf+jeO0HavXob59J2x94Md+w9PiR6Zky3H+
XfnpsMAT5hv2P5ohkMxUeSn/2r87Wd/ogwvx8WlaNzdfC2KIri9zLTC+Oyf9x1lIyBihbQcv/egN
d6sRXmu/tVHZXa+KV82C6WoZsCFHjKVxCbsQUbpGxXDbC+gPzDq2zChtVdIR4yJwp7Mr+wXIHdLl
w8ZJp1LWOv0Ye5wMQ4NwSJS4bwTZHo87t3MyZO5rLE2syUtlSwW7LEk0hh1IOafnm8EXZGbpspTy
x9pNewNbjQVBYeME9vatJ7A9J47EORISyxC9k4mMuyS6/tPnKovuy6Hsp5VRm/xKcTbX668szD4c
Ff7RnL/yPykDsqhf12yW4Y7LkBpfTPS79d+UYaxLu5+9+FXCaAffuapfPGG7ZSqZGwFNA7D3NXhM
wNi1S+oxgcCGHQUYrHF1LvYq11VPVcKrQU2mQ2Ejy3tUTRVTiEys8/378FQ1VDKnUbZn6LGZIN8d
2aNySc6Big4kdzfKUePtIkDwB2qLQ8p26WZf2HLxB0Kg+dOOsmuEzeOJGJXwmBO8/GQH1ct7NwNl
bWMAsbY343kbFfa/8gKczsVcFKJul9g2wser7SEptGPKys8ugd+nw3lVwZAA2Wrf03wFnhUhzoGE
mLdIpoNKV57yemuv9kL0xs/qGNL0LJJsnV5yOWZWhqLbmXOSdSAMh/NLOlUde31PlcJoCsp1y2sl
IT6nvAnEx3vFlMqJP4bh5KS7MSmx4b193M3MdNVEyGx265BE+OMfOK4vmde/qFdfYJlPlk4Ff23v
kN+lv+BI1AdybJEWxScieet5P2qCBWWQu/yvSBxzUmnmgGshnM1Lc2udY6sE9g/8fpuI6ELaJEFq
tCtKyi0ZYEXgA5xqVEzbGH9bolFdIdwD11dmq6yWLek0nnkSYxRIfEBO8p/y2nzg4E+TP6EtLUII
B+0thokwooJT4glPQYNqAsgHHgf07vd4gmC8wJAt5ttzsXbXaO27kBszcA5cRQqCACinNnBovgiY
QIg2cyPIV9W9CSa5Mhz/eoOA1oZC4zYV+Q7UsflggnnsHvChDHypzIwLr3SlfxWN+xw3QqRFdcbm
Jk0bpUjgxr0cy5oJjEC9NfOJk52BvXz52ayIL+eSdce3j9dV8I2GMeKG+Vgj6f0Y1I38gcoteYJ8
7TVYimCgLZXJn3ryJq3QV8fKNjtWmThjdujq8Rwdk5gL138zmhh7EnBeRnxl9qNfKEMIsDKe7QjU
WKtmJPaBs3X/TEAyOkHzR7xyO8+b9Z08dxUsrI9YMwGdLBHHJ7c1Xbww4506c0A2DkwHwxbn1vzS
jLLp6sHEIeQeMvnhN/lwHEitSUuBggwJmaR5cYNV60e0WJSYKirIZ46cv8O9KawUS2tpFRu0MIp7
1ti9Wbac1XMk3BB/a139ZUHiPvHhXBBpJARbUzPntCqmmzNKMb1KY8EXc+14wYwpNzWESCt3/1Q4
MycMmyhsvbM9/hU6luGrqHVgDDMDT9NLt6OoF5eUBPzM8XlFo2XdAVH68I2wWzpm+S/SPk+daWI+
SA+2Al28xR6XAZDeoP6K3Wfa6Y3pJHnpKtIygKB3gfOTys8fHVbbP4XGDveahsZzXsFUVBGc0xxd
mNeEIJRtyMY+eQvJvWExNQXzXtOaFk5DDUgRqlZp7T3L4luA9NCjZvFufLGLM7P19jeHfYpcdgXV
6/SfF9YTJRkCxSSkYmLHA0atmUPaJuZvBLI0Rkae3KN924Pjg602FosBvYVOk17kVVrU8LowWZtz
UvKX5Bb5T9At+DxeGScjaPonJqvJM9xJStU7tFuMpRvfrHFJc6WOrijUAQCthacwzoSrRA871DXU
HgBr9SAnw50X8tmmGzNq4r+TVRyjlP2suQbjuzxFlrzVnN75va78uTOT/WW71t1JNZOi3WMjDPdr
QC6HxUZEdA+pdDuEoKF41zxkHrBIq4vXJQUaagnLMz7/tD6fHjRPFoo93/2yvqbNlaHb7ihAgAJS
EAHCUmkN9AACwPu4TV4BVnucHiCyU07HRgOiuMtzRVWEtC9pAFmMUsLl7CzrDg+3PnGhzgXpT/Iv
cqsqHX612vYX1RuDsvpSdpK9YiPgvxuIbPkpZpaYQhgwgq6jFMxYLBokEk+EHuibHV59DsZL852X
s9FL1h/GNb3ZZFtO4qMiC42GmtM8N+Fh+wiAZm2qHovCrbZrxSXpBpdQ5KVsC+atUD7picRFG0Nv
zMMvEXl6OVyrzJ99KLiE26isFn1nYjYdSq6ZoWORFUrDLys/5UOAhlzcCUxnwcN7yqeu0gJrBVpm
GufpuF3M16dr7xj2vNMq/xQQqM7Gr2J0nCNIKDAjsNAler6luef3NPXTh71nmskHREGy+oWL7hvD
7Sar4WZbL6Uu+Sm9nBJ/awvm724UTXbgPh72zEjFBeyjRNlifDyTLB6U2XS/2I0gxtdf2Z041Vzg
a2JEanMGDc59zYSTXPgSmwn/fo6IP8AbjfW1VB6S+s0LBC1AnikIxAbCn7QuQt4ZaFAOxcLJvI6C
l0i9l+DXwDyWh9AXAEBdbllItpLjqxLiLYyVNcLPFOBbJ0KwMpW6s61fypcT8PFJnWmqSGewxedd
O791xs3F4Yo7NqORjwK+XfOvr0GLnKcn1VwkHy5+EhpsQa4o7rhhQrcHntWc3TBQ21jc/La+o3ln
aj4PK3HASbLVb3lA+6e2stwCiiz9xLmyZQeWIX5ZVeqsMdo1es782wwY2GmMd/HQ++ji04S/V9l6
ePRaGsm2JN+kDoMKwHZQSl5Hf8TOZ3yCOwED52nyO1WSqsiOn1s8E6lygNmLgvWKaNpsrhRDwKH4
SlWQOVeGaJjIv/nLdLIQzabm8GsaIZw/dc1P1KDcbI6BGJtK33SivabQmR0POQ0UhBmPmx7OOV4c
eFtObexH+g5w+Z4UJp4F2aIEpnl87/M/DDvJoV/y+3DxbKzYtaJ63EHJ1665m1wGaNanAWfqS+KA
rBeAkJWSbovohUS5ciOEk76ssb1JFgklV1vbYvNU5PFoIkOJrWrXQ6+Z/LJJBcBWZHCzX1SgV7tp
YOQsffQYt5aTmDVrv3Bf6fCHI+ZOZ77QIe3akprwyiVM4gAvHg27511NJcmLTCdWStCVza4bUGj7
PUKYNu839/9hBlB9ZHykOJipM3jLz+BgmuIXGd3B8p34EaNOB01ojLgs0V5tvRySmPTIQzQ2/JAQ
CYfRzF9C36ml2pUlG1IKSq3JbycKiJBsW9c2ZFJTVM132M0UL5+xiTIQgwR2JuFEe1cRF9yNK8nQ
hGXW8u6E59AhGuCuAsdwYdx+Phfle3zJ9d1OI34IKTh9WXV7A5JVOHsdZ3bXiZl2lWTVzVFU9uNd
OCDu4Qxy7TTlIWkGrIIAEp/PUsmn4FRsWpM1m+1A8Yuz4r73MYPDpRWWhjCrtx5koVCm7345u39Y
HQPXT0Vv87VWW9nI/LZqB+PwO1y5PeFOnemELlwlNmWeO/hJ+YXXrO9fzX9Ffztfwi3LZqGRIy3L
7hVMZLvFl7dDtG7OV4pPuFpkL0TI6FugfqueizDdJLsZbYm5HBLyO31WeCaM6e3aYtFGXSTXDUuk
3GnAU4Bh1a3/AsUXGI43IP2YrJ1J8QVmwfglRRFhVGm6r0s6wEBXWknTkJh9ylVuOtdXhpZqshyZ
F8aJIiizGwdbXpa+Ku4Odn5rX4lEIqDkbvR3flebZGkbmjMxtD5u2i8aZetvAzUqVAWRQ6b0audx
FLfmRaF4kJ3tmaA2wEFJCETlL8G2RT0GttquqmjG43E1DrKCTYbVCB2hUWMTPGZeK9PIKRTd/gaI
78ctjYWureH9OyZU7Ls+l05wm+M8EUt6mcCJUadQOXhmUz0gxI2ZjyHGQIJLjiMd59yrPmywdYff
HUDxpUSP2tH2Uf4ELENQPL9youTjYhMtYtqq+jxjaM/Zv5Miw6d4N2NA1whRQMp4A5FI7Ho2GFEH
qO/lzNkJcF/3JJFn94LlkWzZ1SzxLzbN517MYib72/xo0ZcjQ/BiuCE+ymATzFxeLwQVp0udHgy3
C5uRYZlfMlQcEiIhqI2oIHAa/OUikkE6HYXj9givmTyMH2iLJsd7lmI2mu+6umkQ6IX08AGevPy3
E7Fd9Akre7fi0bPJEhYXsPB/9BYE9SGhH+KKf+vMrN74unbgkuZofFz2J600CnQZba+plbxqjz//
BoLJDRpQGV974X0/I1hOqE94iwS2BWaREU9le8NW2eaIlXMr0lMy2UjQ3a3hY1VcsDCt6F04hBjN
ByYvCqGyrQ4ZxBtrCkdvk+zOYxCSOzA0gVTOtXWlHwx4TQIO7t6FRlvQIiVq7ZKb38G1cinFlSIZ
PcuZTISkRmTvGT4y7rZWtAjAGvAuwekkVJHvX52Y5o5DDfIKr40/DTTR2N278xVjCnCNdw2AA1v7
R46RgPQJL+Iq3cn/Iejv2l821z3Ex9mOC0JoEdQWxvRKvVbmLBRSOFYFMFO0bauykm1rkp+1vveH
m4sTypWZHiPLVQxE5PtEBDQ8LIYVyrz1NiCOphCgxV0PqA9oFeCG1ilrZwJ0E0A+hVaX1e6d/FnE
KIHsmWg/oVOQGLquzNt34l9BNlKrxJ9Gl6dhR4yVmIVCl8fP3TFeicrnNrl8zVl8XGnTcb1KXsJp
CmvJEP0M4QxTEvEZCOwWvUN1TQA+NWxNlZZ7jKgL/xPStRa+R41lYNsTNtz7v1tfd8UnP7HZXJdK
6ex+rJN3siKnU6lYDkl5m1xfEDt8ZFd3szSM8MlZzulP6h2WU/p6iDj2Nyg0WZxwpe41i15t9LOk
MH93y7FWeljuKSH1cDfGJaIH4lK6vBPPmdV2fXrqph52kuvJO/Ul36B1wKqfnxiKAqVqyf2RwE+d
2lnLX00SOaMu2YvNUwK+vhVYZ5SEC2fArNBLIgEDqG5Dli/PJZq7ex0yglnEKmqTHRSZvZQV9Oa2
3SQBhh8mkyZx7Aa1BbR8NtthB+w7FP/DAitGiAyP2O7hL+unUhV7BtrvjHOjFBFQ1nRTCNP1WYGz
3T4EObJgUA8mNofMMW2GT4YvpTE/kwuZ4YSgmAbZ6kF1ndX/H2cg33u2nX904FlpdKHSh3UNfeY/
cHFF5Gkh/h0f0Xe5/tWyGSsvHXNukEi3wWB0vnuYaDx95LVqM4ZizBvZXjAS6Q4Ug4wvH3Wv7hgM
dM/7PbIid+w/IEVcwM5Q6JYvjC6yHF0T19jtEqdyZKfHa6EVnew9M1Y9wM17FHDnFLSCXpWNlnWF
VlmQX2j8wr+FNMcX1BB7CgeZqOY+XdTpwVj17FTjsnne5psx5QdO8te/R2Ticq0PRArUJSBdA8GI
+pL3qojstQi1HHkZXbPo5YOSyJ5KjbR7qEmxY68Ahv04SwCT3cnsaL4mKjUJMMBoW74kuxbF7121
/eVnU64GzOSEYguJW/bhei1vEWm9rTbI23Wx0zOdR4Ahnhp0liarda+C/FZxcU2haZPDhZQS2Emo
j2Cni0oQ3hc/2+Jo47d7bDOhscM7kx2MFndWi9urc1Tf0y6RqYCxIjIVdZxWpT7lnRF2OpAuu6JR
HmLcC8yu21y+KY1O7/vfC+5gBVPsx5Fwz30TzeAVip1VOlbt/aPGmHXrWH4t9CdBWdnzvGqcM2BN
xp8ItcORL5lESEdGXn/TbD5GeZLBFWwSRZYb6TaNz5vYR/vlQCKM9F52AMRnjZ7cMk39g+v++bct
qJPIm7R1ZIHml98lWDwAEW92cAfYh70hC66sXuEsBbb0vTcLri4sdq8F3X+tZFnbP+FSSRwS68Js
X/Ca7Jja6YKDcnWb2/qDiINa3vdrm2o8muHlSsU/C68XXCaXmZ4E+mz4YcpBBikaiM96CjTYh4r5
W0YUrlpZKGH0ENqKMfTCMD0aJKp50h1zYTeQmaAQGcgCeZvqTcSZL19KeOv14/6RwIn4ykP3Mh7W
1kQh63a9HpqaXs5tdMy9wnMSmy12aKVNkVbAkLdDHVncrnBURg/AE1utUQx0kdldlSZTAuoC0iZd
eBq/kmwX+ZES+q90Aqb3LOqP9jAPFd95ZNfY52E8cF1NE6iVkRR2l/uogjZ1GDl5zXt7tyim0y8h
UD6URd2TNQJltyGjNRlRTtQGmx8wvwumutH1wUqu6HGwQeTmAjRtfDip1yVWDKYW/E10WuOb3UTo
f5J0IDThFcuMtFCL06X3RLxM+YX+LX1fR5jjk33wuLeZ/Nlm2Nj8NkYrVN0oSAsnaXngXGgRo4G0
RjNu7yp3ByeAbmeE1R+4K5EJ1HcALNRpkk36jitG8NzJyJXmFLvjrOxfUJOnQnUR92ujZxozGGKp
sAJzBhi9XxB2bug887oez1zBr1Y3qUen2xxFRgB/B8mM8xBEuxam+S9KBotu21aEy6bW+hMxdaf2
AZsTKfYEpyBY0jb4ZUGNkguJgv1bq3V7o1/zYxM9LHykCwVqMx3Rq7PsPpvwaLJeiVdwqjphTO9N
MnIMLKFgyKzsbPoFe/ZhoBiSgvQY2PBafJCCwVcB0LKEFO9sxhHJOTrjWraXv3cKEL7jPC+ESUsV
2veUsHPZ7/fjKd3jcZLzzx9F8Kh5LnnnHVMea0/fZLMYWJwfszCXuvDI9SJQeP0CVoc0niZdpoNK
oQF7VmRd4fPphEdQKfd67k67/zLVRp5v4ZHUsR9g4zNZzcE94F8Kbigv7B6sfAqwnqEzipZ5sfcG
EWu/BC5/pajkwvfqihseT7kMHhWrSxDy2FKz9Qf8fwyJ6NYg5Tos9Ae4r1bhON2/QGQU9Vx2KvO4
NKEiMlv+2XHFQB87J5FVe4Vaf4G8GxALKg7oFORESw9bYXxykaoZN1EI3bNR1I2WO015cVqSA6gr
q2Xr70OTe96Y1RInHjagDjHUWhPEIigDsTJk71sEdI9IkmU0UFNa9TtSjnHNuC1pleeRPQFrEQWO
KeqT+oHLTCuiROd5wuwG7KaCcfqpcvp9bvZnjomidP3Yo/5epbn5ZfFQtJWAJ8IEtB56ktdqKr3n
oyLGVmhNULI2s/Nw9HOu8ylkJ/GTDsMTtX7xaIUutAG5AM6YeJ1XRN7WVa2ijkH0JGESSXH99V/2
+lBzmKh411Tb16XwyGQ2U1ZXb4qdi3L29SolzxOnTKzT45v04wthIUpJWImQT7TygBU9GnkGCh5W
pgvFtIrPDCcOVK+fr1GSYN7Cz3WDp1n49+3SpVwTseYvkqSs/oJD+OCeTLYFF0ZS6sADXdn6Mmb3
2UnG/2ZUmkfx2ew3auVNGM5b0LBzxFDcYnwH6v5VseVPFf0+6pcsZmg1hkC9qXoqWstLHJcX8Zhx
M3P3HH/R2Lkrl6DvvkTbRw1GsUHfilB/PZZFILhIAsaEot08V27RIZ3wB2coyw25AWKIjO/z8t+b
MCLSH0YAtLiNuiXLBk4EG2kABx+sHa2OgGctCJ2FKx/5UCNttb1b/bRhnwhzP/y1mzy1xppY3Pgq
qWMR04tyLeym9fe2y6P7LOtiPlDbMoflu6XiWL6kxukdJJ7MOVMNY6b+rUZ7H9WmK5XMXjzkyIXx
z5nugcszctK7YEMoMmKNkwVqqhZvFfMBUCT4yOJ1IJPszViRu3cIXfOBBtax/1Ju7ht8C4Ed104p
b1z8agyY4A8xOjZGbexQ6veyCZzRbEC2wfXUn9Bk+0B2nBJoCjKNE/68fAJBDa4bZV76eIlXsFzd
SioKOSrmLc03Y60NkI2ykdztRp22H3yNOXFUJjhS3eZfjTcgKsqvi1+HSF/n5eyETYRqAFLBcSW3
HDksG6WMSGgg87VhK8Lu+qeIHNxZ1PR/bsjGQ1LvX3YqjcDNq0moDjEGseWSZgd0niaoBztMEJJP
bWSRKMSXL4Ic4dC1aIXqZpwSIqqPLqbs/QsMOKjDoYDox5b8MPph8Rsek0/yc5EiJKa+ENMJPlFt
z9dqe9Q8+y7Yyrc30Tk/19Cw0mvS0Ze4TrnSRl7d9ydyYYBwuuTA3nfHeempQy0hQGN9041Js1NF
8f4usaL3F8XHwXsZHLpxACi8RgBJO7LkjBqizykw1E2CFe6CzUb1/+r2UwvDpORU5VEzq/3xp+f7
2AITtQl+fVSD8B88Imhhx9h6ff9tVCL3ebabEyECJuAnVCVNo28uAAF1KUiHzK/rfI7JPkpZIfj8
D4MpAhNtQ4Z/GzbMg8yTudggxVa9F/ezv0/UNpidXdX+zAJH/BLVJA1excs4Da/1KrHtAGgTpfVJ
IkfyjMbzv31Ev+/QdUwfmo+MGMFQuCdXZMwVN4vidLTXse97TUAIlV0voU38oQHtVyY0ERKgJ/cF
mK8rqdRf/I7tXwzWMRlk+8/eW1tBPHN/iY5NY1T424TO8cn3t7QtJ+boxTsAVYqt+DjluSGrX08x
G/MPjEbgigOYohzXw1+eN+hgcw0myjaJ8Lni0Jp8aB6jyPwSLxSHACeyg5k6utLcurvYOn/e1DDG
HeMCxh0Pnr1VWkersbWM9d4cUPvgMPs/Hauj7b93rA3iZcfQym9ZetJSghOzAqVkQyJD5Xvct3uF
57VPJkT1rqQA88hk/pizQSJ6wPvQOd64vWGLURsq/KQ4hltt41Jc2+rYdZAwXV89G1yh6k/3FMNv
RVmpzeoOZTDfsDWwzvgxqifayqqOaIX77n1+iCbcnvx2XWYVryoBL6yiGdwEzHKEvjRSNqYsJJQg
ikBSj+Ujy1Ix58TQ5UgE+s0idcRIeBLuQWMmD4cUpAiKotTeI4XcclrsWEEK31eAGNVerW44GuDh
/FsaNqoXKAj1aNLIfLkgOu4e0I3vRRjOwLpbKL59nUW9SyJGqNoaX6ykjfUlXaPWDigJK3wpyBbn
pF4NMWxoZdXp7QA92bTkisbpa/7ihJZ3LrXYv9/ECqXAKi8b68kS+KZgiMEp8ruT9pIjT9uVuobZ
MPuGq7KSw6zoq+j6rDJQemN6DwVqx6B2LIWllpWtggCSP+PuYHbvpXqb+IBL0RXlpQheYHyKQwZF
gHzp4dnpHvYjbeXqagxAVbZFsTV8T+hYzmWRwnOMy855qdVpzGJg6iYuBGj3UT8Is6YsspJUpQog
GMY1WMR3R65dvXyY7Fpr4r5vuTCb2BvIL8Sbo6f96i1VNySwxBOOmywugWSHMcUQptVvFn8CT0dB
w2tWSwONmk8++XSjWiWsZLchIDYUsqLTV618HmsU7x4aaz5V1Yr7tUjiXR88IWqYy5aMjkonyWqc
QP1S1dvNE4lTKthtmXQIAd/yCuItR+VSyDDRVGZEGMBkx04GdpIAKkJsH92WQ5swRPYvgKF9wVVz
hNqQQajWejfl68JZQo5TEuYUpamziWB6FMEHEkRGeYtA0kSB61za1PA0XDu3Ll2S01q4gZi+4gRP
vEX7C6UXEx8vAB+L0yFFH1+q9D160nx86XbYLQBgffiHqwDzXLnQnwpHfOLNgk7LhAx71JNneRzK
JgF8zR8vk+63xx2j2yB+0GEIuidWhip9V7yflPaL/NBFGVUwRYcQQIMl1kXZZ+Dtoh9dihkY7ZZF
5EHh/aWl23rEbB90Q+VGyF8+7Ipq6KWd/KIt+m5D4+2vgzAd/qhXvGEJU85dZVh0ptzuhSlZgVlr
6Sezr7BYM54qEelDV7RLx5Z4L9yN1fGmf22P3zw48H9UvZAjH0wtuY/M3XnYgI6taCtA9MWlC1JH
L1rzcxE0SABNsRAszbZfKVgDTJ2L8unigxOrQAwWr4oGOpRBcKlIUvXQymGhZWmjMeOYRVuHjK7y
0EAfvDiUdx8+UGerdA9bCGlmxc0eaDiHmfDv5bZh0B7FC9q4rWEnF2101l3VAF39eTZffl7T4ck8
wn74KFvExzcwb0qx0uPcW2gO/IjWPWv3xuQTe9QtAPvvYTiKSy7qutCWF1C/mxrwW4aD1yvjxG3k
G7Ky05nwGwQEMEr5F5NDsv3XgxWRTRqCrCrASqa6IlD1pTexKhqLo/+ByQVNMf/dFkFUClClc9Ez
jMal1V9tQDZwU52jOzaSV2oRB4FWzaDf8dloxUnNOoZ6pE9MrKv5AvhP2nacHIs7MvFaLruzkyMC
6QfJIMcEaecgkUAPsYDPcL3G+No5VLSU+nPGLfSGCPQw1Ma/OvcHUbVkBYcZZ0RtPYWtdB86c1HI
9JHb8KjjcVESv+S3NemWzuqkk0eJr8M6n825jSfKU0ZKzz2wSdQPD9dj2wHGqL1ivuQ2r2rW5gGO
c79t/NW21ooDzGIzPn1fxJxt5IG9oWPrynSFHvdK6TL4z04rjq7r/fNGaiDEest2MsXZ/e2WACSo
Q8xf8hRYhWoY0quCMeSjkSojWg1Y8hdBrkvxZHX2eTJDONCGdx1OED0186mwOl5yvaF2bN3D3r2P
pQ6ID3bw6SqlER2vnk/uPjA9W/FOYSk3U40dL/aQOtNRUWGOroAQtMJVpjwBLDPZy20QDyV5ErQV
1/dhRDrf0zc3j2UenFuICIELHK+YnqPtg/MiXsWnq0OqWterdYV4o4CQZCl49sKqKI+C+AB4DtIz
2FLcw+8lb9eoCUw6zehZkqF95P5lwBrBwF706JauOg1BL6DrzmVYSvekib1I9/I5zZxCLsg06XwH
Ynf47mMVAld7Ahj3I058vEskPT9VxjmImxwVCCIxxh3XrVY5Wa9jhkawes+CElNU9WpPgqNTq3Qs
ej/YZdwsmZ6I0dr8RmDGp6XKQyuKYZQmDpsgvDEpyPK/lORoKaPtXij+jar+HfUUYg2kJspgQf0W
THsjpxIO8mlDnbqdkb0Fd5GeN7rYUhW3ms7e1bZUbRbE3YAMhl7HIXZv4SP3jaei7CEpx9Dbie5z
RVp/2YBo6eTaRst2y0dyhagLoU73qHZm4LLswCT45bmtRLG2P4FRZ7zBifaa28rSxlCOVijbIn7y
DCzIc5fpoJGI8EUnxQOK46GhFOriHdQ3dat/BuYBHOp4UGefj7zzSvmShO/DneANsBUcMuBwa3PD
IHjuZqtf+rKPgrJeaQRNDQX8GoNIoRNh/Tn+A1Iqp2W4w4I1w5ous5S2JInQ1ZIK1hVIA7nWbNoZ
ea67urFivnsJyy6lvOqFKDW2Tu2sE2t86/sQpCGLU4/Zvrkc1ts2aYkEOsUFdwnBpB72XXhgA/9u
bezgbaLGYQiR5AXpFw5L5CzR6DMOzWvfrxua/Kl5BetD/fMRqcsyxjnvVN7tRomwEQceye3qR/Br
4ILXtqiZ/Mi17zlVOvHektaz1EqcOM7mq2cROV4jawTNtZp0nGsGNTFEsqkK9g93DdbticLh9zfX
Q0rqFXsI5Zqi0JtVALWNldlJ3FIdrem+RgcE7S7ecYezDKSbMLlYhmcb4ApfUciywrgTcwvaNfU5
TULYkDpBbxacvOlWyZRcM9CN/41dABLN/sAxPZarhi1fgX60v7DAXZjSISZTF2EbjOW2+a0bbB7k
sq7XhxNvp3h9man2ultRxwqrzDSijaYUpDfnl2h3R+pOM/f3kdVk/0ngq/bLib02/6rLJPe2Mo6F
r9hz65MKEYTTzWd+fuaPD3XyVLFfDsEwJCLNhjqXVOucEaB22EWj88j/FCq1agK4FmcczG/BFW8g
hPTeREpWRi3St2PZIOms/kvLqozq2eeJUmpcswrL0+3ePgKdATCEd8EE0OdYemCDDY3gB7s+NlCX
T0le5uEmE+9zWSj5WaffqMM1Oi9fttjUwOjBQBmSpmD5D0g9vBdShR8+rNL6k3XSG3xkOxqQnQ0X
AKKBLHMwL1dwtp+hGrf5S4O1HGRKu4ce3d6HVpGzcpVQUTrXXUy58pLaSoYgLhpo5yFyX5V8rqBA
t9JhL2rPLq3uPTmQIV+ZtwEDi0N3NGdudSbID9hYnQ60j92+VMTOYSPaGkSb8a8z7xgORb+SPcMM
GJvoKcJ6McLwWLftk6A5yWkNX4o+HyL6e4IIDUpamMlm/9e6CxDAJqlayPLEiOP9VZEUxCg7jZAr
72M3Lnp0nPU+dJugR2XALaGn3mU0dpQaX/UpF6rHVFvIlEetTUGB12oVzljMuBrwH/pc2YZi1YIH
DD9/CLMWdmEapZozefesWwt7wK3q3fxfTeZlN6zb+jgulQRngQzU7eGuCo14uYYfXsl5Gd169u3y
CIJPznc6Mg3VG1kC7/u/V0EaPrBDFgpDvlcDzegU7tb9G+myLR7EQHY9qrjNnZESJG5SgIRd5tw0
rO2IBnL6aOHfCT25nzRkGhhhZ09hIAuMuDoXsHMr9tfCJ7JNcY/Ftwpy5LJ+mDvvoPefxeOwUu+/
8le2LLYJ4ZIChGR+opk8AB3ygljB5Qnn1IWMpYHBtFbAz9d/r/rypi0Coy603WQ4k2nVZ9vS8dnu
mRALH1sSXYZCvSlSVBv9vL+dLAnGSdTcEvnj+kkLU3ps4+N2hMpnu7FhIh8Spk9RYo8r2R7Z8j9l
z33DwgPR/2wygfHU8GSCq4nf1MNq1VRrMghOeVt7MHZLigdmUaX7/HRrzPd1dEkwij1AkviEKGQM
3lFsYufC6ZXmg0Fq63S3oomo/Y+tJBR2nWvG3M+3HWagIpnBA66rOYQ3i7CPVQ3X7qeS29i+iKdG
P19BOSFVEO1VFwzDMQDd8bne/1VGhcPuAYq33aoQp9r4A162S9sFhK+qHzobQ272XsuedPswQnsf
mQaPxvfJw3JyccnA6VrNVw/kJNeE0ncYZ8vh6l0kROi6edU+1ee2izSFi8txKMyNvg99r29QmEV0
9j/gaUxdgyZxlinb3WJs2FotqavhB3ayU20hsNAm0WtNds8QDQNon9xLkCRXjMTWL0+x/VazPhWP
/F4+y/7gPWXyZv3fkAAVdJ6Hqu8iPiU5mHU2Fr2Lf0DL753kc53uOfk7tiLkwOYMu7V8JsWjnG/a
kBJYRjuouyk4eCtGLwAjUbaeSIrLq02MPVD3df/RKsjkMTPedxRQUGZ47wG+6mqGmUsdgvrQEfxO
7e1YZLzlT+Znl2co6FFNPuXcW4AZdKXQFzVn6nWi8TphIhan6SXM7ST1D/zTVnEd0aqdpA87p/V+
U1YHlWxLk6Tq3faKFrgUtrQIivHmieTMzoamVN7GqSaSxMSWEiU97C752iTXGoigVKhGkKmKevEB
RCVei3TNxi48a/6R4VxmV2glXZPdpX9kEJwso8aRRDVWJl8OfvYLiC393hsiT8y7O3Q0ANdmvZmS
gcxqoaz12cDRvwppUfv09tQ+1wZ6v2VbHeavWe8OpPtgq/lgo/dEHKbRRCb4+DE/y1cC+pnf6sbu
YtBlYsfKLONNrYIevUhfGaLtp73RLPxUygcBWhCgRt0BaUp/FY3MD+0D/4s+0kuVXWJTZiIAeDCQ
tPlno8avPPdTolvsywZqS3jRwHZjAM9vyYHfdeKNAMf72nmzIopuoGo2jhS0w6Y337CHu0uz+mk9
DYJ/N8EuuRydZrzcdrjX9PhHkvtUZEMbFv5PTUtC/M0GKISJZN1nZbXUTKdYTC4UOEwqhPQyANve
m5tuyZT9ZJ+L4EOcIHbJ16onGBvmDDwGJFc4C4tsrTnOaFt4WsaJEGWh2il/1jitYlrZ5UfJAU6S
R7QCgruQtjsnvR6CjckExeAFfcXkJI2JQjHFAaW44c2nu+NvnAjaGoyamaJmGzS6+z6iscrIPmHl
87Gx/tHXOJ/fam7PTE5nJ81HqJUmHas6hNOTBDOH+NwQ9GM3xyj8YCKJcekozYiNdoqMqRblUIM8
yDlq/u9c4J32l/n40c36HpP94mT9NnlZxImR4W9wuWaxpcl3Tvv01TSZKer8CKPHjLKBJXwReQ4u
5Ud64DuRBiFheC+YOe5dWjC2iYWzD8oJvTIha09icNJZYGIeMPsrMGaigbhMO3lOX8peJpKeZP6S
m+9pMwdWWth74Icy+H2GcOGxD1RwsnUHRC4nweejciPzLWPFODmZxaWk86h/5zPbSEqZYqt6AC7M
MKfiCquMWGoTXtsfyd/l+TejZAIc9bGi2pG0Op1KOVYToGdQvXLO1p76fc6kioPEpYN0U1GFgy02
kG9ZdPHbcCyb6hyAmqr2Rw7h+hA7PkHANhZHuGKMT7A5XRiq4NIVxWYYsZhmS1WQXZxSSWPOp4hr
wrTyQyGRZGERzl0MniIJsySPJn6SSoI61Gq2rsVyWKG8mgN52G29BHyKuWVu03vFns7+YIphs9US
/clEScrpZ9/ghptGe/IObDCNoy4rig6vWPYf+cYy3SiVMme6hBIjrjzbEgYz9HXuBlb/mpg+SJ+P
JxRjUKfvfkNNadcT7lnUsMARJ8a4ZVgjGK/P1bAX5yk4B2OclSv9CLmKR43WUWFhUq6tfHGJPM8h
YQNKWAauMipn9yLGj2RPml8+jza46dDb4poq/jFWSn3Lt9R4Xu1x9BNKVVouDyjv/hyz1c6hUnPr
vdfGwCJFXqjznHU7uqtyhf0mQ/eXWNlnn6aqm8KXuZRBtjiHcAg5Ty5n2/me03B62gAf8Qkcgh9S
rbqQEQulp9UWoRM8Lu5d9a98nXimLPtjYg3asajMYcvIyEVB+W24PJ4Hp7qXmoQSSG6dLgr26ZQP
TOofTFgLNigi2YtSJ0M9C1Vg2DRQrFXWZkwRpOMkKZV/yszTdDOjl9D9RzbRTwWFAU4bmXaMpFCr
6YVxN02eAp676l2siQik7F+nhDj48y619opMGbqMf9Fk8XBa5wj8T4Mt/mio2ZCgLMeqisW3Zcj6
+3BR5yWVb59GTVihPmfNvldSYhV5ATiAv9epD1XB7gfSt3niWDgjoVekxwV+f5YEurJE5hh3CCel
QLLhErHYfkXsaAtPeGap3JGCEapz1BM5e0TF4dhMY5kDtzoxlhoi11TXtTPeEk9JrfKLxh6xScyx
Oel3dGehb7gdys+1ka1zzD7FT+wH0kAqMZf6du3JhaKxcML8SMcl5YPJkMnE6RTJTihcdD0nWGzJ
7o5r19Ysh6K5fKgaU/0UtCRmFMQRKfuDt/yFDguwTxE8zNo/Xdf2TP2Mq1xGQeTGerO5TmWeIfxi
aaOBO7gQN8hNTW6fpayx1AIDqnV32LblFmhoxHA9vyG+KrBPue+RnnENTGRSlfhbcdu7doHnTfU0
4YJy9Qsk8xrqLsGpKZc41CjmUy5WgLuS9Tn7cOGzj3jf/v6iXnL7eMvWJ3YvAm5+AJEICgils+Ho
ZqfTPpOgAAojaB463D/bVy+E2Y2P6Lx4N5AIs/COfui8cHXm5zKTOUUDe8AOoNHQTQO4fvCPpPLz
lD7oRWhPLvPWW5EFfoNWv7+93beVNhfaXcxPfz29MakH9te4tT3/ZoP/lxagBQ+ISTz4XILbJoqJ
ETJEWBjtFP0/Md/2PKNe6cS+lYMSJxk0jKZSQzMLtoM1T0Sz8E7Bz9IMrHOilm5CSm5IJbIUluxC
jGfMFG2OCJqhJXAJUn62n+yFGYsVgoY06d3JadLGQcCP7N/auEWzlExbEILFGGdWyGHohKbzXTYL
vWeZzHQONepqW7WyDr5zIPKoXd8tiA214acbcUcwZIayBbBjiGaapPOnetfgppOXnDZv/Rs8cXii
79UZ2VeZriWvXyV0hAZflUY/arBh0Nlr/IW6LahnFXifaa0sJ2Q9fgm5b2MMGeIjdu75wv6o66rh
8HjycgqaSdhvExuEPhFc5yu/kThdprA/SnYbKPqMyx4YC+LG5JzvCjNosa5degug3VnqoFhOGTUd
pAuIADJqpEW/E82Qs4rfN5tRSPuSaw+hEoTe4QZPHMfKjEW9gor9aNFzLnEdgmV3QIZCFrsI9CCD
BAFSGkEbHjdgvUhWeGprRx1hy/kzu23PSE3ZBcQ4D48Frb/0qoWM1IMnBYbpevGfDAO/Acymg3f+
Wf8SSnRYccRERgPT82NjX5Qob/oyCI34Y+s7v6GgG/imQv8XRgdelW3nbv79zgkxdtgLjMWWJJz6
4m2cLCk/SWkiRCbhGiGTsHZM2zqM6w8pjBTSx86d9u8cur0jk+TOMYuxsYS2J9uxc4fIZzySdsvS
iuZg0i9I+yAE7v5eEEXKS4MPo7vaFzBCYpk5ZK58gvPzUf5ydZF6Atk7qqIoUOuenmHMQIs7fJbn
LGvOJJnr/1CeKztGera6t/cnRKWQM5ajOgdfWtyHBd/HV6SJ1fX+gewUZBrqC5mhWZqqu54haF54
gkkCeWYEYEfqVhjcwuJIGdEZgvqrkffjba/br8ZlflBeqFhPMyLMdqgIvqmvq5koKR9U0fGzgsKW
Y5qkZStFuUhdAEruWwx2ShYN9Mv7/axTRA28BhgWPHOTFv0VSXwww0Z1GAyPr5Bz6Ctj1y6a1Rjz
zI8RsVBomWrNGaqDNJWdJbgABTu/9vlo/JfHboLuqA3WDVR5XsGFEAHhz2/Sw+6Z4CRanks1ukwA
NEvWGsYljXYyN+bzsL2lQihgfCIKX5QHHJjb0FHKqa7WLQYSHM3VZSkYMtDvVHTkpvt4Sl4roW41
CCq6jgsLMYmM36vqDATru3gYoG1wjBk+7NaxvALUtzMFQYfoerwe9Cisrc+l48b08Gb4Djqksuvn
K4JN3jhEnbbA7Bs0cF/hzVV4Lkl5smOmQnjfOxw6SPYKxM7ucUpZUPz4Kw/V5kbdaRoXrVF+WFRa
OMna/+FyfXQiWEv2pc2RvTF7lhi7Fi5NYH8CjZP441KqhmSrgbePqqy3baweVfUj2BYtBQU7c/QY
fxegjVJ/Aeuedjk4iU0/FM5xIxbqAEqdG8PgY49xJPAZmEZQvaWeOLvm8x0E1f4U/njNYkW6h7TR
MV9948qNEenjcfutFdoL0iK4eUJgOx/acJ3gYPDpkBOsEWJGaq3DstfPRp17Iva1EgJytyJFsAVx
r5AL0lYfHPaHsh/Kfhfbis6Xdw7GSN3eqjUoKp/cgxC5gykg71iVWbPaD2zcKHhn+JL4HCEv5qVi
LaVbS4lODhJd21sGsqBWmPThPygwEqdKbpO1RCcrSyoy/NzzxOGiWl+/UaO4SoonReAqPs7KUBHY
3QlAxOk0VM3Pj+7u8BYrM+Co9uGxIQf6kLj6RdtUVbvkkK3G/Oc57nqJ9DcewCmAN6Gbi65RtHNY
qqD0fI8YiF8ymVQhfrWCjmc3WHHtLWM7S8yOw7Q6P1jbDwDikt82CYwED4jHVvBV9sH5p5GATOSV
sMfsGGESb6VWvZ7H/fuLxHZaNQ0nQu00bJgJqrVBwK+/rWuDnt4Yau8z/aFhLQu3LEGzM/jJBFab
/PzZ0WHrUpR6nKDLiICZkRy3H7ECn4zBYjz0QfR8EG9/GRVSAbwmhgwH3ZNrJ8EnNXNnXdqJSBeT
IP/1Kg6STS1qE89k886bnxytB/HcQ7ZSMa7L7DZQpuUTf8vJNTFenYW6xanmKdXaS6JgQ2R6ifWI
akLDPMK/bdpgE2dFIdbll4IKjiKTRsWe497AkqxU55GgjJPkw2XjLF0L/L/bPxJrtjF7ds2H/hUo
DGja2vyyTmlWwWDzGvMqyatkLLo6RE8Xwtgj7mpZHDFlrtCCrLNeacodHDnAu4fyzmWr82al8S7H
fZXquFGhPBxsMFqEG/4Fc4thayc6jVBMjB6KZyY3LYJWn4oW8he02ogwRKLdhsa6mURrqCzZ1oTw
f2521ZSGXG2rpnP3+m1F0f+X2qQlH4S+2ZbSF28BypeU+2s/0TLgnNXxV9vgKgqndYljGhYD/htw
5rpe7QW2tCJJ7oq0FplZxpy8XkJpYJcwt4Pzi3b1EFraolYfzlprGVZIEYnEDcRKv6XHDoTnRcXF
FNGvDaQkxUyqQkOcDh2ZEy74doAlh/hDCRheK8J6rOVHot3Snobz3EK7+/ndIzRJtsvuYA2Nr9BN
iPV0OK8ZIBl5mkkkrG3mGDv1UULClAGjMqBqDQhcMzEt8ii8VY/LX49ImegD1CkejcPoYj+Lewag
rhsr5uZMH67GzuS3q34Ijgk95IACU3XUqVm0iSMVXhwxE3Sn0qk2hb8/8GiEuZ2+JYRi2pSNyW09
ekRRmlyh1Q6wn7tdOo8G1vCw7eRSvkvQrk/m6Zu5oBuRxHRWGRlaybpjd5ozb3GP9/SGp0jrUagp
4Kfkz68yL1eE+FnzVWW0hUPij2CNYGRFrrCGfkDm7ZrPv1qpuobs2ZaUlnrt4zwgyKmcwr9QeCyg
2ZcnHArbpKH0kCA5xOPBnwbUiLI62KS1WlABSo/IqipD+L3czfsvcPK82Dv/gMs02OYmTJn3R2iI
WreZijdYDLqqvF/Qt7Hkj3wftSp+PLQQdfzvE1t+LuGAG9glPjwBf00cFSp67dsGESsO+bqTUzYi
M8r4KWcsILophL3AHuZNf5g8xswe/RvVPoIQ1oiRgWcwl6x3d/dtk4psQDLgxywLRJ3NOfpPJVkr
rr3qMMQX3QHQ9LEYP7vgkLk/wFgU+DwYJeCKnA4VEriiH63piFkhdYoBTCapvKMspYsocjvx0vOO
IRDrd+Ofu1IRQKgKPUVV05iTasDj74nCJGtzNRx3dQMOXpSJXNSScuRRjVV8+yHNiZIC8CCNpdUM
gzV6Qao33ZiP9UVXhXLB3OIUgMdmGCznLRhuZO1foB35LWORjTpxXv5DLt/PhOdDdPDYYoWEpgnJ
qej5xPi6DnE9kRpZp8xRu3cLZ+AjSBAlAN/GTjedCgHtnAgQQZh0KBwvHyF/vKAPm7RZR6fTxAVY
JI4VKxd4cNYMQSsbD34e3lCkmjwAvi+hsPAPp4RXtHuAbMcsL00jW5QQmwfG5askdXqbAH7efVHx
ypqPbRN2AddnE3pxGGdCCot0/+u2MpmZqQbN5Mdc0zVSWy39zt+zeEY6T9nmbBw5qvVRojitKxgG
gfk2/u9Lrl4w2n/5i7z+EcpKO7ZFTBXrN978OdykDCCGe80PqtszZ266IzCdWyBnU+v36cJx9GhD
SzezjC0/KDIJ5l7uY8IO3SShjQACD4eF//56oYq3nFRZR0Y8CYQDrVvHQDRtw/VARlUmqAUYTBFW
HMnAvbnJL6tDDCYah4g/iRWAQp0BuC8/fVBxQ5W+5K9AtgrCKPvuz/4hUBVOK58KdVFpKjBBXTB8
kYk7JBF2wKTKus3lET2YY2Q6Q0lrmZwzLSh5VwO7gBkusdstmf+jO8lB9DN/HtveHK7K5sdrlqvO
82k7fCe+J7lNLN5LA0PNlFDIWufYfWu4GZK4hzzvWq/6Ld23IP0fJoR/A87Y1v1CgFhJDq4O8eSt
vWP80w4mXBFKYE7SFVaxKwZb9EooL4iHWiskn1jaFfyrZ4NCnGlVav4UJLe3VE4mksIITnouXmSE
x0350CJAkWfghwLWmpLS4Lm98IfKvVq5lJuuSQoavOL3v3B6f69vZqx7n1BCYFZuyBHa5TFUWmdC
4CVWxS/e/ot5KyIod1h60xy4f4iFVRhHenLl6fXRS90v9TI7vdbZDOziDtU2gfwTg7WvosPa/dnl
Pgm+M6aOKopqHoxbypUEfEUTEzdfOB5xBmkDTQ8cjDb6q8KzU1tjnxXLbp3nBE7OP9XbtybKd0PM
x+TPVnSPgvmoTWOpQWxnpolIcWH1gE2bVk9T7QmiyxQojgBjSuAesem1cqnNtNqR2yrEtjBnx+Sn
O7bpG/J/BYXCe9dS4sFWLYWnDdsKw8i52xIFSO4TZ6JeQUA9nzbOW3OkzxP3vH8ebM+bniOf+H5k
Upbzz07yIxTCJ8dSODvMUac6rdoOG0PA9U4TC08qd6dntf8lr5GY/qahdPwVq3qtVFqbZ4U7diTp
8I048N2+s4S+rgwqgCjgXY06svu+Ewasn+Q/FTMpUOuHE9hrX7t10lIUVTqc4b8W4kJ76nGlNf/1
AhHgjgzgnA0mhd+xH+VOdtgQRPwuZgusN67B7JQTvtkjsUDhuDlYNT2hiw4+EYM23hUVrpnzdaRj
LVs2rjaz9eIbaR2gZ82oGllTAl1FHgXlTdl1w3DJTtnEGymiIzVrq3nesesm3ztBVvzo/hWWP4zf
3owXOOfB/nybRbZYj++AD4z+78bznHXrGbLnyRUjVAeQpgAdA5eK4WN9vd4lblw5AWwfinAalbg0
7dhMtK/1VfrVK1qu/1TieHMaK6iYm334BaSeR0tmfNr4TDppazKp8GbWzVCPu55EJlfioDOvwgoH
53+hLBbhdSVr+5P+wx2FPctXzmHgPzK4iXLRaTZC5FxVeJZELLSQ3+NzOu3McnEJOQVE9kWjutrh
kzeNZblIi4Qg9VJwI0CzrZR4daQJDIBsvcGbQ850AjK+L44pg3SL6AZTbCN0ZWQclV3si7NcJnCT
9Mz1FKtEIHyI2UCDd9qS2K+4oWy4HXKug6z8WNjezKHJagN+3MnmCh/6o1WUgEhOwOEic7mZB8r+
WNBMETvUEJ2aMrnVJbReuuPZxDz0JbP5slqsUOlc6Sb+YmvXLks3HO5oLTUyws0P+QuXbeaLJ/cA
AhjPTuwYAiNSpucmI8GpTB40r6ZjAdHXplV46S4NUeUVUrPErRS+/2M1yQdNGUvj0ABY9r0cE1Jh
z/2fz3DDPTCE3CbjOcZn7+IMEnORCbMfYE0herELFk9+jUhQjjlnhIj8f6wuATqRNP8Df9enA2SR
SmGLaSz+DEI/YMx7QWL9e5kO1kt5fVMMf2hbLFbJil2KtS2xByzWhdimeC6Yp10wAKw8F3lhODWE
o+Ij8nv0XhF7Ehxm2fUScvSPpAPS9iso6BfZe3oX6q+8dHZ3fJC+7h7ZsI+MKYjOtVvNVtt+y1ui
gG3b6N5CYsU5Nu+rg/bHzRdD2yorjDGO4aK6kXk+OdSmcDaRl1+LHkZp4DcEMf3rIHNwU6xg9ss4
aCGW+P3wIkb3mLg48BizCljZu30xtbguQL/m7c5jkbWJ/2AhNn8Gxvw56pbJQ5rUgJw7G6TlGtpD
bdhcSIr4AetSwY7WHHml/J+Qcp5DfkqjS/VzrbWzDcMZxTiRRytFVmdZuo+1J8z5dIazbhnZ75jy
pMcy4gDD4l91FVwOeAUptFaerofxARG5InX3IXOlhhxpkA72PiSszv/L+gCtW5RfGCgSEbqhlUMn
Q23BBqM3OJZZTleinkSCurG9yoVKZ22bPEiMXaFwZ0gDNNzSQGR6ZWn5g5cmgxWgZCE5sfw8p0cW
fKaXR/a/g4+ha23Jiekn5oNcDZc3D7r7LwCmWxZLzgGJZ+6WqZOETVTPtCtPOe0RiAbNqEvHcUCi
WBAu41BBrZ0Fuj5PKJ/YlZsUJC89cXng2VmCdd/7swtOZRnl15vjDrph+dxWnHF65fpw2lZ4PGrQ
PT7wDNZ57ksv2c+9DirgR/+Gu5LY8+/0NrWqlc9JSVgDsJ0HLT5kQ80I0X0/5Zf9fAgfuvrz2APw
Cgc+NiLJ/RWUE735JCUKw4DGZjbLiIG1Hmdw6WK49PLSrE5dUwWps9zRisEropBtPJnejGSL9+UH
zBbRRdKHR6trmsZ8fiErIVLWWqdtw7FVNv2TLrFhdce3eEL3F6yKVhT9A1i0OoDV0KibqqYnlr2E
Z4jnY7qpvYbBpsWQj6iLsuPdcM17NnvWRMBnkFm2Z+d5A1n8iu3HSz7cA5wvi01a5EHN8ermqOu4
A0RwsWUSniNjzt5qmxj9N4oMKDnjhEJYDLEr9V9fGMMOxw4jY6D8n6+CGpKxcfrPsyjXUTzIlGpe
qdjMKxr8Vd4p2YLh/ED2BoKFK+8hSk1Mb/z3oCMY8oNFy6/uP4gLBzLVg/N9F1G2xsXK34rhf5Lk
48W7OsG2xcmqiNY/Gdpbe6s5tWYyig5nUMOxxTuZhQDJAAr6DyIO1l5JiMUuTn9yExp1vWTBV86p
h6wYep6HdApxkjWIh14LoRp6Fn/yGUKhDY6DZ3MG1TtZ6OUjp8KdsIiEmUL9VseLfGIvHF5aRYVm
loq7eskY0IQqOpvkNOoIlgHTx2S/bK+0wzmTbnI7V3iXNCsop2/CX8wvP3y1f3Ih2z/gWmnwCdfR
+KP7hS7rpyvFaZ1aG33YN/oTW7ZDSu8dcuw1yVAi56rjshz8TimeTRT/yBZUbXdzGEGkNdTrKMcI
izVLwXwbY4MW+8eVNGm9kqmrq8GCspkD2jNa8IFx6qwrs6OSr9rKI8Cffl+K6+qLS7clbbuwKZIj
J7KW6wEjvbL1u+jn2WI6CvonRZBCIRwkRj21784O5mHFHyeiGeh09b7F3mUAig0Gt4ZaTjnfqGW+
B2cO7nskAjahuvo9tiiDTMyGp+7lIBjpNc/RMTSgePf6idAZyz6bN+km9H/yDpK31Sq/BgcVQtxb
/R4Gr1nU/MhKqEfM+un56yd/qseCSjHeKeUicT/mE7Rxy7mMy7wyIYHDFSvf3GUCOY/HYinnyuTl
fyaUoZgen5586HG9QhXZgEuQgtBi6KoTHz9CYI/FsCrmGnIokASO7G9CkWprHESGxdBt6xjsYOcS
MMo5dW+F1um4Rp3GVVF0i/lZq8IfUDwnEx1H+RO9lomlWuudT/GYsyPpZwNfKKQKqR0R+4o7+g39
O2Hd2v/dbdk6+O5s7pZApGEoRGX3pfTWNRw+qB0+bcNtfH1Rl6pjcAaQg07doCzSoIdKUkniawNT
vKBql38XpJV4/AxyStQAZHhgrvoKMqQgd/7NV1DtuTjon5hnho1XeJz7LzEwlm+iX0bnzxa0bL11
ba7ew1I7slQkx0HE+3zXQ0CKU8r5xFp56qgqUX5VCEaR5z/NCl+7W+YnyLSOSjx8dKaASmEkExS+
uSd7RJ9eNg/gaZdmzP9zEHizfapMmzUvaRzBD6rKTeN9XjKey9r2yLVS1WqRj5GUp2K7iCvKUP57
HxXTlmgXczJaCSmP6T7jy8hdvYq4Hb6sVL+thTp/DmrG3UMriBTpW0+P33jkX2qe8/iGifEITtAQ
+ewZTZqr8njB5f1yc9W13dL7SzkN2NzAMYBr6sOdqRLmZHEi0pPzk8bcqJwd2fgPquLuUdWYZJqD
uI3zMCW+cImnluwaHBbzYcc/L902vjNAklmNa0PKuoh9OeSA7eph5EXhMlSEBK2AzlZuIrWxqMV9
LflI8Mw62KH+cZ00xXwYDkNzqWNQu78ySbZlLuhzLeorKZ9WS+HOA5/Zx0wrzfaYNugSF4DW8z2Q
JCv+vFNyd8Or4B5uzg2HLgEfw5UQxu0Poir/tKtmNt6PYtnCr34yYhpvMG3hMg/ai95L5pdVQzGt
VeQdglcdxrHq8wurbjwX/RElKX6zBdQ/22Imgm/IlLXeyeKhgD8xgGGPfxqloeeuTEe8kERxHImQ
fmlpelwTTEr8Nxgp3tYH1t2fP/+SixLKXBFcPIlyBizGb+gc4VrUt4Oh7++gtfNT8igNXJElc5Oi
edldMRCEVszf6YBXr8/oFvG8CXN9ayua6GUhjjG5vyVTLhTvF4BB1lB59xfSbSA6eTCxPCkLsTsn
yox2ZosmXA+4scByI33B4VsyVSLI0yJznBemYF2atEvu2dpJL19Aac+vMgl7iXoOsMQjal09j76s
+/X37dpo2PjPi2MesJfQshTDnn6YDrx8JD7VLGpiNG+zZ3CldkYx/sJfE7+PJdDrkeaOwFohjpqo
YUiTJPQyoTeT1m6ONNFG1cldOI14puUNu1K3u7p7+s4NMBeAz5EF+WLfSm/lIPT2eDE5eZNyv5Ni
zKqp3xvzsBLf77E5NENFilDCFRAFg/HHrrwXjLIwntILF/xhPIjuNnIo7/Ldd8lE127vB20WgELB
/oxsenjmAXDZYJowYYD3Rg9K7jeuR1wU8WZO9liT3iLwy8BuVpXSp66NqAiPBPVUFzMNXdjdZwNK
Tvh77SVnaxTFdmM2IIGwS9McMoiGq0H0g8R/ebkGro9GMPEcByMnOU0RAi3E0rl+u13KlaPx6lW5
nEuDwFFpg/jdVyX3SqQyk6SMnSdJscYnt8BcA4hlzJV6pCWs6MeYXZifB0LQ8VI7KHzLZ4t8/LWU
2LAiUfFz1Do8pWv08ymwtB6Cud2qzMjnjmue95gXRLWejNYepK5xqeQRKToLsNwDdY8PhQnSBFYy
bgmMBd3FYZVjmEy5GseijGi4W74pNzsN5btlrntZWnPR/+Y/BLzvbYcwWgSfT32vp04FrzQf5XuV
h1rc0/GIZhHMw7h9UTpxmyC7KNXiqzHoc4q1riO9Ynkmwge207s4vvMZFO02j2iLeZ1qH41DmpIm
eQIeiWZazwHbIe7RU+7I8acyBJiFd31sREJm886caCcq6ACwaKX3fYECQEcY7WdHgI+Sc04W90Gd
izov07PgGBmt49eu9wQyPx5RwrCbXDrCkc4iawIebPv8e6TcXaARvUdN+PRbhBTCerIcHLYLWHj/
ATVB+GiLQoJqJcBNfJxWOny7yHLbd9YA1Csqfm067Un6/tdBLnVAGrb9oG4f5OAU9I8EibqaWK4t
mroNjc1iraYLad+dWJ4CU3WhNjeuerlkMeq5dG3pQi1KV41XgN8ji6VbjPFg15Pzrdie4mNyhWjy
VUa+DcVMs63lDRLX/AYoAT0BG/a9uluQoEzzED1vnwrNRlBjKuJ/Bk5Umke39LTDVzGtlA0N8KrE
x/3ySFNcuxUwNL6wfQEvylL1Di0B/dmHxJ/LVfjD+pKMifp60bPxkr/ctyFr0+WjMgobrDr5e/WE
jU/2+7F3ev2jpeUsZaFQ3HaQFMw+Y7ZSfpTcLZH+le45kqpPvBnn//0kckVMySBktsCs8hWA+JKU
PXdIWt9LA2tgzWimllL2zvN0soPRm2iMhsgOiPPE/5jhPChabiIxatvfbfT222EnMjIicix3ARDR
7HeBgllZxrEtCqTOksSnL7aantIQ6YKc/Wp6o+BljlsSmLIhKTps0b8pdk3du/I5qGWWQydRySeM
ljkUEmbKwbLdm3BiuMJuDeaNNXz4Vfe94DfgEVMKHsG5GEqUgvdL4uIeaj8EiKWIQcZv5+DloW/m
9qRAs1MV8p6Wjff2K0ascQQ1UQcQ4wF3UFUe/yOPjrOK3pkn+ti45hoJ5kRuLHfR6AKH29Qo5zm2
0gWAaV9cG86fj3G+523mOHosLoJbNF9niDR8iFiXvlWzg7RsX5GA1GztRv9CvxQVFr2FiPmP3nrx
jmzhe5mJz+a5x40csaNZt7+Aia/ClQgblMH13t8si/jN78SRaL54ZbltkX7kmyNqSRgRqQu/WdGb
HRCyxlNM7ytnxZkS+NLOq5JRUniUv77m3sJiYKmYAxQEV9A91OT1FF/v9HRc2D8EtSVz00C5lOkn
st6ndNDHECD8e/Vybd25WKzBezGxo2KoM2lrZiPl74yu8CZmF4AIZjrlPZcG7drM1lsvu6UFLYYE
EZyAGV4L5cW0bIZ73XxbxAOBTienJOYnLKsCFR2PWmcF5oRa5qBnM7ss6kUxJV8Qq8HkN+w7/EAz
HA6cGLSvoWMurDEQH9zKVlgmuJy4MSEf5+10rCEie8jNxi1dHLG70DPyky4Cp4ojMhbUg7cQnLkR
ex2g7M47j/4lOwZB7oFCo34HOg/a3nBA5WazvU6/f3R10viIgOJrkxnuvjDVNC5biOREnXAFBGVC
b+YdhXqLeBFeI3gi0peD+G7Q4cYGNoSaTLrnLIBGHp/g+jo1QJ6Ik/f5HSsVzaKqavd7KVr1aHPE
pBX7VKaQoKKBYijMmeLZkHgwnDClJsGH+VovJADQ/hTgvw/Cbi19D0DrJH3mSd2aMS+lvgICMJSX
/tTd4M5HeURo0ji9hEpqZdS2RwrYIAMSOkaw8SAohWZoHnD2MnngaJXCqcuymeZo96aSNA9sa+dX
HVNU4W2el3Etn07IcSZ00gBFAa7e+ChIQP/4GXMpvNe/EgCrwwujjvJg4eh724fc1d27uX9LgTv8
0pALX6Go5s9TvCndDfQ/+9OU2nbBFRT3Kp7MPVrKTFHauDlt8oyahum1YIPgDjgxbWRYRneJ1e/S
WltE3R6rXQ7W0ev8I++29lB+bcB/lqf6BJAcS59HZR4JkQ+4+VkhU+dDnTkfCr2zUYRyOJUqCx/V
AQ/jt4wEFOS2yL+cYKgzNxDHwQpol3S7CttFWu6PyIWpjT2TAR+qKk2EdBCFrDTrEj2EZaeRkmwF
zfKAMwWCcDiRivbppXAKVusDP8tsUTAZdaKBG2o8f8eIk5ms6+aGVSQKgsBxlOgF5c556gO5XjTE
2UgAmKU+2xV3QkZ5FG47jFWyvBRnMY+5sMOwI/d35PzO1k1cNHsBtX+3T8stUr/wkERBYsF3UITk
T7oQJ4+yM72uqAo+YdR6gIAB21FElViwX1/zEiryKd3fjKGIqpx/EI8Dj2YRMAWPJKMLKzK62i/N
Xd7kx8Fbsww2++GFP0OrZKyubgBbMfWlqk1TUw2VT2ZK0NqMraPkvRfOcmTKeAeiAd5/Se/AKWhn
7FG08WRoKzjW1x05C2sFbM8crYG1vaHxBxI7RXefYnbGtajCHQZ8gaaZ78cwfPXWsdzdZGhijrDU
UUmOZQEVRKqupdHwdCRPp2I2BFqPTo8vAdp0dyA3GFQ4Y0euOqTefj57Ef4ey6XYwXlWXnhbzCqg
M/niQj9hTEYOJY6346yG2uhCZA+/7YbQJxpf4ujPV79/X40lscLrEawEJgTW7E3AOqin+bAyPOhg
l3Oclqg0T4ii2GOBNQhiB1iD7WQnLdHbrvM/DdTiLcKM+2DT5q5f8LqGOnjVOCGtNoue9CPQLq0f
p7XjPSbyMJEjtSJHYkszRM3fJVCobfghECzO+L2SKTQ1eHHLNW7MLSJjWXzP/fdqpo47hqiwtY4Y
UB+S3RRfDPwKQ012Jn2HMgikDD2e1la2hORSOmny11CzNkrksA+5tukCYKaxaxXEcWMve/4dNLHO
Ju/eh65iuIX65YhoYl+bU+FdGAo+5zDUzWhRlwySZv5WRF2GLtznex/SSKiqtCsEyLO5n0+EV9zv
ZxJNzaAj1zQXk0hKdiQhcRTVhHQ2s2yQdK+vjoe1c6AmJ8kfaK+BtH2RGAK6sVtR0GmMK2R1/r/f
BEGsP1Y0SNcT0BIWoDqrjJpIXfV27VxFyQB4Xe+IesgtIJbD82Ro0S0ekBBd2JcKMW1h3xoOHNON
N+FMAA0pHWPsC6BFfJg0Vui1tDv3tDJ4xzBvGEb0AXgLKq/nHso6dYjo/G4Gyd0LG+Tdlo4JI/ba
Z4sPnz59Nwwum5OzC8byI6OQwU52jlowChPmW3HuqRK01RqRwDVqhRV/2tooD+CJD7tkdPDqpxcb
djrh5syxQV4rpoCO8UAyHPIc8ft/qg+NAFehbgeSClhQH2H0jdXuDg3zP+QCdq/lMfbS30uCPy1G
3FZ3Q4/QTl8Muf7tcE3XdiNuOUJERbRFsi6U+ivlw26iZgvMUiHjg82c10tf3/lgZ856aPrjeu4T
Ex1YKkylX6U18r0rfqs23NfpNIA0PLH0xRU/0qRGlZ4Pyklw2EfyeOUJbdihnLOFZRzGrfZTvLA3
GuA10BmkfeKPfTE/5Esgqk948yUckl1IcSDEAXUnQcJplKutt+bL0c2sUx42luXiPyeWXRz0qSMI
efmqDMm2QZJzpVB/SXDuTdybHH6jjSff56YotX3WlUC3KfYgdpfWwLoG/sOEcKVnuX5Im9q/DmjS
tvOfW/fuQ1l3oAkPH8lacUNajd4m/GX/MjGHDqOFq8vxHhL5YLqLgi26VG9+cVuGAQMTM8s71XV9
l5fV/YgQhuNTbozVu9VFwvX+Wqt6KODLKcRGkoa6eU4mmdB29dA6Xuln7CJqpIaeF3ya9bHG4mQU
wZTz2ubrOi7QuqyTNrdQEZhE4djEvnN+28PAyZnJX6m5CjgcLcrmZ5gLCD38MOYZe5F/4JGvF5Q/
iesZ1Vxmp6TfAkr3Qu3c1mOSK/IEqwLVhlTxNGzKBegX5MGq6SL5uYTPeRYcTNX7Xflq8pLOxjTe
8rAlI3A2jAQARxgPkHY6lndouUY4xbz1/IhfsA+D0EtP1t0COGmIdxbyxuapvOwl8uZJvM8zZcPQ
UJm+vZLgM/1K/3xvmmD4f9KUtG2yYNUhKqQuVYe3paHW0itluCcnKNCaRSNbwTGEMHWOtRYrmC2E
EhFrlaGN9q0nE5bmWP0RzYg6eyfzBvazrOusG/Vv3fjmbn4aZoUaqvCgu50+IwHfnJIzAVo/b9qb
1juwO/125Wpxn6iOL3Vsa7cZes7ed9j9fBSlO7TgG+8a4Er3Bu8RssZjrfiVHOAkt9L1sNzdlrRK
pXSdcsjSTJIWGwcPYrmZh9XzrPm51y62ymfHUzgCBKJ+BNiwjyyEt7ww9E4GT64KfZ+QX+flQgjn
sWv1vWd52V7pe31hUet/XVY82bZFL+wAJoCx/gqGV9YqsLTjTqvohL6mjshvS9ZUvkzi3LZych71
BDPagWgMj2lUa4YvNcr6teY8EpvpBsFDSM85jfydPBeIlmIYaUllR2WTNcFM5x+Fy4aWbSjOEsL8
TcaOv3I+/27uKr+JsBPp5ZmSasNW698N/KO56RzysOPNUFpSGGxRg725V3FDBxaJKZ/oetwR0OoZ
a55HX4ibt6/2r0ZRc+yfmgX55ZQ6zrpu93AVgd3vhfQfIGXGBEmSGRu1l8Nnr0bhCJZjj9knhjA0
ZH4fUuEnXjxikkQXI2nzDdvATGf4usXwjzqJui6zhb6CVOMiAllGedQv8RqCC2xM2b5lTAvwO5Fx
HPymXNXpcdnF6B20157CR7pMwDYbYkBVvebNO0O5e34mP0fCHt4uJwT8RaP46JdHf1hTbkFYjAFq
zcoiwBEi0o1oZ0B07SWv1V0+Bk0QCJdYRAvY+/tqB2BrcXOcZQ7HJ7DmwwiikAvY6qRTcyT5pgYq
Cmi+0sc2abYOFJB0us5O0h89HSfTii0V2o+Fo+I+EAiX5CNuiZiExsNK7y3efOJCO4NFIRwy+Sua
Yie2L2Ox7woDmHGG32BjeBjRnLMo8RmRUj8FgLbLzC+Mzd2Kalua5c5V2+8qCUGfmrgVhusW9IjA
N4fHq11NINZz0djYaRevSqJQMoAow9J64IQcz1Zw188geMNdjSuCIvrBTaJbCrdlxVeg6bxaUIKZ
Sw4nrAFmLZYouPaIQrjFL5ba4AyhI34VjhIW5UFuIG8QoRLHHsVkcH2tv53F1s4EG5IJS1L1R8RL
Zb2pzwNBAPhbbK18LaFTcOpSGf0lVrj57Jvtngz1FQ3cAtxugze+6XQ2HVv6kwS2oF1xKhcoXhx3
mXsKpkfLYHrM+sg5/xSCUXMk3TGkRxLLbszJh7q0EEWTyycRjd2kUrhmbMeAoMEBLzpEhLAG5sXh
KYuRWcBa6aJh6PW85O//y0oWkZOXS8qxuplcoYzLLmhuOdy149v/nsWU65wMAaGiejYkP5KB6KPJ
1L6vsAXerdQ6AAzopBVPeLqpA/IxDiPQKJkiL02XCYMABUJSbfVxg7bp3nYkJr23Lsnw0Bw5Dc0N
5TLSg1yw0rL0RSr7ocAjvEQQlKdUufaGqaJmH6SY5bPhWAV4wmruJ1QRF6xvVsfqdhvKck1u0B4a
LoVER1xCZyYUeihPU3uza9HrRVhrCEo8z522LbAy+pRy+L9AlRzKTO5eQzYn46wu6h6kvHTtE9cC
gpgXDy5viEUq0Fz1UypzZcLTBemWnNx+wyHPOa2PL2DXCNAELiFIE/N20bx8JzsLd5ZG2VYlhHNw
V2cfMf1EJo+LO1oQZeJ7kdqWyOksKQIBT0ZSES69nRlPCBE0eXqNn0l6Ng4Bf11tOpvJlnlJUfWF
rURBlkYobnQyZoi9lAhkKJ1JFUnBLdlVn31cAAD2/pdgYA6J5ooc065IwMLDpJhf4qYQZbVdV+K7
GupbA9tR0sV3YcLFKaubC3QoIqDIdZqOBmnRG+2hNqsnRJ7WJiKRYNRCd2ivTYW/SD/5wdBuziAG
NQJXBufpQJJqxtZhjjHrDlOM6I8s48oWWdgj4Pp24po2uGl907Ms4WsSpVZEaWxeOA9jVVKK/l8N
YKzMhiAFPqwpILaOsk5xotOdF+U1tfayZWyUd50rpIBusvOk9F689j1Ssah31a7VjZEJpqixphxk
fLrv/UO/77sqwnHWdzb/CDIyPWsai9x7DUmlO+Bpe6lixuW9Q44f1nnyo+3W0adradmJ0PJDpj98
ih8h0eGAXvu9dJHH8jX+FlIzP6ZKad9nFXL9Ygn+ekYKgudoHm1j0tB9BV3K+H/3ghxgElNWKlEK
ZUGakJ09qbWquMU6uUUb8CyofX0zRgRAkziVycJG2TeACed5ga+94cRnQKgVHF43KDg4sKXFh8Qg
w9EwHQ0jg30ONU5fdRitxoL1TtswKfPhqPuRpgPbKvL2P+p0xyUnD8mj3UCWLbvAcI+sx7kD5l4S
7UhUT8wzIDj7yhcVDpNNUOVHzeHYs2h72Ak4Q8q+WtApS0AQXJExoRmWcG39Hr/E03o6dMwFla/O
oSc8ARRVzR3p2So+MGvm9lUi7hEStGgQjIic1uJYZsZwAyyoQ+0rgqBH4YdXK7Wh5xT1DJA1nflc
b5LXPyr14Yu0NSRnEG8dizv3D5h2aCG7toKu9wVeuR7IWh/bXwJKywHYdCa9pk1fgNRsOouvw/fK
1NeCs48unRjR9rEp4oA7b6t9K+RU9DRjdbp8FZh3NkVjKUvpLkCVCu3wVdkpfl9ZHez/k5Jc7wGP
L1Mtiz8/pwBrmvIUgZj3vLpmyCG4RMFxarVVoLCvH/LyTjX+I56DReHEvUynkkSCCzjJgUHBjzH2
okk8PcK8E0oE8Ua+FiiiJEca3od1jz2fvvVV5fjW8qj4Iuga+ZxJKax1BiLQ1Km04I8FOPeCMNXs
J5jSZ5ybr79g0f/gx9xlHoblEZ8iEdLLpDGHK/CHltvNgLU7SeIakm9eU5iKobzPVK6GbNfQ03I6
YQcwPmqR1eo5vSPsE5vrd2zqLu3PkJT7Bh6NTgjxpNPyg10xDFVIY6UZT7KlMGbzu8pM3draGmzs
FnUqebSk5EJCnMpgisiPDJd5GmjVu/r+16psZxkzsr9na30hREoAb3o4HniUfxqXXVdax7wsB4wT
WEjq3XOkRS243ejdkLSvxweny/rIU3vDxGuuaXBjBL1GlLbU9on1C/62GCQt58MMYYXia1WwXXni
9Mgm3eVmR/7Jx9/vDIXqYKpyUP8YZjfqlLmd21/k6z6YTlQh8cWUkJc0tl/o6lu/fjhuUnUoIfCR
VBgwSQXgzlC/GsROIWofbULLH8dkAPtSShDNKDlp6w6A1dN8tYPcw6I6mNqZhizrZeKl/OuV1tid
/PcsAwh4DRumJNkDPcVqgjxUBbBretA70D98VuFWO43/CfXhabfVZKEfHYTRh3PmlHvJWsq+BnYl
Me6B4ZYgsYJxQrC8734y8aCAxI7PtPFssLK2f8RjNP/ljw4ytIJDq+4VOcHBL0OA+6YQECJ97dH6
oq3ew5+bOtPbLfUePR1JGMjgKpxofoNxupfNA0m3ZvcKecUXLJGNqSufMdnsChsWk/i5FSOLiVbb
AOOL6/d9trLs6q5DQU9+vOB+2letZnsx41N02Eg50ZiC4xrgsd1dXafmwHb18xSxjuaXM+7OHbtT
9No7N+/M9SDvbjN2PtTRviE6e08nOWaZTGcGll800E3ABO14YOkQ2pATWmHAOWKFn1uzrcexRkPq
1cvZP/IvXjyWuNT6AIF05SFi5D0EHGi+sp+oIC2x0hCOweSum991spwq5/4ZXw8AdpPDbfqC5ykY
VoSwLnUxoBfwg9XXULUW4WjrIRRVBJQqkrcOAWjIhbIhPg2Vty9+sBmOrjTwj0/gj+zokd9ENzLv
TBdizIMWivWDQDmym+i4Ld/sKUjn2qbjZ+DLfHezOSYb9Fzmofgew4me0SG15O+63LRtknYTCL6j
Tu+NkoC6AUUt7ZvMSyvYEMQebFtlxXCvEEoz9NrOMurIPMK/LOeHlpuxdP9qStn9BKnEXYtaLN3Q
zGp6PdKKMHQKatWq7hhQonToZDhdwBBhAxTIWPXu8WiafRbvMhU8CmEy1cC9g/QyPNC/eEXXlvd+
tKDb5IKtcWYD3nDXGobYBZb89sCzhK2qPlc+7fbz6FxRpfy17gBi8ImiAEbpGJ45rwfdD9ljzEtH
AXfbQnnrGAipS9XJuvHog++bNyw7fZlx8J/Soukt+GXRzB8nwxRtBI/fgV3E61UjccW4DtgRDBa2
BmwoQYGs8ftRUXWYw4y7C/w/A/8lCz8Go8AL8TvjRZiuDZGg3hFfVb2LHXxKUsaEStj6PBGj84Q5
I5VioxJJNgxabxTgQllEhsKhx++mnKVphKEZH16Ar+bcasrOsw3So77EUs/U5jQgNdJGhNaUUbqI
waFgLdKjBpMvlQ9f2M8M+RBjDg8nrnb64NhU494YeA+TsZPJakC3JSr+GP4rC5uiqQ+DVRECNBf3
0jWpfofn/PrzTCWg/lkttU6v5NQctvb1tDm/b2zAecs1mtEmcAHJ0/1hxviOvm+BVODZr8YToxDT
VFcwFi6hkEKNKh3PpNLGkC0q8AZWFiqp1RCeo9ABWiI8Z5ScUuLF5tg/6H7s1ZA7gRjN5eHhycjS
+TVv1Luy1d6JSB4W0ifqWvimy0/dvpOy6+4/vqpcQTchYzqHwybg2B2dxSmaIAb6F3//VSpHEJQ6
ulpjONABhzAqZihIv7tAQD+LWOMM1YfEYNdPEKfxZmBQjME52qvxVN0Cp5hgYl+pSS9sBvqYsJfU
zpCYe2ov/cgVJ0yfODrhUT4g9SnrD4koUvs6W96U4B0T9cZrBiTNJE4/2M17k5s0uFm9jMSD+ETA
wcBhAn78Fl7FjSnv7W+VlU1nNpNfmAi6CZ5y+RiM0hY7O1CzAnVa4vuF5mF+lOLTngg6vZeZ7p4J
8QgrhAgU6E6lP2MRttsSddWKE2UgwTfENhh7wxbHHD2DnQBB8DaRfikY3g3h+WZbxGjvHM2OsH3p
XNqEs0Az2P8RUUTuXYQ0tPuIbokwGgW8H6yanw+Bj+6/xjznqRFHimlyAMNLM4Nknq66PO2eNirM
m5U+tpt5A62IIA1jY3Bl42zTmDGs2vTQ77cKkE3adi5AuCJwEeXjX/RZBNqLPQtbfyVPicrbZojC
ZuTYjuY6RsIivp5pRb6tzRGORv/aXew/Ot5FPey2Vcaxuol2TKueoWWfIW+nCtGaXKRB6Z93Uy8D
2kpZBO42VyKd/hiwz1XD/rZHfBA971tHzYC8vt2aH6q1ynqo3TecWHMKOALzuJhhvHE54O/nkVoV
WjEI21HQXT5mY9Z6cDgk4QRGTCfC1uDgScTsCuBCOTKgzvE4lJ5Inwwxkw2XXj85wmcTt6vNKa3Z
55Q3aZkh2p3MAEB3AuFPbZ8ri0W7rubB4rAuxeLIi34ft3AkDRf/gI+FUSx1HYpnyMmauL2kVeV9
M3IIYuemaBe3lW+x7vVCcQXE6yJI4c33ZLX5ZFaXYPo94gy+p3UHuYKuqYwMa208adl1gsKk94O9
xiiHAM8o6PJlXHS2nKL7rHO+6Tv8QUVgVOHJFktTBsWUdBhmmNvn6zUG2R1H9t98Cwtgtq06Hkvd
ELQXCn9Bu0yavko/UEq+H1+M9kzwQwy3JHn71aiHY+rPm94Apo/D9+wG7owfKaQsu/Y7Ya9giHLe
iD8brf9cl8x9biEidfS4pw3ASkawiz52JDUkSMkI0ynWQ362C+zrJpvHJr1tF4Az0AegwxJ2P042
alhQYXLhc7uYfEuN/8wDQhcUlqP+9Um8NqNdCTyCrf4a+9bITENPSGJnYcPjJk07JLllEGcSWf7T
9mioMjpIrZDVM611+/7lhoTQn9/OHSMaTozD5/b4awJB/YrmoGJO/NGo9OuaGitbjAYHfc24NHjL
KwHH4orNDdRpd+y5Xhg/M+VxExnjOJAEVFLjjkPbrc7u5EStEUw0TZzll6V0jGmExVHefYTFLdos
K13sftidyJJVTsiqeMqmltXvFT2B9X5ydd9ft7C3JM4RjSUWMrarza/pUIALxoIFGb5F/BfvuY0p
GvbSvjOjUMvJoLOFRlv2acKS5cKPfaQ7hUc/Imk2SsA3k6DyV5tCb3WvF/wAH4Faf7sO2GBkUI/c
Y5JgRpbS8kfWTglGgBTTSUqdLEPtiAIvmnKD6lMZ3nsy0ceODV/YyFEeSTF3h2F5W6XPGffjK/i+
9zT5kXD214l/M6TTOsFgFtU3QhYo43iRY1lKJg5t9v9tz5Cp6pbUHQiId5itlrg88X4Xf70dXri3
4hZxleECz3IFXhI/l+H/ma1CVY9pKjqs8idpLShxOEnooGTzZUHfiHNzBCvdnw+vA+NBrhH+e0sT
ESmaFpc0ZgUTJOWLBuywZsHLkTcOy3iVBgAnhbOpCYqoPj2PYyluY+Omn0GENBJU+1SzxOuFJIZP
xOjG/TUM/Biq17hfJVt9o1YSb2LhZk/3rOUQ4v/uDnd8LJ3rpSUXGgf6ovwdEaNhCz8IfIXUrr5f
lOIaK43zlG5w04S1EcXDP/4zJKRAotFqTba5LS9quIAbbcfIrSS+w+JRvG89o83Jr19p0hKD05ad
3Djz74MBDgf7N+vQZIehL59O5wt30m7nHv0v6rKGjDPkIkS45uC/yH0FsDdfhkdTl4bw94Egxpgh
fXCrnYYRQr/KhJH4EjZ/vE6zbzlQMwjoezJTBmtN7vPyze+UMocnCbHdboQT8Bw2slgBpaqKYseu
Ll04zERKkhJZ512EVl3VO4Nv9wqhu0r/kbdVhFBu9IRaHki9+7mDn/+7hO4q8p7132L3HH04tJrO
EIKQ02Lw+kEkI4xsTpFXTeDeKRK6U5hz5+goVufbPW2s/864TMstpgnFV1GjEeww76uIeRWvb59V
vuYC4vAq6dOxbJ4MjI6Fhi0iLseRkYgCho97YidI/7XUzvH8bghYeUErwF+DkTsDGl+agVJbItKc
K+AqsaIkMl8jBYO8Ead7b0Zd5LyqXBtaTFC7E+8EmNxnFIqSlbXRS35upQfRwuzdMBtTiXnxKyAn
9O8ixM4y8+33wKiQ1s1Qwy+5v0+bfAKGq4prUprh6uVQn1oAxIklQIHYiGh0fSh3//bVnBBsja+F
1EkmZSw8LqYhGSt3YF4LvOkbrxJfs51g97lJtP9BCGpRZ6kEViI6IQdaOQfmlFNlHoyvYZeo3FS6
Rl7wuYCQGQMpNqNDEfYVFwpFQCCNwamY92oxqLFprhjMPYtSY/CY47GB5642NQxOmt45idMk9VWM
prjxS9dTLnMCkEja3MNwF50lyV87rWHK/htcYbIYq5/1a/w3MkSUAk5BRdKio1Dqb+1ur733i6L9
CxYvBciJlqLvRcACBC3tKfj+1cqbFA6ftIhZ/Akx6vKELS/C38Os8OPlRWbDbDp7VPmg14z9GGCV
2+x7nlWxHZIN6ojTKNiFGbA1FSiMqsw7PVK3/Z+8b4S/G1ohFSq7ewL87ZXfIFwjQsdVMjuLaAwW
gWmuo8+We4cIC9ZXzdAu5nb8vdLyOwxCdvJMT8TzGKVhxJG9i3SRhelLO04ogLz1Kgs7rC4AaP5I
dzm3nJjZ7gQjgIPfWz7qvnwMOM2ZE8QSiLxrsjY2G8bO8damEWZZ+JSsg8mfYH/mJWc0oDSDbRLA
5LT2wuf9ditr5hdPlBAZt6TAlOkb31aaEgg6TMwGvqiIFf0r33tXOFiH46GGoOafRsHWPS7mz4Fm
yUBLedXTjHbSnBskCZ05owCzzC8Ctd3FO+1b/5M1cIctNinzfPDues4pwXalj1rv3I3SjrXreL2a
t53id/Oy5vxChQTxC18aXxeGiIbawgCe9jyzayGeQjHQOmiCeR4fzlSutBmVxqP/mA2GEhxmUZp6
RFGJCuns+Yg8I1c9Z9rmtuog6I5exAn0mEIzZ+naD2YFdzCEY82sID4E/LrDi5Xtx6g3q5Uzsk5P
3hyeTp3SnVcoGE3+kUiEKwIq4Fnz02uZUar1kifwdQzqk17xwrlUQ+oF61VQMIo/k/D8Ye/HcQIl
5Q89svAnUrei0YKK7ktoLidennpWr3KpJrGk3+DQw4qpaJ/A2PZfeL6z535TASYEeUYZzlqAnQrT
O8pHsGJ/Z4O96L10i+mn3vXM+Atb17Tsq57P56ygqln6vOc0/mFIkkeqCMEZGWCWWnSKhHRBEjNA
Fax1xM0suLppmuk3GMQJFjIvfQY8829CX2ZI45BuwRq1CVbHAbCR9G0ZgCdwOqR/KFpu+6OlAjpX
9IHMCe2SFEqC8R78Ce+CM71DiMJ/nuhdbsoQB3NUiudrJWbutIV+Ce/xybeVhaKeruVEsAuWr2a3
9Xjs9E+wJDJNcr5gJcyMDN615aCGOSq8FglfrhSKyuC2NDA4fWof4so6Y7+RY1IUmqgCQPmV6T5e
clxVeixvR4O0/ZABJMt9fL4cXfk/6KtcACmK5VWkeERYgeKMLjdBx2MW7+Z85tutKq+1usLccjtp
KvxT/hYqRu3dxV34wc+R8/+ksWKUbRKasUDqrfsy8U9TJxSYVTtjgu/hgauxTegWnBFqZwycgP6k
IzOIEyzKWI6HOQOk+J02rdh+Pi3fEG7PeXOJgVNMnhgN7LMOqCugwR5xelCth4Hac7GRJWuApN+/
DYV5YKhEnvjgHKvK/zoXTNQGiq7PbCMM/cC1XQ6t/0PZ17b28gMQg8wN6R4pW5rGPrx7rfMLTA5U
zp3yhrM+JK6XDaytgnlZgexBL3XPGyPaARvN7+ZM3w5UZp85cSCam02MzNkzHhmJPLdBGl92ttpy
5PMV3HyXOm/erD9KtFVZYCiYQQ960sg8II5du3ZtyDuwy4Uc9PcdGWYJcZEWOCLaadYW6Leo0qNp
Ap9KynhqLs5qtEhtlR6X0UfOXfdDO5tnbUEaNXcaV7IMo4/dsVcQcO4SJXSd+oTQvE5g5NG44oT+
bQwTPM/jo5zkhiw8BhHhRpSNxK46/Up/X2kN1og5+7kseG6RsOFLSCJdWSqXUay9KnKlyH0z5fWg
aqpI5/oj1TrsIAtrmfFpFNchbUHHN2E6ACZ8A9JRwvz3QTlrAkBBAMsH34fyCcEMI707XTRSuHl2
9XGSCtKdFVeAuHqzsTOjHDAR+7/FYLG54qILnjYM2LSsjHgNQcfDlHprFv9cq7c1UCYrtidSgss+
DGB3N+cd0D/qHsbY1mOJ7/n1CaWynxW7qolIhWfpora1hMleRLt0jKSs3+7edKlJBAnksDwPXK2t
YolFzU55JYCPj+QMRhykDDCzNo5P62n2nOVaji7X7pVIeINz4jrY7Rl33x98pvJ013/lMhbFZ4kx
TxZr2mfWDtGiPB+ncgdpOtrp0uZOnIvs1zlWv4YA5Cwaz//WueG4d1lqMek7S3l+LGH4V8lxwA06
ziI3r//SWCSFpyT5b6HDGNjrEFGUj89RWbzgKHf3taYwMRcBYVxMK9VPHsoAR2zG2mO60U9Fl2Q0
acLi9WotlAjHG4LxDkoLqfjXnzLsIHNDNkHnikvk2tPA2Y79gMgyoVXiXXEcsEKnrizECI+T2sYw
aiMo+KbE+ticpl3H1BcBmDpsavx71QdmYkEaEpRR3uJudW8PuduWmmTqA7uFBSgxuExXpky5Ji8P
TL+tx4it/Bm87rrqpAT3PJjo6OPGEgctymMIAHOjBMqSyeB0P37qQQD1eZUQvs4Nv9ClnwuHt55/
rCz2AFi7+idgt72STNpumo4qL+5FeyamzJLFZ0xQPrbQjhQ5gsEhw/m3nHNFUZ4tbtc4QxXmyR1k
bzRlh+6mQq8awd5Nonv/hljhJKyt8GM+bpw60iKcG46NWJJNmziDjJQExwYQp9Itj1OBDiCbKQnL
tCRYI5HfcDq6yI4r/FInbJ/qG+x3E8aOjPqAYGUktklreF4kGlOIJjtAvA9LEkGho3HDIysxrYaB
dCt3xWq6Y8yVMjPkMk595qPWrxIpYUZEq1EaZsE7Bzo5X9GkVxvRBOPUpdozlNee4fcq8M2DIFeY
WUGBuCt5IsT0MXaie7ITH0lph/PtPtL+lYzG736Z+mOJvuaAiiYWkMeHQNQga8UX1F0fxzx02gUB
B9/vhavaVzQADhol6sNmmL7vFuwNTjka35bVfE1QOLRggLtfesvsq1OZyRgEnAEDelSiRza8WO40
KFF6yHjOb7sQlztHZ32YJ5gI6VdDMWY/IFSy3uYJU47LA2RluSN+IywBxX2le8IA/JpO3lgUmxcX
s34r2B63Q46veLnJDFMQqGUdTnW3ZiA7P+M6ZK/y9BfM+LkCM81DO7dH8rcLpVaAffZONr557WUM
ylLxtE7UzmmgLS/9Q63j42mF6m9Xy6N8AkMAu0UqocgxNp8WNGG5B3avZqNvuJpjgSH1n1Pc5aIY
7LbYBI9P1fd/p0Smc1081AympuGRKpNkm/xHxFQ9F6/W0IU2CzlN6aeoLk6oWqv0GsMS1EGCDdwC
Yb8b2C7r/k1jPcdM6GJCU+0nsp0QXnV+BoDwURZ/ug2+vuynT+UzXiHJjJWZJi7gcXcNFVHIbOaj
1N0v+ISyryFNcpRA3XCWaVZd8pvYWocUWGRP8AbifOPQHVp+sIO1aIrMuPftjBcRvROZNjcayJBS
EAWFl1JvvOMvmTSqcfojjaGLeQN36kBuWxJ6QM15p4lBMfJozRlaCrxE4wzg9DT/eoMwRYpJYY5Y
SuiYIMfC1Aa3ZiB8Nk03/Gr9CbbTDgvaVGS8SwER7PNmZpaOvfD5Qe13UrvNj5BEMWK2Ih7l630v
4hWkEEuhDOKVa2afUVw7QWDLTuN1n5tLgBhsX/CfEbjixM2xNC8rtXyL/Ay0IWKkPrWWx6wYXt0+
IwMqay1hvNPJEGYNdB6gcIYLNYN87P0TBRlMr1cH3CFHJ5p/eN21r+hQu3RdL3d9sDFAm1diQ3KL
lo3hoYiF7IYGCe/jARDIpPZPpAdsNfcjng0bl5QrsSZFee3xX4keJFrK/GC44b3L92Yn4qpF4o/N
2aSi8fqdDIMtRAvIIc9qDCSCbUqq4Y+FLeadbvshwSRYaQZeYeWxgBbqMFYerMZ5UL9HLm/nBRMD
WMbeoCjJgZZEB625xD4bRNyfgLM/6YXE7dyeuv/8+Y4dKtu9Py/6jpNs3JPFb9e24RbD6+nC/bCL
cwo4hAiqrws1mFUX28Pdo2FKPKDiwS93TfUl5ewrtH//4W4wtE3k++gzvmH7s/Iw8MLqk6/0Zrzl
YlDwOry5hVjTuRKO9hqmVKrrOs0LgiwViaZAgIPV33zszm8/QmJ/JFsSLlNKS9Zm7e/WN3K7GMkX
HA8YE+UqXvDr+GZbnIPLxc8RiUzufuC2JZb7v6ViHs4t36LDU7i+Itpzza2XuG+z1A6ID6epfLI9
O1pnvKMksAMLUul/MC5UePtD60fERqtsGEUXcqtHvMLHytKN4iZiQc22bwqNfblBZzuqSl+hJfsi
ng5VHLbqhds1gwtuvRc3qvLPUjlU/Xo86kEjYDEBoVK9DjWMcvSrmnENtaUp+Q793GZ8sbVeGaRo
1tQUTuJGhqZIZlNg3IBf2eOw25s7BTPju5NUGzFukUXVh+MkH2+oG9A08C0ma/YLs4J/7B7Wj+3K
0jn6Wt3xb1JQUhIcQ2qRav4u7deuvkHx7EqwVcpjNGAM1uqzyFU15tdsV5LqinyBkyRsZHGAOJhX
M31nN+DC1okUpVYV+dWfulps9SkZn+N16/6Znd/jboO+d0NMqmIjasjfvRQg8CjpvHjdp5IPgh/r
VPr58uZ01LCrcXpvGVyiNjy6CyeOgwOQqoO6EXcoCDHtIPmAnY2sli1WcAFW7Cgt+fZnyLU+amgV
pnUOTeah7wmckSWjbKGPFv7DkrIJL7+zTWxMccEXYQAzX6pvaafCJ0IvjTevIRaM6YNSIFCaxtLp
k7wqUyVuMbrVSZgLLybnQBRmwjGlmW5pdmfPdT0edBzaVbo40EQyZjMs63WbNlRfubEM2/aMDU4Z
I08Sr4JPUxUIspShbSb/1v6rHs500IuTbdk8rdQYuJ52PpoeAM/PcS/FL78ueAjXF9dR8has7F4d
npHUVXLuSu5TnJi0UKCr/JVjgTN1i35u4TzJZvmhmAF/td58HOIpPK/SfuL5i7xB9/pm1GrJXJWX
zNWmitbH/XI9gdCDVAfyyPm/oRKgzl2xKkfX1hV47VpUYPZ0vG5gjJqdxEIVXkgucCWeNRM1yfND
WpfOg6azZPsrm8ie5x+XFKTJ+nZ1Z9IYdDyRPfVYKH2J5z12lkKrDIgpoJ15783lbbZYXXoPq8av
P2+8uFoR+ocnAMyf21zA4ar9XlNINokVjGCH4eC/Ul4Ge3fuvUW9m2ZVzkwhSEN7Pe8RKhusndPh
E62lAV54auTnaubdmp1/q9qV/gCqwRdbhj0x1kCIV/IUeGkrB8ptbx42OjHwz9Q+s+f7IycnzSpY
kJrIMMb5XzTJYl+5K2tUTjeL5CMwAIjqrnRVA9YTyr+RDchxIpk6kr7tFiot3QIReCdPa3FIjTz+
qqqT/km5rCNyNN+A3lZC6x0vV0JsSpFs79F01osqOa66QNyW0nRGNVu09ziSk0qu49LiCAvE+H5S
TWLcSjbLv6DqR7lu53WIY18j0Nm4wgVAg1EL/+IiC11DB99AqRZRYUzTzPPQj2ZDXHkVUdCyQLpK
LPXdTGqccI6J85+xSuiBtSz3hxMZdqxNgRWW7FFvVbl9gLedYvZ37f+CIhJyxEy5lgq242vLyDbI
kApjMpMo835shTqYzXREsGSYO6ZuWCxl1IuEXzg9FqlPwFOhKbZII7bBYH2STD96Zn19ku7jiLca
x8x1mbIA3Uxh5ubFD5J6urwW2he7+1qiuS7dBqdtFAJE7DPCqNAkSVGJftpnztDSA5D1Az66Mp1c
//cBtLtp2MPe3aBR1Ip1USxjG5oX9RBDE9xmlO67H907yzr7Kcy8VTRcwr76tz8gARQ8T8sHBZCa
HKS0wx3zV6w4fBS4X5kMAzbLF0o1L8JbTMBHl7HZFTc9dgufK6clDmczznMtLMMnRmDEpFLC1CNm
byXj/RQ+59hJtpdwz62f99jSts3ARPyyKEBjTkkoNu80/cEcTqRyqIqNO2ctHXmLTAMQN3ogxOkl
GQKsjFrItkfHnt+JOJGZ4t5eDJUfoMcZyGMvxfzuUWCWAiEdVYsZ5W32HdhO2kBwKim/8fRw4tPz
yACAQ730yqVQt9UEF77pk05cR2SjffMVcjigivP5YZ/LKkgdILwcgufiEWYPMQ9sjy7oLt2oKyfh
NMVC+JgX26/55EMc7bBC1iQ90dNZ6xQmZMiJoSwBTK769vPDHrD6UtPQAkz03NOB/cNhvGBiozA8
CSs0ymhPyWIhWg8Z7AhkI2mOiaus8E3CXzbTXQiQE8UFXjh1FUYwD4OCwPrjUO46nm0TmzLf2Wcm
OA4/vKYlhL9tFI8rRzJGVDRKg4zqUcxTQlB85noxy0hZqlOynhfZxf0X3lzo3bDM14qWHE8X6qD1
ZBLNV006Uh+wzDaYxiZmfogETL4UudSAVxM4ovmyg0+acnVgefvWD9U2p+UOKCC18gRQAYzE0PQr
tcDSovKrJM6pYvV/wEuQDi7e060/D3FtDmoFKYsBL58AmcK0MKqcWf5dw0OsxW2oV2kSxLw40pU2
y4iIlMkDI4FAGaOxkejQxYFh2tkDMAygBGhNcxV/8RjIHqgJjU9ZkLYcZLAbYw+bH2CZBVJRjM6o
FXG/WJoPzOHFX31RdiLJKKaNt9RJad8m8OaUS90M29BEBkLPuLtHPVro6zA1yoDxH5LTaO4RMf0P
hLFKq3QzPQ7YO+pfzayKQnPS9ilyp3F0qNf2a7vWNKFn1dyrNZjYk0vLgRlLKKPsrhrB2ozIHlLr
MYQf6LW9S5ADZJflfLw892ZZJdHhQRpYFFnU2ygGNsfYi0PsTTkm1ehMYmNGA+TLpPJ+AfktmpfV
f1PvU6GBIZAyZLtNcCNjIIxjGV/GLNqH6I1EXfHWJhmpJyQ7pdOVUaND/4UwXZKS8RfU/7H6zsld
79ZWdEpQuzTRDKW7foZhKywgajJdIMNRB8tSSqvSpb1R8TbEo/p8YQrHxVhGQJdNarOcVD1YuxHF
IUiIp/puKORiLjiBtHNX6WR4tRHVLK5wHtz6VwBIt4pn6e+BonmTQJq1ISZjGJAdBJ7sSVfyubyD
U2iwlmKLRKTPLU16gaMmjtCj/GvmG0wNWIzcLMt+v1dE8vEW4ocn2pw0VYrz2YJMJuHNki/RtjnJ
kzQG9AZY0lkbDKkwNeYC4AA/MdHcyH0P4xSuOX/4KUccfA3OO0IbF30Jaa7GyIq57c2gD19HX74S
lIeJzuNACNhQYKs/YwgxVLpSAW4rCLqnC0YB+1k9B3j4xPptdSK9kMob6VmLFt11G0fSYEPj+zbV
vZSMC7HZyFPyDUTHB4fOIwd6eZ4EQ6a/d2xTsZqSGcHaWsg4jV6dvfSpS9wPWHj5uHDAuSBqQNtN
DtvJTNXHRCu4PjbrvCJXbJ4aml6T6HKGnUCdOlZNZ1FUwOqeeu5Df5/eSSRq1wYHYryRzhlkr6yF
5Y/90luPpzIQfMbhY4oMuhabNtblrG5QResZVsTcC3/pPLBqMwreK+oUCSgKXlmO8hcTI7GQO5cX
B3f8j4ICOYQH00+ZWbqoegKB0HZ0XYEkSkXvhRRH2enzbzGJo/zGUgFFmWOFUStQ8rSLmX8jHUXf
IJgLJu4E3IGtpmzvFSev4F/FgEo+j+LucPB6fZHq6KcIYvbzYREZ9iqpXl5XjAJKSHWRb3CddbiJ
iYSIiGge1UqJcgkF05vdDcEKMGe3SM8l7FkhGxmhgQxmBm4xbIgg5oHN9fKzrtkLHbMFf379DQrH
srFYDqhGHYqBXwb/67jxcngYWuIW3Uy2U0lIz5Tnc412XqdmvjI4ymzuMo5auqpyjSVn0YhmjW6W
GXWxxYSKucHrLcFJP2ut/vObFcJXh4KjOqBA+wtZEBfJC1RW2QfhQddND8an+d01hvMbT99/CKTu
R65SYl4u5OlC4z9AxGG0TezJdJ4h5I6gnHNUCpjBxL0de2YgHOA3IdH42h9bjcopyA7C89292GY3
mYF9T6iH6Z5dL2mqzbb2mI7/e7FwFTp7C5cr/Jh6hfs4StrGf0TKWtVUmnSI6rGGKHRWuyhw7Z6j
QBA+7n9y4+9gIwE6Gg00KG/l6AVqBub4eiUdqv88CcTP5qcXkBUpXs6sdpNOlAgdYxmd8RCCT4GM
d1+dVSwsZZAJAiJzedLxxjmstQyQl5ugAg5tgaa/cCqzbdp1qnGVBNm7+kRx45B0IKow4k2OmS70
qfeJKCh4WVgly82PE4fFzGk5bns+g3uMub86g03BllvQu10g/vNBAyResctIzSA7RlLkkhQxPjID
i3sdVvv04qqhKCBmQElsKi76bccj3uFSXotRtt50z6m/IT9jjWzQmL+9nYMejRTpjVEwsM2LsXCP
pcR61lkXDhVWwrHW5zLo9wbF1B3lyd6U8M8rbKmhoIo4x6bfuQY5OEZhjh42q9qVnvJ1vV15+iOf
W4Z6r+nAa3+ySgThzO6nPeZ1kD7l1yUiLOIGYpKn1mfSjhsYFiO8fYENK3zsfnw/1pZ1f3cUveKM
agzpLmxSjNP7asac+AdpezVVJcCmym4JmrHphc/rz8GTzZh70HilTRGWCOOlu9PpOvxbLuJDtRw8
SEY1niW0DrmWkXxkSfzG14DIjeh1M9Ezzuo4JLg8+LigGZupXGxDOlmz+2Lv8DUShRKmQbQbBIxL
fmspqelCa2ufROGiBp3jIvJ91U1twqjmrpkVi3eDvhCKo/to+nCiS3NJZ/I6pV6aHytP0iYELzUC
wsXKyJrUvbxL61jfAAi7NYY7vwviE3NTxjhZzQGlK1Ksjk6XllIV+srf11eXGs0TOJEgsxHf4z/G
P6nUMwtOm7O5fNgVVddS6gpBRvEmS4sw41sjwS3JyxvN1Cwdwu2WMUVZ+GjzperENkHgwuV9dScW
Rp9yzgMoZiC1sWZLdaoEB/ejLqhekrlgW1FA2GwYwmNN0fzwKU4kBQHvQebYhlAmIZUqwDgKlQ8r
r94lAoENzsS8JAF6WlNTK+01mALWxzPN46aZumhZQ35f9ywiPDabwuL+GU2ND3m+d4gRlSyxH9pe
ePzW5xvW5AyQeJo2AjsAsvWdihauHJjunA0KZBOllWfeYZZ/Fr/cFsfojf0jf4k3UoXkM7O16faZ
XwSiOMlAvHeQCCs4ZtvFdtP787OnRgMlz5f3OtEwzgzlbDQgOP2uI/4KZTeO4ryCjjxmNDA5Jfbc
DU6oL67ymQjxLIKg5BsM4HVDIFc1uwVw7HKYKQZegvSdooTYC2jrZUK0tpEchrkb/VGn9SneKZQN
vgwZyXEdTuOQceDOd54nKKyghwNwFGOPz0sYpP5zsLdf/MLnYYjfvG9oUN/R9CHaZlzdcV2CB68R
CUyRlAssqWS52a0O1wFEuUwtg+s7gca2IEBFgaWcW48iIUFlr7EKpTSSZwF0NV0F6Mkua+b88xIC
HSVoEvGG/z8k26GS67WInqY/f3FcFC9K9U1HM+4PcAxPkpiWpbZnrNOuucu2Imr81J6G8Pl74Ol+
jivuS9rvqoLpGdyaesoNg6ZR47Nplasr5YFqvZxlbfOgwHDOd+5e/xdByK3FxY6ORXHaok5Mbqc3
CX6LkepMgmv6IjHqClpi63Ggt8nnULCbQQTWsV2yhqFDPdi5PT+nRKvzdCYqD8ZxzzDg8FyaKkzf
8uZY56Rql2qj31HokEdF7xhKRy+/rFRpM8Ep4GFJrn5ZDlH6sGmqxmo7H8hxixF1aHZzaOoM5MEj
RwrsAVLN/yoWSh3LKS2WpzQ/0vMYPsZ+lIz1wXvXzUXwfGFSteM4DYG6gSq55BqU7GMqSa8Dmsah
I92DH4FiT5ECrUPAInDsQAotb/gixUxEob0uyiAdtHeZsfeVXV/k5ky+DYIiXIbhCypr02OBCrcb
U+D/52N43gjHQmuknntVg3bvDAgqujwkmkcFZ8um2NQf+VT+W5kA6AHplwkp6gtOwYTQdSYq8ZQs
LZeEGSzCKV1hwxqVR6I20QL0AKbf2LQGnqZfGVIp676VrghuG+SUdJjWrtQm2I5CcEbxCkofgpgQ
Z47DOFauYiiL2nR7xRrs/mFVha3qAz5dzZqjXvL+hEgMQs16kvMYCcP3mQ1xn+2Tw2ox+qNDTIEZ
SmHyLs8ftBq2Estjl29YE1eRnz7y5zzBnDhfpTq4lLZ+CuXAeKAVnWnmsKPuItn/LYlV1tBgJ8ic
bATkkSbOKkP22UPdcpe8ONV4qEPwO1OPIBJ9dLMsGa8wNstS6gXfV92B1szJN6eFEZGWTLKqRgVV
NyMHhlIzDlNTJN5kiK3sfpH4dmtxdbPMKqEVpScMYxf60t4aXX1qyKEtCz2chWeEGrMxN6YKqZJW
rG5QV3xU7oesabCGBOvE8d0NW/H0qNJSBX6Cet202xrq9mYyAJmamVk7Lh52Rfbc4wOqaMXmwDlx
S/GAfxyvPo/C7897I4UKwu74a77KC6kHhnuj058Q8TMIwfaZFm1FCH350wWf1Sq75tGjUTJMxiPD
F2fxD/C+k9OBzkK3VLCSDqn+9ty2E8DjiOrsaNSUWDkkQgaQFfGNAd5QGtE/zUc4iCilROsKRhxp
hyC6UAed1ZSb1tgBRYjCV5KdabK19tGwcRwj8h2fhQypVIIstTOuoQVeMOg2ospu3opyzbX5kI6x
vYMg+nzKA5c/zcOpy5KW59kM8RVLxI9omlqYo2d/JdAvG5vDd2VUIrGqSicr+vbjfAKt4Detbm6v
sOvO4GoGYf74dFwuSIJS6s0OTboflk9OlEWYDYH5P0zTLMv3XIER++Y65a7H18CFJEQtDH28QBvy
/MXBDBoLYFeZiqpEh5wUbZuS5G9ELxEPt2C3D7RtASkuMVkoEdL0GnTYo28Tq2REII1d12MjNQPA
j5Dq3D7lef2Ow7qSp1Kr+C2NsrbxsMd5uF6zw9CDFILSamJqYqg4JRWPgvD3iuGitEI+zO5r4O44
nF2TNx63LaT7LQTbYVnvWkrr+wKD0mL1MoNbAr6cvrW/M7eJhMJLt14Ds470TeQra30bEkmq/lRc
/0rFPE2yFXPl0hpc8ZhyCpnHuZSAhEB34aNr9Zi2SHXzLzr+V5gXjrWynYXYKqxSD4BgTZDSwxXx
ZGf25HzEhlazdc62v+j+QKwhCMx8onajnqdasCpd3wN30eF5hodBL5s0DZNkBfQCuIHUqej5Vh8c
YSM/947m2Rl34OkvFZEfoT1szwSoTQHifro2EgeduZnDFjNHmoN9+NieaCVbERu8FJ5A8h5v0oxK
Xp4gHnToZF4cMWUrusbCC54dNy3qRanLbCEUCQAC40TJ2hxRmSv4YKdLWqn5NLH4j7bCipYRwYof
jeQtfA2ULKy9vE31IHZYuoRnojrYJz5BrZauNCgHmTw5x1zOgFzVmDpcs930uSXofWzWSurueV6A
AXFrwbgtu/ARq7r4fNJRpV1SKJuH6Vnt4lAkOfWkMxmCffQJFtd1uathVqawjJR9kp8ZRHmh6Wj5
NblB3e+M349XPUjKC5NWKyi9VO0NbSKDSAj0mH6coMfN33IZx3NtgTiGvhE2R3vfHU+itMJaDQMU
k08VMn0A+ZTsb+i/qJ/15Yo5W/XUys9/JtLuQoX0y2kXyf1S4QkXpVLJ5HeAH/YuZIrKwSOyxZRM
BIBUnVWJPfUKmZrKG42CPTXB3Al0CUBSW/P9+WcdTLyEaz5Q6RtIO+YU3q0yZwyWuvvvvaBC9TBC
Ckw5TXKzeDPBiM1mBi4IyrEhmjZ1b6mZmG4xJ99shaK0fw/Z+s5JbtClq/BRv2+ZTUTsyK8wsI4t
zp/w3OHu/xkxd/GCuTdWRrOdLp2ypVQU94aHYBD190eHAVDWAMQDg8fqow5FcLq+HWeUF6liciBT
P8JnGWLaVn59NY+UgZWduPGbeA6MHHTjiHKlc7D/UyrzkXdKFB9QfArAMirx8Uj7kyvSiLIBeWKU
KpwRveLWryBz/7xrNjZXW/ANwK0MUtBaeObF4Tblqh9o1SFCvfdS9J1RrkFECqqi0eQGCpVE51B2
E8Ca0zzBzYBw8GkbYb0WgT/ZVViGzatsFaelnUlpVegkFAieydITu3h8Vatd3MmkfhWg/cHzHUpv
TjCM6Am1vB/ub9Ia6QuKkHoOk2SfjDeTwh1pMKaAvQ88SO+iQEEFXBxA12gjni8W8WZCrGD/TRYx
iGwg1r5Z6MTI691X8YPpvZVwt9NPopbMguGiNY8OR5SPQcAICpGWUSiqghtsy4hJBb4dYAUbX1CV
dFDiUxi2/bUStZ8cHc0KO79mSn4VVP2Xym3Y2fLJtFHHZziZ73luIhdzfUpFZ5kfcEbLOIhULXTL
0IXnOmpDVG0N8i1t3lHzVttCjKd4dtE+VXvStABgkthVoHGCio23J64CXRx7ywsvcEEzK/xqziPt
PgmTy23nZgWh5JcDQaVEe0iURZIhBRwucAmKyDOXGQ5WJ9Y2MhhNvqufscUGN6hoi2YtfLnDIbK9
5OvP4N36N9RfZ/d/dBpwFALzfnZXdR+W5HildCimNOCuipi1GeP83tetQ3lEorM1+q4hHuUYQrVJ
6lrj48INj6ms347ythrnJ75XpDFvC4oJBszrPvCBr35zDV8uAQUDYXvkgZJ1MI5qruuyZc4r/b03
UEk+qw9MW7rB1oojyza9RTJQXd9NeMqkof1rJzRZKvxwR4U7xBMlNagWtWdk9wefxbBILV2jVeGo
e/vKzfmbeaZU4qwNfuwTszliSL3pRGMGAUJG4Ft7IIZTT6AdAR5i7rMNv5Bnr86VgOnbKzp1uZkT
O6lPTE/7nzdULD1xPopH1+oIGxoVUDzx9Zt/uzVvVBaN+7WT52mW9WxCiGilhf/gNAAxwPi1Q1AQ
cgpZQBG3ArOicAB2/LMe7hnlm6MgITSPx0vq7Ozh66ZZWJ4BRR00LNtOVwafeKLzVqXniWUVci+p
uf4yeQPhdReEtnUbujGumFOFFUrp4HDcgLgwiC2Fbqtxh1thYPWznhpCJqQpkYCNdOIk9k5PJs3g
i8aHf8CARbYyysq+sgkhvE/QHe1J5ueqm3Nh+6l0KShBcupo5fUy+V29rs7EKf59QPyVN/piEFbE
03sdJqkN01vTX7TB9F87Io5Q5FJUkpU7Dm3ol8y9/Io1k2ioY/nLIRsx+wsGNuyT0XN7OA3AGbiL
U2FvEgYcg4jFZGtLZq19u/xQfPk8d9BVD2q39+OXfIkwnBsIgOYDORqloDhHYN+ij5opOSCPqoc2
b4DdoVWRM8DhJUuz2XWBzL1EkoE8tlr4BUgH6asSGV028KSX09qUbP+pvp0LIapxHcFU02ToaIVr
vCwBU5j3H6q/juLFZKR/vy3gOcpnJHZxASbbjYLfzBhVrYhbUAFE437oce/tLZ3GGfJzLrZe4pp1
zaR0yx32xL9D2PT2Da5x02d5S5NdwWMYyDV6JKzqEOhS8/G8DxdtP3orqISV1cR73MHUVvwZ5P4Z
3Qo2x/d/99ILiSGUOYBiTWOKh+a/9U8lUO5/5HR74YHyXq9/K8TkWnl76BU2rOW2Vac9igWlAntM
X0VK6kj1V0Y2EPUdb6via0zw5Lqs82dtBCIVavvFtVx8ZBzS6P3P7D1DYPf+atatCf3PkhuepvDf
6XO1838vz3BkNxO+D4q7Z6hKRi2e3r7+dfhLIw5RC/lu5lNh1k7kZbBG4t7E1HdIP8JK67jnbWF4
fhtxA7TTj8kuMYStddFN5TBtZiAVmJ5iYwvOwribLr6hRobQPiluZevmrD7P9NA93RwrIupKRTcA
9jes8IJXsKR23UXSd+wBCBosCILCPa1ohv3nNVugSI9bikO/ANFcY9k1sugZsxq5JHkMew2Dm5vx
10tSz6jl6xZ2SSQ/GuyOtRI7lGqjISYyfwMi7vrq0NQMpSGSWrrEpaHmZydzQD/FtZtYjrnXGLmy
fbUBqm8TpN9WaDuEW/58L6zlz2F4NI1raeqtL3ta0rhnjTjEJCwHhYkZEJiSDy9riLoNDn7idywA
Qq9bRSHEhqVOwtspbd0qi0KZxt1J6okg1CakuzfWkGULbsuVAVdCHRkgrEulbdTjLrpxTYhiNST2
E5+TELlc1/ErIc/Hxg/EMWJo0/AgTesrqt9u9+aXkcbArD90IukBpjHDXAnBY096IgWydt+BiQgr
fcQZvzrGriMKwFCOAwt4hJIC0pjSgkrXCrSRqeXZjeJOcGSXqs7mqTDRwlUeAyATkurhZTyi0Wax
QVAmJZ1Tb7aeJv4spjIXkvGB4dN8ABd40/ypZNQCP6BjP07rUph3NUQ546kAxrJ235sOpPDL0Hmj
bXTk3dahe7bWTgPs3Y3L4dYmsGk1CDyKk48KW4j9GB+3YZjYCkhkXGGrM7QHfUv5zywdgwM/92m7
un4KNWpuD+w9LTi/4A+OYMqmgafGqkWVWHy5UQymofHrJCsTL/bOPtNGv37hlA6ZTbg3BB5M+F9b
3NcOMuo9vnVPRhf8MLJXqjalPecftZTyliHlYjTnonBS/h8JIEwyX6cMnzoPvVDSmK2VtQLZBteO
A93QoVAt0xHgN01dCki6/UTttdwGfXIPCbRsjByiXWFB4qdLC11lg+t5kEERZkQejWNpTSCGBPvR
FgaVRiHJKTayBscl/xL/haMXNNXJm1xXnCgXxWccTNeH7zsCulDk30K7+YZWzRzOo973OvBBoS/Q
T4M5VH40dk6AkE8t7vi+xGBC9A+VoGFHU3GoJkd7fQBVvRPTCKV/i+n1s8yf5vHlWfhvB+fs1+Hq
z0qndU51utEBHmusapTtxbGGIvywgZH1mc/W6/NZ6oT0wfBhzl6FQ6f3e9mZWF8LPOTOIFNC8MUb
DlP6EiTs+qwQw1coRGcP5KbcpHSbAcpENR5zzwMMw+U8MpXPDnyFrv44VK92ioEp86EaLdbJBIlA
2rKWkC5xQR0f5neQNa9V6ocKu6HYcrWWESaeZjKMHETNVrMoUY/pZc29XrVPp4u5JlZi9hMxqN2l
3wATtnVMEvuSLFq4YURSwCgQ+WmZY4zodd/cRxJt/zlhstzURyvfrFelomcHcrYsaZZDG8gPEsqk
BgJJwcRqal1AIj7N+9Ku1iGFV21VaeVzbPaBv0MZXawcVU/p64DaTOJ6aXxYg6paUJfIf1gl4wTO
721oDQC1qS5DSr8WYIQ4Z5b/GPVEW58r8gssrifvk36CJ9YXsQaYybsGxqufAhnJl60lo4V4lpLE
6sN3ZVUhNiwPFtq1pIcg3uIzIJzSfZMZlvZynFy3n/PAUSiL/NNzqp2isPoE4tMMzt2E4ie+XBFO
3Prs4nb46mUDg2B3jMQRKOdIbYThisb+N6RveOpIh0YKACR3kR36/OUFiFw4Jz32H0/RK6+jX+Oe
nvXqTG2jhCjaIgq+W6S2tSrXR1z3fO4g7K63X4CZXT0EcjWjfJBDevWXAEF+9Ofl87GyqKrc9YYy
BIDtliuOtFFGndbJxr9m47XkJYdOXnmP/GtyzxsyQURPIsIVDXANhjnlHW251cC3+IClcWpv2pBT
Wi1E4I79FIV06RxYVU5HXnkLsanQkKl1w62VhAxAX3baH50ceUmlkzNKlrOjGrlQSlDJ7sVsfyEY
HKdQbsK6xJAvBmLgdTYTCqmieVT2C6Rtm9YdeS1kH7KbSdOEHiKpBaNVAZaYKT+2IPXk5OrNB7V8
qQsnP8wX348RRbzs9+O/jaJB7CN+bTQjyNCIQw3b+/xzx0AsxzvDFRIBkLqXoKqZidsVWorV4QwC
hH0JpXtkj+92qtqETjnegkDqFBausHtsGGIlRVYOOOwDBvWZcKqFi0BkmWpjCCttskb4RpvuJauZ
nrvW2muFaol321+URiut1//i46dB0vQADUf2bdu9fs3tzc7fOkc2f88DCiHTF9CAWQQruQLQbWoa
CLATBxZBQdd2aLiZyxOTdaRqgr1vzv4nY3PVHrkyKMrMgogT5G+W4JQgdm5u8Vo9Phj5/irImlFY
L6H6doxNcnkms15oqmnUvnnj+kRIITkZ5lXHWKMOru37wP2Mk6AH60iJEU9PWvdHCAhy/UUYu/iP
jwiOT/MUq4/ZDgvD8NAkE92hxIGhzGVjtR1+HMQXv+6GNLbkXgjF+Er4KANrKQkoJlqP7HYyDIzh
8Fly79NEBYQNvvFKdNvoZaxFito499HoqE+4cWcCHebbOnH9ZA/nKSeYr5vnclyd8l+cSfQ8/Mmx
TzmXgx2ySHpJAwj5XOru25To5M+A4ZuTq1HFal8xndGF1ECMe5k0IpxcxhHvGu2HKZs90nN9d67W
ssHdZDvupJR174i5XzU5twIGf7wkiURhNpOAMxDc535bpto5FPyCyvdpMRaFq2jXRmqLXwikdCMl
gSwzPyEY6Q59KmbHbc/S3Hhsu/e1Hn01DiSBtJDEruDQI6eMkbGZ2zWOoQwoie9MzRaWJaArnZB6
Uv55IiXwhGHyKKAm36cdiu/SGeePSX9nSwl1k1CGccBaM7E0bEkJHmLfCjyh1Bq23UWzJk/zl8rf
ygKj85nBsVQu/+/x8gNkal4W5mMBCKT3Gd7zV87qp4FhIZ2N2cA1tqcrXSOAhBiPZbpW1myEEewg
2sHw4SJJN3nL4+U8aH/c8whZByU6hqtI9XeCXY/k1+xmCc+mzbjv8Pc2GsWBOFYPNkwvC06TXTgk
sxxTe7TXJbQ48sqZmjQooO8rYnCl8cFaDuxGTjA1+hxZUlCSYYDq2ccrLqb/QVjWGzDMhHB0ShHM
LUh3BieNOKucMNYzPny9t/xJlDU1UfRUwMrBsC60gUjNceqHwcTB8QMkdCIu4Ub7+qZP5zNwJVFE
EZyhgnlrWHeyY7KRpJ7zM05ZPRqYh8Kjflj/4z7kWtIo6KWtH5c2Vk9w5H1yhY3fktlbA07gNi1Y
ZCMelcg2i0m7OGFIowfpjHB/nbKIGu+AWGAbXxTakutWQIJ+vmAJCijLnq/ukyoM8LaXC97co3nD
znZUR47q6xj1+G8IXfmAIUkTrZkEWIE1NJgyBQt2dO7AIZC9n2keeX2ypNMe4uLquxXbs+/QQa4/
DSkwegG+x6u25v/LLba2TDUVZpySwbU72R2ewF6tW6AAy6eLkrGWJE0oALPlcbIbqidmVFH6YJJq
wDEv/RyOvL1gHdWe4meBCruI1CHy5FgofN9OceclYsfRSI5mkmamEF+jPyKztHoyQcIx7jiN5wdR
PijPUHhVrymgz77bZ5N2N8nUQvtb4oviHdSLT8cIhMTS4XxsE1z/YeI2sTz5rPT1RBdlt0HMnogk
8g1BdazcyGHnfgIOLRBlGxnlDh/7sjWQ1Qk8vul9qM7yONxdBMQ86XSfoz8OLR9NlOmsMcXRzUi6
plgV+enyQTtivnbbEPvIFIVtU7NkJD5kG4W1qMuz4k32j8BaLztbIToaENvYvm2TopCBarAZrkga
g25uldvxY8U59KxYgo0skPIOOfEgYz89jccuNLxZrctHq4XwAfVh7ruKFltmfH7dtH8E9DYlQxDX
/tbdlpx/HmAwUkt1eEI/CqLkzvzEkJKOo4EFK70PbsJ8XQxas8em8uVzcGZBSJ/C6NHXilVLxMJx
rVB3Mh3CL8fCdP3776BjtruosI3Qe1pS1GF8GRwLsk1fO4tGmzXabX89AbQkgQMSkYTx0OjAGIsI
V8e+LO0j/hqpWPa6woRSwtJGZBQn4k7ebSVB9O4Om65RLjJdF2qvGVrFAaihK9sO0/4Ibrargv9R
NxyJnQRP9u0RPtt5IMbCcY3JT/P4WxpU1VZMFq8xRlqGPIRGXxcTVheOKACu8Xmpjrn/7ND4sgOP
bHJ6E27Jl58jwVz3/rjwK6xh9puQSO01zEjIrw0l2cjdg+umnaeKHCqAs7gAe2iNa6XEDQc3uVKM
2NanJz29mchhG87JjUG2imU2+QXNbo/HnT1cgmpH/Ht43K6j13evELSkrlo7HcFhxo1Mf/ggUFdu
dnzMijTYKR1kxoI8tDlDJ/YrLQHSpc4agDJuCPvrPDGSCivW6mwzfCfhmuZQvpYrjB3JTb2MQ9CO
N+2nA4PjrjyfjPt0Qy4ilVgOPHY4VKw/DwiwygRV2PXDJDAjodH1jNdQv6l+A2W6q/ohQHtr5aNV
s9ZxahjgWTCg1vTw1hnJiiANmW59E/z9ZsVv5Emt8NUDW4rqeCYU84smARylzPyGZhbhVz/lAjXv
WdTwmsVXi0Cs3fjURtd6c64TPBBG1F2N7dtEL+GVyCqz3xvIbHyupwFetWVuqnR/fidHYzvQNavm
+rNxIfE6ffBxO4RTR5SckXV2309zoMbFcMAOvJQCOyI5Z4lqrLpUaSRoS9E0da/72PGLhVfECVp4
K0/6kNsWgbRBkhzIOQez+TxO68dZtFqDoSTwOxJgqIPaGBazlxIBgAg2aFZWYGWpTCmPyBkSbHb8
gVNbTopP5i46+fgguOZY7E4501WflSwkCSApO5jn+Omo9hY538iY5L1r3dHEiH2pAtS9el8kv/Yq
y6KclpfjUc8lbVuCsGRW8fiRHrUwxvCuo/+Ff1i5NuDwuod8kdgh1kMMk+Ds/06PqZXBq/Jg8PJ+
h/EPjwZA5EVoqxa8Ka3zSJ1SFuk7nIVaA7GVw1XsW+t3DNhd39xCia24rLVbzqh5mJWd+8rhlPYN
kbpr9YwssJw3hCCAhgDk+PU6u2+h6kumryk4STUcBexA9b+SzCxuFMZPMjFjrs18TcfMEIdg1/Vz
iuL8Jgu0acs1ilBV16iGWmqSjTfS0yCyHOzGdKm12fFYo5lCtPr2pJG82m//eiI7AgvgHWIMf64g
tPfiz3JP+UFaegbvnEZTIRWRPfy5LM4l63Kua2PzAjRqCymY/mi2qM0VPrKqZwdQbtOJ5/CZeqxG
KJbFJRTyU/5cTQKuG4QWPGnWvdNCohOC9iuqSSsi6hmYHvKGxJCjOdhXR1Ts53HQJtxCSwXtu33B
vmURudVos8zjUmBYXqtfCL4R8dVeJPLpDXb9h3g82ftcvd3a6kcpB54KdRxTOFVi3C/PL5nIqy04
/xc4cx3B8d9bIBcIvYPEXe7G3qy9M/lHLhS5i8ay8lQMDu0Di9VCCjKkTk+7AelZtXVzMkog/mNe
iFL/3laMeyZXViy6CYoxHRdf4PunCyf2mY8VAqHVZS1/Vm5Gnj6QIY6eeQ5uj8Wiaaa9j7w7XWyl
zolKFxlb/VGifDPqR6BjxlqfZp+SoI6doDimO7o60h2JFiMgV67jj3AXjTU/HT2bwNkXxH9N0aDv
81ERB7/UpBUVeqeBrkurQodnvsuZ0DPU0TIC9XdpHknWjJQervRUkw4/7E1fzjlmXPJeTRPEbAjW
Eh+PpMpaqHQ0CDmUkhfgWdInxnHxxcN5+Xe/VTt6k1wVOF019aX1yc+aBZSdZ2H4LQqV3w7UWtOJ
Obhu67YbT7NBJBgUFnxP1RO0OK8n+RTfpr331OYyaAN5rEhYwfdR3opWjm+2iGMdRwXExaMVdx1s
lCFelPA4c55b+Ht/Be4IVY+Exe1hBggC9FqebpflAUkoZfsEBJAHdTQLOkm1zfNMqc/toDxEwxgO
bPqW2PUI3Aa1DwQ9uwQpOr+NDnlWQ/pxt5FcYy4sgiK9RoWFLlNxqgHyLw04gvBwyTrMboflUfgt
JckJpW5nKZ31M0EDdea2K6QOZPF1rj0kx1zaYRtdem93EEQNut6PN+lsPOGkiAjByjwscjpozHZS
0gWeXr3fBu3vTOpf8Er4zeHQfXe/0zhEL5oR3gFrLutq+QqTP2oLqHhXo/K7iiZBIqSZ8lCrgEj+
1bBvF2vO/WCBO81N6RA42UiB+rTSFlR1vbGxLi98jpO7GQfiqj4pSPTVN1L9FYgJWcucASQni7SW
yvupJ8b+IVV48QDncAhnHXFQpblnaMFPu/bYKzkBBquXZHS58NGwJdrBA9ZLEKeK6V0V8ouiNBAL
alDWXkFu+SB8h96TXR8fypWzicZkKblyhdZIRHrU7EpDky5fHMDv3JueSBQwWqLEPvoypMcXxwJ5
hSBWp3i2xnOap4+1RzGm8uj3SsdPAZKMYzyOyhTnd0fioexK69FOLWitEdxcQB6fMMESGack2DMI
AgIVMlVR2oB2z2Y6ciWSYzTdRzjNm0V4j8eCSTuLtnOuhxpLkUT+BIjuXQuAtnm7fG2j5U6haE7e
WWvE3hmwvkOcHDWaiwY8A2j0xRCvDejKCZsYCfb1LJjJ5UL/AfsL3Bqauo22GSt2UNm5Hts/4XY3
3DIGypJ+bABcRmpDH3e6DhfEC7OdO2rqdq6/XW//LM9UXwGYHSxYfVSXcj/QNLG04mEfLlaP2pm9
SrIOKrgwa5Oeaquk8v6HdCswV2mt4IHONL8YC+M6RHdXyfmnsdLBf3UABVv3xqM0eqJ+C/TJAfqt
2/EvR14pUUmexM+dq/J7eREIwPf+Wtt44kSYxGZ+tBfJ9oX4BLSnvpMqUx94eqXTiHP9wAV0ZckR
h/Ego9QwiAcQPnBXLCZssf1Qa5nk7zUIxiXjhw6ufUFFkKoxqbKgkK1pw4StoHPV70n4aW1BVTJt
9/hbvF7o4+1BKW60ykD8PFrrwEQD2OZLevHWSalCGNu3EZNEayIpUK5/iwJ1qzoFKiR4jGHXEIc8
pYT4ZKgeM1F59vr6YdVyKNbkOGg6+jGXU8glkGdq70ISVpFCO3nXuJhh+SiUOaWONmb2z2utjYb4
r9uQQ5PJveUPH8dQsC/jcWlwlbgcKAUcypQQakVQEXMbvmvwfpLnev9sEGV0H5BqWP4vycjyq7o+
qv58EHRp+1jGWwyo5eCqsoc3WNV5umMDcVLRzIGJtIcqWuM8FBeuAs5gjJczbqS1Lp26xbD5sHpI
Ftg1VSL4EVi9Wia7pWulvt/pYoqVQTzD4NJVG/q7CUxQ+sxzv2rbN+mZJxg/NQzfKF32g8VrfEzz
6xLrjCdKq4lgSTupPMD7JFFygVQ5POuv+HXPcCzqzuA5xECUFomAcPjDadLq3Yk3sSGP+54s+4JR
p92MCwQwPOPNIOob9t2TYPwHhmwdjyeKZeYlkDJ/iXH/yL5hN2Sglo1fVPPhsDpYV//IFEmJVJPx
KRGhLMwpZMkXStBZn38ja3R+qDxdgl58kXfG5V/aAbNgV3vURVcIn5m2eHhYaZIiZmrCSWyubekJ
CFNMDlIy3dX7xWyqCJukcM7blUmnpSoSe1d2U/SUuPywKx47T0uPLkUJOs6VsVWyh6KAm+hMkxKE
PiFedxvB5eNEaSv7LIfl7wls7fiIi7CZ4MJJ00IxtPgyZG/gEkIz71TA/eTtZ1fbImG3Nhgwp62y
WrPLw7io3CTe5RE/ZOrVTk2z+kjiKABoFABGOzf20DYCvZYWE7joBYpmHbmayCIyotJDwnX8di35
bDFxHez+qW3LIpC8aC+qir3Z5j7v3Hs6oxcWOxgRr0yrl3NEj3zeI/YdhSHPQwF2pN3IHqNaqjn+
HeoFhTOJc+X4wFbzJK7ud57gfY0PaJ3l90qHrRo3T3DFV6gr/KdHoXpqKI9s0BluHmt0hHQKeSsQ
3mTJW+yMXD10Re+kRkKaHh1dCmydMQloUtD8ZoU8QkVy4bd2mtukodji5JFxnZmOpT9BkqCcPC4E
du89zKwJmwQyBL1UYS8g/HDT7qmb2wYci1tpQdYFKFqVHlWIv7M096IBoB3RrRzIPD6F3G5U0UEE
tHOWNZGVnsQ2CWzC1m3Pt8Vp2878BRnaXcgAbU7kE94g1BUfVo1n4obukjn8pKxKf69WwII+ML08
kWAwAhwiEQ0N44uiVN82abPeo7Aw3cgpHQWOJkr2Wn3Bvm2bIacCGt+cYLpALwXdj50FsAeM6Rty
uhvvU0+tRuRbueXj/PDq88OW+FSIlhqR+Kzcrq3xIGdZSTPC1hy07zaHkmxbDntqM/GXZePNJl5N
EOwPUQFo39imSVlLctDN+55qK/OMe5083WWScER1VvZRkmQs9562gzi74vOBz5j1q3/d9iXtCWD6
S8aIhQE3G5s74wW3SfJhVoCOUpypchf1VriK+XZlEt6bAxonA/BLDXFheoCiITjuFpWPsIFP6pgd
xf7f5beQfb3g8h0NkkefjnhksPr40m1fGyhbye1fqY1Ixh0sAoJd4TJXIa8GmvqXALC15aXonyNO
W8l58A43aYZOdBcOmA6Ey502YGys0jKNTV6mBs28rGMafonxqwNgSZ6DjLguV2uNHzK+Hb1Upyu7
vz2Z6xBuLP8SCOxSfhWbUtnUXBZcQWlVYdofy1tU/FSf9kMamyiHK7333Dz26q6qUexFzmjs9QJZ
gE8bSxNRCZbx8stB7hBdRqNfrAtU3sYhXJ/TVgtVc3A/d4K+XSOqBBSrgE/VQ9IKPStTuzrvkm/K
y3W/rL6Wwe36t2Q7nG+LgBF51yYHrVNPbYRXzuRgAVdZjsHEIWaWvdHBySEPjPKwEbh3BJ9cFrxM
y4vzTqm41zKH9CwRRzsx+MvUN69yJ0XhGG+7o+BGs/iZoWSk7V8eQZEHIn7w52kXwHSIv72+gCLw
JwoqoPHcTcxt08oYXvgvMIbiUj5i4FN/7kXMXXR3vumxjbJ1cveu4yoRQmlYvHuVClS+ta3Pj0W8
WgNDTyEHPuY35NdNQkpwY8P1KeWhm2ZzjFAqxt6wnVqmD20RjH9JPACNul8ICnRVZ9w13oF7HVjQ
SXil4ZGiWjua8iX+4Amv7WMexoEOv8fmL/v2sMg835k501hvPthaSljvk3SQ2/6RA9tKrEhRpWyS
v38EtY1iYj9PA2aUwnu9ThXhFsLvOaOs/aaFfaTcJBk3YcysrNebxG7W5Wwo3phudgYIpo5Kc0+9
vUopbp8gX5CDpeTKixjBzjJgkMoV8Gj6dcKYjzqYtpOUkyRCFPccv/WOVtp3wlRVaTQbHQWsHJu+
Wc6TqKMbhTz4lYbxgF2UE8WVT3+S6P7IuKIVCtURfwroOEveSbJpXAEhrg4wlKigSPkKki/00ulr
IqXamjUaMQoC0JFPT6ivZoW+BARCoqE2VMmIA6X1ySST5AYjVPIcYLWeKiDxrUOTWFRx7dozmtF8
CSfbxFR4jLrG6veuo8hu/Q7jZCCxQ9tzXsAmhYyBtDyp3n02K1ibxXdFoSYSr6R3IstynluKhNSX
KO/SxeJNTH94a4necDZ4/lZDkSO9mUk9NxY+8jIyDIusGRT5QDwbOqtH+EJP3a34q+oEb+gS8VMy
LJzlcQkiddM5yWM8F3piBEZs47m6pvd3ZoMqoBE/4FCLuQva4q/0OO8AYgCuyLoiDqV8DfOBbDwQ
W3EyV1gfGo3pW1bTZOoJZPWkOG0+YJ+fRfAZkjpbKLbKxxxPzxDniTSJCIm2v1KmylRDqday0pe4
aMgAXmh6+KLN3LFpPwbmObc+tTfiD0cMGEEKuVlZK157/qDioZ9v7bG3t7uby06REzlBauST0UDS
aWt4vjodso1RN99f5IRSeroUwOS6Z/kaz9b4MlJZJtpMeYM+vqR3tTem2Uf6npIOM5kHw3Qu5xA2
JzAShoyYSWKjqTe/xvIJgPS84eKaL11aEb5Y91iqV+SX4KT+svxjQklRhgbNcj74EGsCrW8GMrbA
v4BFnn5PtNig0hRDAwJAeIeuU25IvbWzNWs4D6be0X2YksMznwbAvjfBsoIWdZb5FaMZ7UMb0IPF
hTgn5E128fw0im+8f1q5oPTbCJT21uSF8iHHLTrTHdSLT4RWQkAEpGXkMnxny6qWNYKtZGXgQX/E
094vVGPv8HuEXE89AV1LNAQzOLh4kA01qSNGWsDkT1aaG/bFbDe6+M1S/fYJ4QDYrqutkEVx3KRA
UYtt/NWQGJv+62drlW50zeJ5S8JHANajOrem7CRug/D64w/EQ05/f7n74J62dAdx9BthWFMowCyO
SJWgHxtUM3T/kYcBfsSxuZduk9ahK0W9PDSt2U0gJVQEdyEccrcU3MImKTCZMduMbdbO+B/zxQjI
zDVXzMrGjqLJKh6ptoCEhPQfW+1cI7JlIXRushVTuj3RAT87cRpBnX3CCTAjE9vMddjmTSFt5VvH
xmW6lyuEoBtW25ydZqfr5uQI9N1Uf5jsl5sgKaeUyqjE3hUwFXxed89rpedShZnHh212PaZUhWJ/
PHcSh3HSCqwXAmH/G6sQC3XnRRJcyHmbnAc0EAaAXckiewyc6YrJ7V1Cy7whhd2wjYhj8GfIln4C
s/NXBa5Lv5A8KIQNYX3J/ma9Aj3vyfuLnCbz7bwi9YVKhxaRhFel7fv+KIMnioLtUHW7HR2kh/mq
D+AnsLfsqmC6hqv5+MUlgmocwTuHIuCpE7dA4ivjJWCMImN63bpuu/GXoRCw58bYOFZKyAH4FK7P
zuUcUCDzklDePsw/kd09bZlNy9kXKeQHTNzsAUnNaZUysBFbK8NLNO4a6RIAFm7B/EAHtj6pjn9r
0KyEPuPgyIVZNeA8EzVCNiGVXuREQ3VjKsynwG0yuaAsABmEMLRxTWIVc6lW1eAxjnEUwm38pdSA
35LAvvBs5jq77onwdaGIKO65bzUUVHdZidyl7/xwWcRW82t5/cHa8ZAnv6LnwBliPUX9xq6lIXbu
HmuDGoMLlaZaNZBc0DLs6BNFuJk7wLVbwo0iEVIEDD64TPDtuu2PV+Ah/yk44ws9KE/4o4BOBpHX
BRsNLv9YRgS+EjJNeQpdY3m+Y1mUDP/kUV6O1GfLtZGCa/kwRU7dnPXdMdtvoaAVXxod/Z2h4Ocq
LIDmyYDiRq3hRzioUASTRS/TncpHjW5PHCtvKmtEoEJ+O+BnrZlTNJO7f2OVy/8QW0hIwfZ4UYX9
EnHFwYVAg9h1zosXEsCiFga3qZXdgxybolg/3Ksht4s7tN0q3Bd+53zYX0v9Hp0YPzr9MxPwQdEI
NDEEv8vnqPSbHOocwJfTX2A1R2ra5/dW2THhyJ+gwq8wUHHRCsrNFZtYSwcxXW9bsr/iAd6duTDH
0yYmuRLCSsqR+HJAUIdbMKdtwnN9/WbDqZrkdd6OfkxXgiHYsoL7PUQc09tmdVs/z3zeY1RUpd4n
VV7fHD7aH97S+1jhyil0Bvupw6FpcdvmZtv67vEN+FJhIyWli/Fntq9tvrNP71bDskHO5Xx1O2rg
DivLIHPKus4a9PR0Qmz1oFYNyfaUloUqlm95eGcNhI04jJT0hOi0YjDa2a1CEHmAgNSp+YeBRtru
pV34LAhmVTiSyDhTL3JF1TokEuD5BQYiY8pLDYzSQH8LNAQlrEj2TnpY5E0kzBAU8nIF1nkfZG9h
yzI+oQUg8xS/w6LHqh6QCpLWVtI1TnWye848DedAz279jmPfhv7BhEv4dHtlPICLWEsIZXNWSwpF
fdlLNFKGQqc5ZrGE06kRCI+sjzdRMmjSc/SoVeKBJ3GatD5C0A4Uxx8qp+4TT5pN0UrwCnVdfGXV
ZtTLR+6BYjvjSWxZVmRhIBicl+S2WvHdf/NEXEKVWT5QH1wvNe3ObHwA8y7iIk2LyNwEEpKtMIAl
wCMJ/aJ4Nyt8nBhjyCqaBSdl1s/qRN1vxcjdQAuQtylq20DQhkN2n1zaevUuWMtmJL1x8XmZRRF8
9+ZMyMI89PdNxd8S6RAzNjagQkbRnTsvaM1Y/V+hotWBTVVtogoOAUqRiWCPL+v9Pb33/VHg8QtN
NoJqtlAxIfUccwpTRHRFkiT+pRPTI2LDSSKQrYByi6FCcMRnCAWofbinDg/9IamS1aNNNzyfVs7T
VaJrsJjjZHS2DN+7dXI8hpPDt26/rzNHY+eawae974seGg7V6MzxD21QsHm7zxUh8qC35dedqBDB
4GgGaYoE/ZmUModlH9/Fq39QEBbMTXDgPiCbIW/CX5W/SKoXw31Rd7e1XT0CjmnbtHy7PWdEQcTI
Fq9YE5D5AUqBwdb1CFddbKyfFdXtxWQ3p1KZ1R+Z5EgHb+XralTqezpVk97N98oiDrwu4w/5r0Mq
9cMqpfq3sV1K2xbxbHEAuECuLoxadED4beNIwLB0psIjr+izu3Aaaaq8bkpwWSXUOthiNJRXPZBH
sIqXLoMlLevW6+k2IppP02A2RGdM91IlSL62ODmPx4FNp7RDmLNFrTipXsAOnZU5i+q89rcptbfk
YoWdakll4ENpI4pR5dBH5ZYPYs7XaBd3pvu2vb24npHA/Z/q9Kwv3jCzr3Gd4aafzOMCv4YWhqXJ
d/QUqA6C873Pyl64S7hdnMRNtT891d9TySgH2SW5LtTJuyCCq8UXBF0e8PjA99uvkoygP1U8Npzp
mcQepdu9NFv6lkPNsDPr4UjzRRALrNn6lJ/TgcI5fWMURAmhpygrSksbJyf47GQHtnwuT4mbsZy2
LoeMWbXXyEgGDOy86rKPJ3OYx4wa5sXykm3l9oFM7xoted8wgSfToxgVtTyGvrrVZM9uJS33p2uH
jzTVgnqEsXmKqQvd7BhPKTZ00ZNfJsuI6E7RLz1Kn03MRtRHr5oZudjyxGJBWXZ5oE41tnP0sNGr
Jq5gxrDrPnaWTHpvorap+oDr/Vgo7nmhtLSMfWL4u9NbpP70rIO6JrwoYaLofuWsd1iqWD6gDQCt
9XJ97Pex8x0rKwpgHijIMPHo5MFinGgoA3pTL+Oa5yrA46x+eCyY8ds/vj8ju7tqbc9jgn2gHlu2
W5zSXtJLRA1qOHAXeOdLBoS8hPMVo4OQTHzc9OAEte6gmnwjwXsS8Uyq0i1hYsZs35SUT86c4p/n
mtb6R7RDlAdfrGyAyV9shJGcYlNpgAVJesUDj7U5yJrKjuw989+AYUaNsKjTXzX6D/j+3Ft8+NDR
ech5bWc2TshdKHwjzanvWf1hdED0PPKHftkKCSfB+s506PBY7ZNzrzdAq5BueMIqcBwcqnNxxFQP
4Ho/kfFlDLTsnIKZ6cGqd1QcKWGUSFyoxlYRt0yCRK+ZtEbT0ZYlu23AGy8U1LOf//3hIhP/ocu5
W66MLJdfe4i/1hjNRcrUj7m7Hsii9NHVxVCzlr1bZgK7lYkkyWUhIHBzPtjWCmw5PEPbe+3OrMT+
5vtaWLpp2Ew9eT67mwh9ItB6JXHp4CmopMGd6anTurtGfaQVs5sQV5ujONiqRjsEKQk3Npt+lmgx
K590lxNG6EVVeZWHtMXMiw/146M5XJZG7/U0sk9/a8vJ2bWG+bnM3hVRxagb6c9LKkV9G/WEPkUT
dSYYiT/9LO8dZ7G7vsMpYfJmscVF/Y8x0GaD6hZ2ibKxeywdBzy+isl2RdWrfe+nzeJbJxzXqqoE
V2pOZtFITmV6AJgj+LAYZp1G0bA/tHFHguILvefbMUJx4H4+C9MoHoYFWt1PtBS/jSoO0dj1xeZi
z5Sv6ffjzNHyBeUtx1oIH+nb3yIEppW4sA9uhFV24DBHSxdeuc44TEw1xe6I02lJlj06zlIEpGgh
NiHLEXU5M7rimAMB85TobaCSIPfO7d5w8zL/UCUCkaWvxWUEXjnjzKsvPaOYl5n0iRHcmZLqHKni
kiyJJEROJ26k8ENoIPKsUtXPzFOUCvTQ9hwuvjjQM7tMh7kUh3vCCxxxrd5htgFRWWRVQrB7sZQA
MVK2Mmrjhd/CyL+6m9GmCEDtoQgPo81aEOVRwMMV/Engyd3Pbexq7Cy4v+6m+7UshzNisnk3r4JA
mTSr6Q756KJXvBp+3tPRdQzFcvCRWRLDOV+vwnShaAsmcJKewYC4c2L7vxKxYaO91G51bW/RiOz6
cKNGmd8V0q4gWo7sD2Bb2txkGDt3CD+3vXWa5QgYNNs14y4QeEPgy32pfxyjGRMcHZPDOdYuX2Rl
p70c36mh01qwtG4lEykS8K3VNMT+m/hdD3eaC0E8jbM/CWe+5qrYEC/2Nvnkkhn7boBcgyzoNDxv
vynprDc2xlp/Dqe11JtmBITGl4ngMjjdyCqXsTXgOlrKtpM3QCiUUWtCdUv0Q34IvM4GwECf65Ru
ABEksz1Q2xpKTUk9TjvsTvB55NSmoQHCKBAw+vYZI7CA0ZjxfkYchAmy+l7GVXei5vuj20NnLhjI
8B54ahaBf/IP2PJsRhjW+yvGYx07XpX7OVMZ59bol+devlsVQP3hMpYfx80JcOopd2ZJiDOQaLdM
VUVRXtGeRd//3GM06jjKYajAXDNDc3i4IWHG0I2BUVHAYBliX8Fg8iP9Wbvu03JRtYF8Kx0h6SQS
DxshQxLJSaGIfLKu23qGKnD3yU3Yjju5yvORRw8yhHCLB8PMJH3gQVt85l+LwuPbXgWgVKdhOAZv
F5LUO52RlkiP3wh8ZdifNs84SwckitCuFwdVp9q5rC/VDM4P3bwj121Ug39FRbG5+FkqN7PWQVyR
jDofFB0JAaVsiuM7GZ3eox4y/rbuXM8jIFQaXEdj7YVb3Otr+9NFMPJUODfyeHfwp+Cj6ekRB940
Ffgd/bVlejVRtdhjrxce6upk4QkfMBTqoCh3MAMVr+ltAd0TrIdoViZ0/zoPPk2r8PXN9ZW61CxB
wqJrau56kRUIzZ2eax0ngS+Ws0ExtBjTDLMIG9QKyqAdlA8Dxa+37V6Kw+St2nimU0/bBhHdVLIh
oktexTLam1aalIAWynxUY+xd+wl8nWGxYt/OD5+B3U3UeE1NbTIghD/QL9gq6iNuQw5znIylCw4t
xo3nZ3y5qNpzmJxVDWehsJXGk6uhzHYBvqmCdM98AyXMJ7eQyKEQvGp2wV/jCj6SKg8Fxjmm77Pn
695U66BtAksy25suy01bDaz0fZ2xrJDA94feHMjsG64Gv5NGpUI1rkqzh0/ocMdq4BXN64MMDI/G
NlOhYEslMlS8n2slQ6mvSYQSJ72l2Q9wJIWwYihkT8JlfBxnLESCsrvbzUEESfZQcFhFd4orM9Jy
u4BuJgHVEkSggf9HL+lpm6fpZANC27I7zl9AFcc5Vrvwk2BxQh8z+VLjiURHfmFMqKUaAd227Zpm
OZ2B82Owy07NMLfZbj6kP1eHXcoOlN41lOSG9IjTfaGlGKKrywW3SPBOjljDXSUw50HPyci0Gm5l
XkWbV4jYRoZRLRL9IeoUjw3CAiasp4PbJG/GoBUeN927v0bjfk6f4+qZw5+W/IjLGQbbZXM5Isdj
wuD0kUpb99bY5VMuVXpfp+e1x83Xf20rWwNJZMkx2I5nTWMgPXjY7/C2IUBLmRZmeK60qWV/m1dq
p6oLwtmST6iaPIk7gU1Jy635YaAaHIVsq0H4q2GKnBmBUPKgVmJ1AWs2MYs4OBlhUZ/QU6adSpYh
VRY6Q2UVE/vjz71Fzxf4cvZL4Vjm4oydNoI0VpE1SeTn+27HDszzYy/WvUGO+tvQq1yg6WXL6ROv
kokefrA3kPKhuTFjrtYPM1+M2WAD0nPNwwbljdDcG0pecJEecIx6qvX/bSzAQ6qqLds8aD7kcAg7
0PEKFusSmEOClrRbmt7yTISUcpAKWyP7V7YOOCUJcoDpdXh3ByYbSdeeoKo6mLD+3X4Q33AEfS0u
oOxjPDFldva+0w7+MAzxPD0WxzHfBldExgFW2XB2Q6kIG1LAzK08gWGxn13QHhb4pXK8rfBpIXcg
twelGBrHsAsZx4pcGVIHpzHWxarB+beWgfsSc+f9gfor0BciZvMOq//P4CjxgltMYx2iQsQv5R6A
bp95OJQdtKIJV2EGnloslG6bf24iomdboXYulJX95tsUlAFKoFQE8noy1izGXFSw71wPv0pCjGrV
IeA3chongzj6MyLh787Ltmnm7bEsavKOIctGNvM2t57qwh6iU+bKpVw2KN6KYVhNB2lvos7kc7Kr
bi2p0UrS6whPseITW/tOi5b/+tIwUyBxTcAkVDntmRIsrwoduPo0AS2L/OelkYjFlFoO+6WxZmEn
Y4C6w1LVdmDcLD7dunmJUoKra/Pa8ubi9lEKiIbqaySpJa8/jF/Iw67VYPg277sHdMqCNClv2psd
QC/CjF1Zbo+QLGperG2AtZBK8Xn4U5dMKnjB561pXBtecU8DTQpniEoGV0g/+515jDGsefUVkcHh
ohenu7kcGm2poeQbHTQKRveLZXldPS+YiX8mY0f1ycwgw43Pc+1K+KCbQPkvDu+bwREL5xTNfu9F
cPzJk5eXJ4lmmJAeFvPy1TDvIGU7gRYGAS5oFWo1AzlYndjaP3pc3Cpj4GJvsp5OsgtcowNlQHMU
8vF9AgEW+Hcd876j6hkNXCimH8AirCjdZHmbk4pgvDz+GU9+9r16BZ+dZgKFcRzVCQhEB/kSI78J
5xDOaDFOGY6iCscngKIeCAeJ/cFFfFWaW7KuDr6CXp+4NapA6R8bIwsnWa9MqJRj2b3UvrjnxT93
C3hnHXekNB4hPxzqO4/BKNLBE3rJEWYfFCzqqO4rxEdqr7dXiT+19444fHzCpZIW4no3wbah51t4
AfW/JlWypQS8aEZo/i5Uoy6xRmzLWSUXyCGXNpj43osS+04Psc1NwF9wEDG6VayLcMOwgfi5dkS4
ZT/WtL5YqcoElKO5T1PLIG2+s5trwrl3kuQR5V3MgbhqAp08jWxtZrnTjXv5dnjCPXUl5VGir7fH
k/AeZ3eBW9Qm8P+h8H/zps+vhJrN+I3r/EZWm64ItDSlezPNd+4mKfg3QxVha5w+nT/BLnXSt0Nq
xwKnJg8DE3SyGpvkwhCfISY0zFebalJxp2JQZ7Z66Ho2DxqnnRHCx43lFjePWSrF52cB+YoQ9hqd
piq1TQO3vBQdjejSfwVGXfpT0+om9dQTwx24JStvK2ZgPljcHWJCUAZ7WNFQjlNxsK/z7EfnD3n9
hEypCsNae/mXwzMBNucIw7ZefE+bT+6JGjehHxvkCAfc5onCXQskeYqTTASkAzwlZd+Dh0Hose46
IInhxy2NN3VUAiW7m8cwpLHkao2MnR3f1MBngqHKXab8SdK7j2/pS3aJ6jCyCTyiGIxJkYYe1VXd
djcqFVgwlbCRJjSw6I7AThhcCnsDtj50PJKxxfFh7g8C0238wo6Z7/vQK54plKwjhsCOHJSgdWmd
yQz+7WGt/jZpxYuPN3bkxdBZgbwhRNuI+XNXjzjENmjCxHi49t/BADwv+9E3a5w09mSA2m1D8XG5
S0ZhchiTxoiDWJoVxAjEBND3Lu3qWwHxodow34Q/lGn9NSbN3sbnhgHq3A2kzqV0OxSkhlp5UwWz
5r0KCxxZEnL2Yn+hmAxaZPniVnl3D6EJVOKdE0ATQgt0rjrlX40REaMGeRdLtrxCqzUUL/2YJHJg
5YoIgeBOuw4SCkLp6//7m+DcZnDdoqmEZZwE8ItFwiv+lpnU+hC5LfqFmAvAozIr47tnKXMvh9gD
QD/FxwpEYPwMBHBhuptVGUuUqj69q1t+NF8zC/GEQd76jw2wCXPxjl/yvuzZWCrK7y9Z1Z4yNHMC
wEp/Gk+GQdco5uwWKEa83kjp9OJGVEEO4Qz5b5Wv18VQMPtphZxksFB9AzYNEvOuBugL3lYE0hYI
M79ZNmMYtMXlhgOatrcxwnzOC0KwWaFwgIT+LRKRgVWaFo21+hfpkfqC5n8f73XvNOSPcVl7lwGI
1jN/P0YFMxm/6FvhfuCd6ExOlWSO87aKkv7pcFVAp7XDD+O0Xm0qWNgrQNjeXH3qRN3tSHdRzV3D
6FU7BPcd84ksMAsrvD29famMGh3OwcZ25IA0xWLl8XjjzAbvxBGLmvEGW0Mq7n02MQRSAwc0+2mx
7xjOk+O8ONMKIXdfYQbY4dwnwPojBzuRHl0jkDhy3pVr5ylnItoVe8oM0fwX67yhbAoXwym3jzu1
AxvCtpbnMD+tl1ioJswFyak6P0oQY6v9ujQSdiNWXzhZuqwborcM0X+kILBohfDbB0YHq0wPH9Cb
ZvmAGp/7OpKAmgSP0gzLHGBZNOZ5Ck8NMgvROxY8++lcLi2aLXRJg3JC3TMZfZtiSUuNXnMVUvJr
q+omoIqIi5RzktyAeGIISkHbRw79QCJVF4FG0ITWcFDv+nEQffDnFwlDF48jHFdNCH7dZpxoXXSG
krM9LAFs7JJdy0nMoKLoiWxrCH7rjlLdGMEolr/ScHOZaz2KlKJZ3lip+6pi8AqWx6q8FgsNn4GV
4OehsJCRrMuoKaqez+6N5DXtbNA5bYvuuI5yFt+nO3Kpgm2aSrZu5j7V/RFX2yp6+6N30kaxS0kb
6WgPZohuILzVdb8ghjeGzml3427tLMAvTewf5nBWyuVF/MmloFGcvYJu3/2Cv9ywRl51uqNtwD4T
j6Mb7AH6sssZ7MkX9ytdXsrc7W8D6mBR1VD3D7YtJwbnGjhzaRAR8YmRrZbxlct6nQGwAdsi+sdT
YMrfzl/Oyd1PEvD8U9NAeOBKMvZjYqQ/PkFFuAtnMQ/oMRps+PJTtnqpS2CLj9HiFRqzQYLnOOCS
8M4Wu6OgfW6R0nnIdCPvIDtJo+MmIPHtJjkj1p1HTUmtd5QcbBfTWJW5EEF4qC81MKyYDrtfN3h+
OBt/k9E3KC/2IN3J6jDNwAmgbUzN2mSyTuCbT4ZYHQvEvkuOHsj/Y86MdR+79r+evLb/1cMTobjf
2BJVjqrMenPIfk0AqukNrB7je/cyWZuaj9WHgFMg/czRvdIi32CcElkL9Gstvu9a3y3sD7DG9vP6
0LuusCY2TwDbAabsiWzMJ0CdNAQQ64huG691qIiRCDekk82tFqXVGpHSl3jZxERssuOSzuD5K+ja
qk3kXI5+bdiL9tL+0O9pKPHXGp8hWlfNjMyRicyevOONIyk4xdENaT44h84xw8qa5Rt3jjhwMume
eQu/vElUO/15eYz4+ggqrB8sNZHj8Vbmr9jBuW9dwHjCSoAit+DULxhiY0uOBssHLBQgSyJnYZcs
+pbGdRc+7lbmsj/PszW++irrO+6TOBc38gNIjeFl4EgjWdexQBpv3X77igT1hUcWwpjn9YFLgX/c
4NzuDI5animqfKSAre2u0RPEHhSP9ZkznGk7/XD5PiEAC2B9ywqwWZye4GNNzzZkpskHS2ZNDish
4PAJEoKFM28PpmhVXqyOeeWwlHl1kFNKgzVTtZ4gHHmQApB92ULIJN6XYEmY7VjLwjwm31xEq4Uz
xzFWsHg4alK9yfDe3N4j1U0sTwThdoe155bh4U6Q7/Ce92dil2Sxt4KuQNiWYxnuUsbHw/HG7cgu
Tra7pQLMluLT4eyRO4EDPmVkl/EX2gaAGduWJ2+2HNnJZwzGF2B5IVQ9zG6Qv352ln0NUOZ+R3wI
X/DrWh+aYA0kuZGgsAMtf6s8FNi854612VvidBq+fgutyyStrLGAvus3oWhg6AuKxS6GZrDqiXDB
G6T6Y9pxxfTQ/4fUbV+Jv98pjOP5Ev9GZrkgCZoVXjOUl+xQmkrRONb1KYTF5t1II5+b6LDM9K66
+dIVi7CCh6zcuMNk7Witu0uoQxZ+iyWGydywpuyvsZBy91pcX7XGPEIHYYeD5TLHNLi7uZkBXhaZ
V20Y72drq8yiSEar5Q0LVzvXUsHsK3s2bLDbVc5PDIlrTjBb6DZRYNoJgAFm9IRVrCmF4K9y/Sw1
rPoPeg13r5w9rGaYLKSiSc+FowblRicbmjzy98872b6UMSx3b/u2wu3MN08SUUEsm0bmTBvB/WT9
0ldWcr4IZOhgcViNaF2LBnQw7RshYJA5F4g+Um7gZf6iNkIEjWTF1lEWdoe8homAUF8JLXidd7c9
vd0PXAH+2ZXRAYjTzhZQbSZy+xO74hmPYO87KoykEhqO53dOdezP0V7Qyg8xpnt9lhW7aVP5nqEU
rriEN3d84IzYFlfMe4sfqcytZ6dM7aQQU0HZ7rzCHdw30pXu1/bnYpsNEq9VKLEnl/qTp38P39Zg
FbLLi0ga2KQuUP51BzQfdUTpMkezcmy5+/QPgWiFllXtyPVySj6OSCWNZ2RomP+9kzdtD/X1K3AF
JeH9HHRwXTF4k9qoD7zSbQA8NkLo1tIQnoJwXRKQaDNK0sahNRhQou5CNCcYePvnM47KtBvHmTYw
OMJA/SXyfBourQrJDRHVgUhPXEdW4dteShGilTo+VppBmiCVYozXFoCRe9mn9Ih/tvdGiemNofo9
4+HB8p/2XffbchJshPEk+wsdBDt/ygllAerfXFIWC4ggXZM/sXKVqpb0rPJEgi4EvacTJcnw0FJJ
Drohb2P5nKmrbu9YGU0Rb84/hsL2lKvV1iAV98TnlYu4N/3iR2s5IwiRXZKKElAlb+47BCpB/e8t
DLWjFEogJE/SUV6lWIdbRPcvI/T3y6W1+zrGCHPyHG1s63FL+KYsNVE7NJlv0VLerp9l+TwpObHH
WC0sE5FIyafRLY+hCNEZqvinZ5qJITovD2kJZIcku0ESz4vP1jHwXeHS/d3CfMU18nHzQ8EyUqMS
fKn5OYnWnKvZPWvEQmNzwlgVM2X+rlXTyYY06kyoTevH9y+A6Dh++KULf5NuDC7QlOKvRW2wApmU
whq7TMRFCVxrQdXX9oXG4+NT4FzJsFQj2Lcht1IHhuO2pqJ+ga7m8GWnR1wfhegKhotj7aSQyTgb
xzyzwBLE7yJXHp+lu0iesnVrPSdSCjgwA0hvguHy4i+vWs2symdowtAYwjrj8oq20ezGmDBDwnMu
8H9TUUvaB4yT1hz5EcNE9u7NP5gNRgQe8kq2pUNizj2U9b9F338IafLweEm2FaBuU7YvcWxnpuv6
EBOf64SGgpzKbiOXHt/2gYF9prduFdOXaXWSW5FeCjExI6G48t4DvE9cwY85/QRwz9b60DduIY8C
a8WNDQnCYEUrXDRqOsgJTLEwAVSAFOOEHM5FVqt7bkNsA8x9nyuaDEVN2BiNWmR2UB1Bpj8ACeti
c/NrL66pFQTioewweuTcXCnsqt0vO656rs5TDV4Bs2ZwKPr3+3pSAY1o/F8HuTI6m8J1/+0cOStJ
hD5qB1E2iDebvPw/EdDJk82vQF4RYIdpxxo43283j3ZgTJ35Ez4dobdnsZsBjl83F9n4v3vvbdeG
Clfv+4SwyVd6inxP5IV+Sx2zEVurso8bLTPdCG6NF41tq/tjlyiiqOhpX2kxOcICSfpBqroDz4on
XUsEsvwTfOAkV2m5JsXEPCUh1xYrrIqAnqosK1uG/7Q8A8DNabkka6qybMB4Q179+VQUGlaHydzd
3a08ES56jWjmyyMvmr+nFyYEZGcxdu3PCeD2CO0Tf3pb89L/RFeahmvV/iyrCPk+AjG5/wPl8hge
C6+jk5xgWmXqP1hhDt0jUexp2O83wDRdzp7s35HKWPmJqXFF0tGWFOB500IrU7bLBjq4euLOW6hR
uvSO2LiAQyk+DNeXE7L4+hmjnBmgRE6DZG5DpCsMud8zqZHLVvbYTyEG5bl/ixJTIWamY7OTGloi
e9YnOnGCmNlyr5gu4prncQIFMueuiDuYgMCz9vImR0GdQdmBkj6KZn1KBv+7s4+NwVItjDcav7GU
ugxjMB6SGydx3HW/FzcHmlz3Zv6ibQXtaNYSRA/D/hhppcD0U8h6qKTjiyr5NyQI94D71ndyffg8
+7t4b5KmRXjQ0vYT5DUHOGOWhOW0hDp5og3RvPyPCeAOldNJ6vfBuea5GENTq1Sh3dIgNL6fjEDW
mJYKLbqNlyprH1u1aWDSDVjNrUrNPwwWdcvI01F+il4y01MGZ3i78vaJfqKRvNcCMvxAxvvMHwSe
NxhiPaZ8z3cHULFAD1qx4pazHyeewGCWQvW91dXOUa2R6fi3vwZUAspyTRlqDjtMHDip1Cnh+b1t
KqVrMtiYkgodIE2NRS+2xay0bgyu6HlIvpNXG8J3hp+ihK6lCq7bKpydDX0XdJuwqalZLwrQqUfx
rcMIt7T6s4yZJBk14XuBHjn8D2GJvYHM6iCI5lCs/CkZLG9lAYXh4MDHZXkBtx09HqP877p8TSco
rIxkBk6RDfygoRgx5hqY7pisT9REBjV6gcD7Gu0dRNX8UiozIdFrj7ySZydfwbx/pK3ydESZzm5l
Vh9uYPnx0zfTYNIKBLt/pE2/k40lo45Gpy78aI8FyjVCr8oUEbvjfJIcVKGz6/Q+B4B83hoPfBwz
zWsH5y6k+7AVB0i2w8AtnyuNa6XtTUyjuIbnk3GisGRU8efEVPF3lBZI29Uqlfra687qDpv9wILF
Xul7dwJclhlqokHiPk8b8Pulfmq6l7Ums47i8RatLT2nzGgCUDf3JVue7F9Qy5I9nejZI7PMY/LB
MnOiU79s5Fc4lk+m8AMu66s+CHHPyudhkr2C8PGYSDfI1lTqOzjDU4zC22pTlXr6A/z8dO6RSj66
aM4tUBkCnkluDCLmn04b1atMv9QIkbwZeg826WwUtt0k7ZYV2R7XbHDLQxABh1btQfOqzSGtWuyz
FaweMkB9y+npXctRpl0OnpGzTRNlnsSPkhqCofApeeEScM3uhi0xsfRtzdoMPSi5U/VUlyTGP1gZ
HhC3Vm2ppGdYYf3d5T9JlU+E0mGyi0UVfqsebSVPuXut+BmDIp/sdJWjpyol71POvaD0CpUay/Dq
63MAXOJmRgFmf8TKaT0V5KZM12vcWM2E3bNst7kkG/wbUGqXH+psC5UnAM8eYFb93a2yT1GUWBmY
1cIYW4KZOUI+Lp/U8kmUCTPqRzynNCy+ciJbip+9DclqlmdvUJ2tK6+RW1kxCHu0gjhvFD4xdUD4
3LXjoFU5FfBpD/Ea/WaOKWWyd28e06s1iRC+EDARecEjeThyfoQsFBEzxFcM6k1IZPNtomRnJKwe
dIg7upZ3MdV1TuArwMKu9ooDmT1RiUnEFhOlUuDKTTDEMmE1ml23e9d0QUnhExublDoqKyoiHj04
Bj+xRR2loQDCALUA2wNVdmH9/Nea6TFzhh2sQcR+sOcDHATwV6yF5yRaAIgFzKl++mLQwXeGwXb7
LJ0fnfh+o9nwWzuJfT3wFH4uVrr8wwN7Eu4sviy4Y7nX5X+05ZdYH8ZI0e3AjchxYbFt2dzIEcpe
2F5Dgid25Rdu77FgK1e+AioSfSBvC4XxLwXMjpPujDMloStKIvq/uUGCqBBTMLfkA+BK2KJ0Ytsb
NNuP3QsJFfA9vHVmXX2Hiv+wlCup3YVbmXS/bOkjl9W/Ly3V0yRWu9bXwIK5OYRraXJMD/fGohfC
icMA72I6fUqyOlSErqbUbBefq1FI0DA1Mejv74os7vQivsXPA4fYO0o+FBeYVMeBRs0npakBMjeC
CVOVkE7kittMWI1TGR1KDVWI6PEcUWT20Nw3soty8u2XCLqD1YHtLrGIssUTUexyn53GXaBgu85k
hoC1lO02/le7TUmEnhvz7JWWsKz9XTNA0oqtCI1Dt7BEiLK9Fw9hy6MM7lY+yBiEp2orqjxVy+Yb
5QolG2mqKuIbrvx+p10YZsC/s3MLcTFfU76/8LjR12iJtJHUASB46hmQCYb2tJW2LLy+puCd6j9J
dGeG39S4nfeiMZz6yS84n1DSAebnh35FrEzaJOfGA6iGfgP+MNaV0iz47GSNExhw6Dol4NS0JbWR
NHT7eePMe14mpWP6f1X8GpFXX3f9WOYxfMneaXS+4p/y2wp8lA65Y95HIct3vFNdSGvD6qRMtqWn
YkoBZvOo8V2uAox3KiwUglCzeyDTn20uX5HdeAbZ/nCNviO8ZRmYhxcAdwlUS6pcePiD/GWhye8M
bbIjiqERaoVwi40bsXECqEe+YvGU7ndSIvzxDxRYUf7IL+uReeAI+MoT9LrM3Un6nFhGcz5mnf+K
5DjMujCKWE3aI0EVintqEddv4QGX6cb/nmv2nFd8OFQ9hEzaETu78n0Mu7EEheIZMgx0Lewg5y0/
GfDCkWSew+t8TX2QyP4HAIG14OmQgkBptzo4j/Ze+Alwd6WjpdiQWSNWxzYO7EqOEExXkEh/xFtA
UZ8zjxENvVpuOs5qxoTKlb/+o+//QqTL4oANO6XtjC9hpBmS/0FOvwgpuv9LKtKrwx5NAJl/JZtb
bMUUpZ0SpYkaw1hJmLmqKVRuplLrouO8OeUIBXc/uK050BQnLSXQvoBv4wuYC/0vwasXzu55ZYJf
y+IORHsq6k0srjRlKPxqNo9bhmhGlJG/AXltvCtrddLgkWFcJp9TtHNxXF6mXH7FUbmzeGGWpzv4
wUP1SP21cHuO4eXYhbvaBwFS0B5wF8Ae6g37VPWWYEQ3bCffX17gFMKZqA+J9gspdsJnkCiCaMVF
1YteCiVfIygs2vxkdBaCnPJ/yjoUbvjjvWEo9aBT/IN/Qek+bkB9AYlezsZVi4enXLBUCFuHFY//
dLOu4RBOAMrZ7ZrN8hKQUdNZE8im2+7It5JbfnPq3niBxWDUNnYRADNzxLodDTBJO98PLsu2rZo6
tXC+Mlk3bkCGk/Q/nmXJJlfngQziTdHDyJxijJtaUwzCRW2pUcds6o+aZVNZu3x1+ZPP/ydcBEGb
A6hZHoeenb4DLRiXxluZxMgf2Xy3CVag99Vu0flhMJYBsYFHOH7RP6iyyDXTJEB8SqcBRXlsiqwA
ny74ZKx10gFVzh7OAkoKVCCdC6ujSyaHOGM458HLreXqMBx5dwUJ3iW+BMVrudBfNzErTCZ4xRuv
/8yqFfaYiYjrvRlM4GxJvQkekEsUl4c8kUxCO8xDVK7qfau8hjiwIbo/kxSt3rANMgZgyO1YbaNZ
3F+poCqClK4eZosWM71Pd21LgaMceP0J1FFsrIBDgXUywLDlQn8TSb+jfZyHhg1wtG1AA3jfOHcy
wdtsmzDrpKDegY7j6N/tHDxP9nMcUr0GrzKHqNSi72YDU1m8K/aXD0535YpY6JfPii3CefDoNohk
NG8/ulbaeO/Mrxx3UuNjtHdfsMkpmKnNWItcfe36AT6SwBA9LH4D18BCwiLkkvqJUuibihvdsUYQ
n+Q1HZYuPicF3dPEWoASO2gNmUA5FGUn/mSLLnklxtRTxRLZG8YNPijXjA6hPB+iVttiOcOjh9uh
bHvSZX3jPmFmWGbH3uqFSN+fJZHLB72RHbo8b301znQsCy4a4coprpw4YqOoixnh/u+uLwHoazWU
wO3J+d049efoWhb6PRANaLjsP05cvSniJX0T4OODfGWbJ2NvyKhe5m1MthHs9v4SAtGxEJI2w0D9
kHyWZEEFACstAJdxvB/1VoEFzxvv6f7QnOILMYtquLtC01Ox07dU3d+aB9ToOLiVsPwefsnjytvv
WjpJx4N+hKU+nm8D9w50qhcr4enyw1tMN8Z7/ap1tgB+HCauMymOxTJXuJcQ9fUIYmCdCGvzMTfQ
vYWm11r3GgWocakCl9AFCCqAKTD1TxMjjjQR1+ZxCAisBhejdeYLM7krDaHFBW5AodkFLyKkDlgY
4ZCZUMlQSZt3I/o1RWk5UMYY3MaHmvBlUj/V1MnpxLzLoZluM064oBjKZ04GYBphlmggm3p39jO8
Z6jpWnIGFdUsbDtS/k7pT3Xsbrv95MxPK2bI3W3rrvLQQDFLCXjho6z8/shG4BJzZmJlIxS0DJX6
0Gr3w5dHbkcjQSmvNeUo6RVwLZgT2Y0dxJVkDBBu7nDKjQ/M9XB6rUTAqhMVIAfC53Ouc3ZWnP+3
us1mAozLosyDvzzPY1u5KxM/XygEucSlBdaeec21qy0KpNmQRkpj3go+su2Poxe6AfLB+bTCTZw1
7WI98mWIVF477R1Ug6fY6jl4VF+g2wPjEASondBDwyFbMaf0FYxzUrfn8N2RIxip3oKNSmmsW1ki
Q5v8K1MEEed1hXJEybzUMtOl6mDAtzmi8dLcNmDlGkaDH762HSo0KvgaWzZgHWBlaHIeu5208Qpt
KyQX/kMftOSSPPQrRi+WuodsostjFc52jb78i6BsoDRVh4yGYNsfAV/+5SKR14bWBJZBIa2ehWmZ
Kl5OnK1Xh2aWkiJalCtAc4HUuQF90o3xzRPXrMIj6xfSkkkzyrwykcF/ytHDnc8TgdAQE4dtsmDL
nYeperZRd26aBJfh9dgckBAC9WhvxzQ162YSAHTiu9i6DxHhg9htD2oqceAV7buoMvT/Bb+mi/1W
ytvPtxunWEi6kLixOcTjFoRZh66SU5hIlc7brC7pPNptwgLyaJvy/spHD3qhwYE7jQL8VYpAc4p4
ratH4X8Cjj4ZjecDHaqxa7UZArzHXRsbhoRFjJoHQwHKQ+d5RcRhYd4/g0Skg5AorxTeDoeAVAxZ
82mn1fAwTHh/fufYGEKVfweBvb9GdWf+QcYmaKsU4olJkwUX8A+LdFUJp43kP0QoQrqztqZxxXws
oFe737a9WRQ6KVTuPgmnMm+YsGzJY6ebbsonh7GuDup71i9NTc+gpU/2Hg7EUnPaV8/BOo7pJj2M
ci2ju40XX3cLB9iz5kU6AszWjmpkAzcHbo1ntz2xG5Pk0duZMBi1+AbUjRrNSZwy2fKQ7893d5w5
AYO9ZTYv6UMWYReWDEXGyfI+6oK+9yvqvwLdQEP7iwrR6MopRcMHlmH14p7JoVasS7IPyLeM4WIy
Yf/BldVQOlFnvZX6ia6OqELbCdEfqgTLaXvnhWjUUvTt7pbcX1D0fp1i/MVRX2XEbh2Fo+ToVayW
4ud8bn2cHA/z3N054zDjhWQ34cE0XWbL7UlKAmg0eCc5BbtcOQWpq/dCaXo0747tEUoWCBfVDSOy
aJYOV8H03ssCSPP9CGw1V5IDn2IEXswoWvgjQdwEXb8aW+vA+azGYBGmGmU392zLLc+SqBwtwGhI
3ezdx4C33h6dVN0TTYi9THw7lAC9RCO7Dwzm/nDJBfHWAq/uvulAAzmeJOukl/PCVP09ZuHSmbbI
eB2yesAz+rcdtV2pNGeseDKub0dg6Vsc/pKuOJRo3/QbQtzCVYpsaYJu9HjtfB6vVL2M/QtdMsPB
cHMgq3pFw60bs/tmTBlu0GMS/G/E7SOVjHhSW9NH4cekbrQXyWpiWItXIlsSV8zyLadTiP71sRug
4+BPC+0Qk5CbvMtPPREr8sMwfkoPMM4NXkYr93HpbXJCIj/yh0lIBZ/Rz4kVRNqTQG9KS8s3BxT2
zvr1I+KuF/scAa1TZHG2EDlDs3588lqQM1Z0Q3h8H54UHdOZQ0iB0eXsdC+Bm3aiu28vGVQlPuM/
ehy7EnYlB0+XXFi1otEOw0/Qv3gxgJ6v6GDgpNcopwiZ82IHosJMgjz7HdWFWFQer01HSw3d/jJ9
Tnljkg/JsrMiouwS7k8E0S1AmqI2mCWqRegMTCjyZpsCqGnywJ5TUzPjQfRxyhKtNSemHG5IQ/N7
82KKOLEQDB3bUq/upY9GKzM7QXl/MSBE/0MqOHuDhYFUskOujGZIIyeeqgziSqAAiWS+xxtFjmB0
9TRlqo9ZxNn8XRFfCNga4V9alpWM54KhArBN6tTfkWpg+LuIsahImErFC4ML8C+NvZrv4so8ZjPL
KGWJUkKfB79PayjQ2hXKEyB23t5gpiVkYnKF1P+pDwcVPtpKh9fFlSn8SiNftJCHHSHnC1/9e4B1
ck5qeug2W+UYHP13zfzjZlWiDCI4w2gJuAdxQNefy1jxvFdU6Y0TDul2X3enMuzhcdDqZG5dhKPo
vyTYjYbDrYCVkkKBJ1hJNK2J7Zjo4iGiEpuRSjfXFSzXnGuYwmGYQtbYRalWI5GL4eAl+xpvk1Tw
eK4lNPaGdVyAkNOAhY2JVM9L7/0msDfWyGX+9/DkqTvVcLgsIke8wsr4thA6crrrfHnIn94DJBqE
HY2cT3MN4cPBu++vn+gCj4oWldlXXdbngwAsHwysZ3lF3W43eXJfxLqe0WVfMBqGz4vtvYQrg+bT
SxGu/ICijDtzHLp/GO0Awx68WM6bKWu+hNQPPAb+ADCK1XXDpSIllAbokrh+sDagcbljLH7SWMcR
l9IvGo186lrAXMFK0FSyANOwwGsnnXJ4vbfNhwymhJ/FZW9qoXWI50mWhq6XOfiUrglvlpyLpJ3Z
58X/stanctXKAGxX8KvPWP1rqBIK5+DzohDOTLOI5HYAjm1WWf0Dj670YGreA9B/fmtlGmXlD8pq
439EdpmnrgZvmdLqV4cuBZvz9AN7YqdtSe/rFIGU/RSDz5CQHrZhYDqEwNM6rK3MSy4suRQVN8vo
O1f09lMKvJbyfQ7yHiNNUb/lxrsukOiYJJ5gL+9Kftq8nOZWGGjXgz4LHfoJzr0dOt0vXOAajXyE
yQVlnN/SmdiRt97YJZJjENlt4jEDxyxLLya/fqbAkEqm49da59lAMzthCXGFLDBLoQo7qW3txi9d
gKEMrxg+ohdjxEmfGWQc4ZHlNC1Q1m5ylCo54W8uQIdTW0HM6BhMz3x9RAOq2WqdyRPailU5XWrV
g6btKevEsHwWnubmhqlR7Qpvh/TFqBhzo9kRfSmmNcTUzC06pC6jvtS38ykpKJsBUni2Aw8hQd2q
KYz644VFgh0jJJ19h9xT8FyvHZuCDV98lj35CVH9yDRcJhqytjenOi5n14BVgwA+AlyMKCGZ0Qy/
MKsQ+dWtauwJhLQKZrjZb0D7v5tuyhaW9AaUbEpiNaGHjPEMCTrOk8mET6DeobU67mg90vNIsplO
4jcPoUnJ6a0nvDnGCGenVmL59SmrT+TgjvejlEIxHbIrqu3zDzORPoFb9DTCOUbnl8hgyeWYspbt
TrHHZuu/zS0WTN7TYBqgYCxMpTaHAItXnLc5Rlhtcd5ufg8WQojXrMoZqT5cG3ruSR4rIZJ6mwJ7
J0Uqs1En/wvvoplyuPbVte/uSRg0ucYoUPQ1o6JJJUNVUAN5QkEpDFjjEUXB9XTLGjAfYlQ6PlC6
AC2An4BbRgLg2WCdpO6oW8RGHvVCyiw0jJPVtE7nNSYqua6ARMSzqHbaDZqHbnvxvxqLhlrUj+Zj
dh0mohejWrl4Lw2JiFG1YUFSmr2FBrGUsAwwQkCz2qWt8rQc2wRmQPtdqeSC+f5q/+zjlStObAEl
C+fODtEc9dkBSqXacweQX4Qhd9bEKIukvnEsAdXrrrheKnuFQKBEdcsI70DkDGwAdjTfAaTRBlnf
dig2//XNUUqlXicDdEQaiszh8FZQ5LJKq9zq5l031Mtw/voyXSLwE2CD4Ht/uDEqhr+G/0V06Nsk
s9jqy00T9DZdB0HmwJ+Z/3Qfx2NVoYTXQRJ+NYbeKX9MqsJpWfKnGiTfaBWy0WHTc5yTC23rsHJ4
UD19s9WLIAWJxN1UjZKFLRQGauSzzgiwa821VYHYN9JAzi9V5p72QCVQ6ZiCqRKRztShckiZtPKR
vdJwWfuPnUMpW0yUz1PBnyQ3VAfY98Gd1KPXgwoF2Xl+VWqTTUXkpX/0xEV6bhGUgFgsFO8rMmOx
sa74HdCVpQpsvT2H/7Msy1gRxP71wQYdqh7JDWn5Gr7wGvU0vrZ6KnyFAfLHy5VJ0YUJ11mOTzvp
flFbYCqYwWtJkM7NomtXGyV0XO4mThj78SxM/eMz0EpCPRyVrW30WOlWUMD3qsPaOZRbjfRO4E0/
hQxHk/TprpeUKYEQzJegBoMYWs8jlPXMRNedi/Mq0uEe+VrlVo+LJJ53ae0Ukv9SceF7uqMu+GTV
G8I9Y1O2CPtE0s4NzgxhR934gf7MCpBRuv297fS1AHzyJ271qf/PvxSUax3wtto9MLfnhShhveLd
Y5iiwZ5cqqU6ZMdIuMvoRuGLbHZhGw96AuOfoRJH7ECJcnv+oPBQEOOX2zNhGKoYDCcdd/ZFP3VD
ISyRQsiiqFCQxkCR4SXdZ2LSQv+gpfW+nBCKOyYkH9RNjnY2E3OtivI6DCnkgnZIyUzwJPZ2yTPl
7oWPmVvCtMXPVNzmdeZk5rdOwwzTjWeb3+i3Yahe6F+99s5lKF+vi+pmQQmMovw36QL0Y/Otd5HD
lTh/FiEI+yDgUvQq2Vq1PTD8CmoW3/mqmx7oBce0basQI7cMp3BYa7Tv81aa/jMuD5J7r5nve4jA
etRfcC8YP0kwUaqfzxIXF57xYMkplPwcNoPC8UdA4D9/SkD9e5CodyV/FtwaQz70IHHqtWpi7ZKQ
WOx9OumEHYnmfYdv5gO37Q08xSUng242wDprfp7FQ+VK12deiOxOtmaJhocCqhy4D0XbsFTHy/s6
ANqCl+jvzX7AxoKLydYX6F6cwOWGdLNkYcNmjIAtDMzwfABNeKYSeB7PwxRiSe21VWRx96K3lktM
4bEfVBcjtBDvzZDxvfgrwe94A/1Nc9YH0ANj1M1XYuGGDnIscthXZYIEj2tsbZjVvu8Bn4bsKKx+
XNvqi/BLwI+HkH22X1vxuyVGjcsbGJ6TAUCfdxeOuqMv5ZGSmFg9N8rm2uydDCwMKj2kZLf0sp9D
QoVmex1Nzo9+ncD1vB3qMGmQ0Cz3bbBYxAsX77N2iK5NsLNuvc92hye8Alku3ZFhsCuiKmbteb7y
44+8jzq1x+O6O9Y/avFvb44KPr/hYjbDlkikowGiMO8qeLuGaVn9P/vL3rJztL1aeFhhx+2zwnCX
2u9XtcLgoAeagN4hK+RmBc5TBPJRWz0NDgW1QAhoQAQ1MbqoFWZu32KMetvVWbt7tFsfeAqw8QsH
+3N31qizKLoEzipmu/4+4x7xwy8sKDiNB1HgJsRPZSRKX9WVArKwPOR3PqPfsjRZgGzsF+TitsIi
aS11UEOeAyjQSbfQImHhgmNtV/Znom1xP0z5kfbaGAhfsB2MCWhsYK0RcGPiavVk9mzBnEUoUXwp
0RYNkoSgtZRgH0D1UEf7/lizZutt0cpN4V8qb9Aa6EpiB9SESA2Ni/hX+6SvUhZtYiXQq1VsyB33
jUS12lE4dgVpxvnEFyAS9iitB4/nfGGw67xtNxRRHcyQUfWC+T82k5fiWBbpidMoSy+Ne+8yTi0V
iQcfhmr2REQO2SYY4JhvQclbkyGADxOJKd8wZfxeGsvRTJajpa7d6isOi4YY020tJEcxK6xXUbYr
nDvesTl7VXh3qQWKXtvmI8q33iYOP+X5savYbH9Um9jJZznCzCFj1qk0Y+C+HUD1k5fzdv8ri5yh
fqsHk+E5v/kV7stGka6wIRAxbRrcRFlUZUoZthbdP9+aEPZfFX6ccd6ayfkZRVnT57p5jT5F0oRk
WRlm9VJ1w2QwNhj33pMzWFGexylkKmIJxIM9u3eVQ5+l5a8GDbtsAHKJMxKB9Q82y04y0BlyPWD4
cIHUTWmkm7oF6sJqbgACqwd9xfOG3DPgcB/eoyq84VCmLf4OTFUrJ0o02hj6TrOvvYImHBKTCCMa
YVymx/siIY6oaqYlnfezyCOpZ59ww35ubw6L/S3pHbTLbyf/tmlP/4H1yQzbuNdaFQ4d5MnJm10O
4EFDMVhcQzT8NDJjZj4BjYQnVlHzVENdi88QpFgQOUB/Oz61clwAmQaro++Iv89OLMT2YkrOqINW
I71wRYuoc9scgCyDXo68sAD1HqVm/OIN85mJmkvtwOTTXOu44+oIMqwiNw0CSZwZLIOHYGuRauhD
mnFnGisVt9FKEG14K/DxItk0GTx+F22QF/7Vv95lumwQ3JMBUg9f3fCo4nNmMiEMoWaFKLCaTV61
6ajhmndscq1vnJ3Q1jm1QrAWYnQbxP+BQN24nvKqGeadU9Oss9tw3F0IK8AUPyqkXtCuhBcopyC1
b4ZMsfUJ0nHlq9WtEtXDuM48x2tIPTegOxe/Cfzw30s8cmCJZeH5BrP3cs/nPn73WWHulvGVCx5K
Q5Zfs8YahPUYh9SyNMSZe0gnzhyuRymEOHptlSUBXdBspKcteNXTtSidtxZCIrnv3AAhdwSejGGY
PySZQxc9FbAVoo1QLnlhcyvwnvZS75n5Xc1JDv8ilm61cBj06tlY7iKacYz7mfaah0fPYTB0VtkX
VjGOAsT93mW8jmU4ItPvYkb3j3gt/L9Siw9ko52lhl32aejMeFw9on07n3yFafUL7nVnX+hJMk37
zcMn4ZrhMtZI7ILkLR5dJ/Co4/EkUkWw0moZU9cDJWr8ICM8ooMNChfN4+RENqPK42Bi3vMuvuqQ
y6FIu86v8YK5r3eADyjpXxw7KxPJf216th7aqP8i0dgQeXo9s5cjZvvRL9ST48wv2nP5zxrx/3d+
GEXYrk8k0v4EdxzL6JhBDkoaV7r0NA0l5f1OknUHyNLoMlU4z2GSWsfrlHo4jP47Ct+aiighCGH4
FxVH1S6EPQP6S5bT5pqopnNhShGsUGDrdukKdLZdxY0uP7S68i8EDN9vG+VyLR4826T6xA1//92S
2d0QDRo+XtSmBwvEysHzdjPAKzOnGsn+2VwbKpyBv8D/Y/aIx4OhyhLBsN0C2PRluOSZffV+aeuz
59euP6r8NwAJ7VCRGt79u+gL14f2EhKHuZMSSqDpZA/2/AWmboK0UVyisnBPJzEyJP5S6jgyWini
nUw9eNPCT9GgqnhECOdTg4sG1MHvewmIemsBoSNm7KyK+zyWaM/NwCxkn2fqYO99sHBP63BfjiwA
yg18JZpmIO8FSwNj7V6gOPXqS6IXxUygtIz/znAnPn8pB3jax8mEAJrFNQPVT61G5ErtdWzeNPqz
Gqd5ih4LjK+hBgWsFFSXN0eUv/hJeuR1YdTXnpAbI+bsdXd3H3XnoSqIcq3LraTd0fZBZAAtcLpB
lfOVObazxM/V5M2d+1t55GROcPneUePC5+5Fthu3UEHR5rX4o9lOJgsDNbRmj2W/qb890WJNjGUq
fx8Llnot1FyODM7lVGxoS0BRSiByvsRcGsTeFPpzLBdCuzzTeEz8DlhQn6obVKtrr97COh/hv+Ez
X2lc61a0KPArrGPuX1cZ41Atcow21LFoUMlQ7g31u1aEgk1R5uE5X/BNtuClwnXe33NYdCHQ68yj
voW5iQvL5iWkO4+uNZM8kNN9iabH3FF2XZ6nCxcFD+T+57YDxQ6j2jOsutpeo+OlU67WxbXfNUSC
8idXynKHsHIR0yGFOD125/e31b4jwjJBEXRCLQYcPghTDUC49pSIbSy6PdMiPbdiUkApwLMUkOHI
5FdgSLEZ6+tYMd9V5+tm1+GgCaIWNSrL5uA4sCftr1x9CzaQxVWNEW2kC+F31lVMiqd9VgPzM9SK
XxS1ItUajJsMZ+iy7+x3HlrUQ5ZltyaZ+ZQNOj6EfXiEBpgYaWCDnrTMFyGDsNmICBCVEAqYyhtS
o4333gN9AI0UGR9NGk/EixxDHD/lWxeKUy0HtiLRpzSoRVRsWpQzAvaNrOSAXLJ+PtYwBSmxZtE9
WzdKCd9+Y0GX29OlJACFYL8R76Gny2q4l12+lxjALvjEhbkItbdlMW/rZ1j+xxJvir+dN7th/h1h
zFv0wB43jIgbotO0iZ2i90pfJI9692tOSsuF0j4dXjSvxI5A0Ac4ec5F2d3UJu2OgmuswYY9yTZm
Zj5qIiqytrwW7GWdF1nB7s2a/iJYr6Ugi7TC6M8eQzMgbAZkRTnqeLFRG1Ts4HXpIb395xEZZnb0
Fcyo7ncw85uPoF23AiBc1I4HluQ3Qqt4XkCEp0r1lNpxqpEQQezGNGWYYZ6RYnjhnMTXyQMT5rng
vYgePb/QxbOhfKrMxMVL9fnQ1DErF3nGXoau/agrWalTSi2cVA5/+XVE4FB/B5Z5nCEUuEXoSdvt
Nia+Ug0N/ebtBsmySmRE+97qqLWlhSWWAIM7gQVPj7v2CP0AeamJLGz8+eGWr/TValurFAS1lmPP
qYzptc+WEFaXH8JscMidfT5GNS48KZlL0TzPd4HNbjG7tk69I+VdBTczYIu1XtdxZczOa3nko1aA
O2/iROD3IKO/FU0+DbDgjY4+SRpbWApsuHlmeAg0eYaV+rLRtpGLKHfCuMmRCoyxudB4A+3fQ20k
jnxeWH/GetlG/+WEqX5KYWH1HSTArYonZQiWNs/47OOVBSl1dqwsEhQw6QmoTuQI2FapbiJSyvOm
mdqYtQ+RxmZ0zF1L+YICyPU8E7/QOECwo4nadAPk0Se/fQlegv276xXKJj3qGQ9kuwGa2GrF8bpj
32PffCPSJq25IbTgtm0xqd0jOBz+ein5ziOZnb1xGzHvruEtEeXv0t5+7HNXAtT6qLbh1/9CKgB3
e/FdIjGFZOWOerFFX5sism/CuxzKx+hsAKkadj5xG4S0dYYAOo2T378A7MPfhqoBExi+DxTH9tgD
KxwISH2hNnC5a089tn4/arc4AmzDIJ/P2UwkzoHJUAfPDqHs9UK8qMxUfr2HJFsY6BozgQ85mG2I
Axn0dsgylKKyOzCUody0AhUz/J/AmYTdnxou+l81ZUlilAbTd18UoO86A7paXEd1fe91dF7OoFDW
pgSIBx1K7wRPon9bYPmP5wxSuiNv0ruCWHItkeltUgn3MPOBQDnnyaUDLb89c0C4ZraiXN+Pj0nb
uDkWYAarNdPhCJZy7YeFUuusGaD58z3wTe16Oex8XnpgJfvJp6066PGuGrEdwCmnuTZkQtelsOiC
xh88coRTavy81t8+0E6HsaolrwSQxBaCUrBKH2V/UdP21i0HVYrNv1KVNOM8IfUYRgzR34vHh4OL
Wf4XjwZnG7cArwtYYKXM3SE1hWnST3R0sFb4ou9DjY5eQxtSU0XW9/+IebTNSD/UDZYdb+ZtqsAz
teOuuSTLEjfToBR17jKFvvCr4RfWvh0nkE8U+xnbQB5aY7l1n7oj0LEtzJ0pY7GOFXrch+bSlt97
LGpXkgLXl9quDwrLujGkJjLSQNU/ZV4Nx3oTPhBKiPgoB22MLoRz87mEpix001IPyALhm68WCZ9K
yO89XD71ivkMVY6INTZQqXn/fGFvSVhcJmNAJdXSyr0n53YL5djMeS7VBOjrtkPvrcWcUyyTf3La
WQ44bazRR96cMJXppxzaWwfEj7I7Skr9umE+WU3nPBsgFWG9HIh7FP/kwyRtzbu5OkPC/uCxtHMU
+DkJKWIFLiSmiCPKlHDN9Yj3VM/lDdd5wkfUsLb7qAnt1occGGQkr9J33ynbQyBJgK8jU2rRJO+U
/aAAP/dN8GD0WM144sflYsvxjFMsl3rWoYn61JF22XSEcuvTFbxnmxNq6qKdmxdXqe6w1LvEg7Pt
kOxUAZ7WdUq1HxQvuUSa347f9U/nxyP0XyTFnxY7pghJnurjUj6RRi9lxsqUOhtFZZAeTWfQn1yE
FfvXBqLHVTMO7tPyvR/W/yZtyZkGk5s9jya/x92k24VTfFW9IIV408fCh7wwfwoIqeeYnPUNcX+j
F2H/xR9deyBqmcGIjvznsFanCuhOVd2DYjyh2Ytu7KIPjpSFbbvK5Bof9PsbFMSKy3rm3hddZK2T
H9A3hC/DgG3X6c1+JidxiWWkQTQM2aje4gDWC+PcLKAxf+xSY42+tzIog2jnsIvxVqTZjAgTMFBd
O7rhB/9d6cni/PQ44S5CKVXigV2IzqOEAX8wJjcCV+ujHD+US72MjTqksZSA3J1V6+yeagAn8EwF
CCMGzLZKGTZm036ucGoiXNN1AHAFGmSsieOQJ6AHGEpNJF3VfxXqwudi3GNxv1i8vXK6K1zhacI5
Of8NhHOcSLmAUm8QAPPPjr6XEdjgPeP8i5wia6CFme8c3Qv3UKFO/CHLrOPahyqgeBUPL0HQk5oN
ESTgmhiS+32f013RP2vssfXLxqo5lrKupVJt3J5DyYYANmCPGSnZpa6t2w4KqFAOALcHzVIxXenH
5hwmRKox21djLS7pzXkKX7FfsMOCYnOTyiWJPQdlJl+zCQr+tGBHINtRJOeSThqwsPFUGZMnpdcs
9kT0WYbNSWQicG/EJADtHpIpymSK07GiLzEY5HyGMlveQy4GZdDEelQAI77Uj4dYaJdk2nRMBuiV
pO/3K/HSPmx5t+Td36Y7qZoI6eT/cDfiWEbvt+ymV2aUTqTmNn5KNdk7AfrqQk9FSZul74lJselC
PqukLVsn/kzTVeg+9AiQn8M03ptJxzulBd9rd2+kGepn1lRltPeoQ1WiCLvNQJCnEE/2X+zXl4xI
/dVIUha6i9VCT6rKCmBFCmzUbJy5PUlUpfWovUesjkr1Mdb2KQB9S5+0FnQR+pLO34eEYbrJYaOQ
LTUiN8wOnxQ+8htGdQNQWhcy9o3FU76xzE2+9JhG7pi4pGkjG/DEK3peeVxcZP5qVaDenXPmR07W
o61KdJnFCgp8rsBEto4W2lZDWH8bn2T9NiihktMMQu7b1axTvWhm3LQ/GFM8HKa34Zrk9ui9MksU
T1VdMKazg5u+2czyVbpkt0ii2SdkGtXUjLVvbY1fGVygvW06Mb+/I9u9vvGWUORKz38zIDkG6ir2
E+UVlaXK00S34PnWp2GWyDbsYEuySUdJWT7wYepCUQC/mJ4AqPcUzfXOveBllUvlITeYUn12ERYL
CzSCr1o6LLfOBMKeOkQYF51Y2uilKCoP9VMxO4PQU7Qe1kTfO4FjZtx0DXdLD2ueTskVCIA6cBoY
4uWizeUZtwhvqtojOgco83xuHxidgONdA0c+yuDjIAyI9mNwBdmVU1yGU9DUYhJ4+AiPKFYxs1Mj
iEb9aD5DjGbTtY4xTEktH4gbfYOXW64doXvPgXvTxC0dChsveCM26G13/6bGE33EmP+x39NGn+PW
hsp8d7tYjChJqb6H2RahODRZ9G7ZaBCC1N1GVdAARViyshBDNbbNdb3UpWqcFq/PCYyROriT3K4j
YcJGfa3XzNdSQVBlHe7jHY/Rt3ReCMcxYY4PUgD2y6kj5NU7itgy7rMGg6lFLwMipLIc6b9irPyR
r/nUKx8wVm5BkMcn9k8CTRtdAbBzksH89m3wkk5I7F52KS4ZlJYU9v5bjegV3+FzO8maHJEMo5SD
hiXJ/I3x2g/nK7MNKAeIBfno1Hgq+YZMh6dT1bExXI8trgotPge/f7TWzTkFplefnq8ZD9iklRCT
cPoLunNtq++2oEgacGHBwhFY2qFwAi700tfDZTfglSEysPZRN1/Z9cHa0obhm2CVVVEuxvTz6RD+
66jxdOVeX7LA135/N4P50Y9awvN+TY+3X3oG1JWU0ZcSte94yPUoW1CSATJ0w8+noy9FnPWaAoJv
SCbDCh+iSDDF/pqbyraY6nhDDjbKdHVfSb0c5TLc4FREDRF1c/bPQ/9jPaH8tsmZwQpDga2B0ThD
XMxYzaPjpfnQTXJdY5svMf4tqJ7yJ5DQ4fGXxZaK+VH+tQQ47z9seQwoBt2RJvErT4VXKC7q2Yfb
/vyZiZFSiUCdur+Ar7v/0hZmhK8xJEH8wTFvfmOYl8D7mfmYGB/zahZz2Qta+Bil+SHJR5QAyqr/
laWvX8XmC6hBAZ0FvI+d2MLlJNJsbSVpfaccYxjviQq3oI/KZLlXnFch2e8mSxGh9QhXvzYAyoHi
Nsnm1v9J1QVAkPFVqc5LhU6jz7RrHaggOkJcc296ihnTmqP8MZT9oauLPkyMOgxibrPwuYBZ66ww
zw7dptsVrJOLEWZcEAChVS+Tik8adbXpn4cO6HodYc1YUp+pA3nQYRtFS9QmrSGj2uM9oO/EJeTa
zoKv6Ra0+8iQr+ykkf+FYC6K1ghhxbzwYgEIeg8dE+Bxq0rP+DV2W7Ak+b6ZXRVxIE/3Qc/vX2Zh
s1DR2YDUDLw2NiVrT8xh16eLblJNmOVGzwq/AhWLnYuMXJXfWg/7ZC6yzK+hc4DgeEwCi/kt/qt6
yDs1QpGWKMdZVJ6r65kUpAoNFEI8NahvM/Fr1aSW48gaa9qYehsSVFPZS2Z9lkUYL+kue9zoo6Xr
wVO98/DnQHl9QQbTYD17hUVQSxIRohDIow5CgYyJe3umu437r386LB2vpAz8CaxLJKqo1IFbjZcH
nDJhDwxSEKLKR0jY7BPQkAK9R0cerWDkDViNcxdzD/HLGHZaUcv/U7L4Q1MAK/wa7nFeWMaXvuEJ
eY2Lz8DKZ/6vercOrAsiaAZop2RPrPiF76AL1m8kDCnsZ1porZy+FF6Da8oVh34iZ1hBhUcrZdWP
iHBCNlBDGPSfCGOm4vMCdfFqzGZDijHCiq+lsZCyYamZ5ys/JPZTAMIvtJHM6M0GFQJMWgdN+R2B
7wJ+Be40XFW3ZNaRVGh4Q1QDQlPAllyfyfcY1KZwJ7p83h7e4no+RxoS89gbm1USda/bR8nGmHPR
9hVTrbZBbeRIfiZc4aYGGkzLPBZqI+6l9cnzC3FblM3+SXQidHsN1UhuByeoqU033IEKSkgQdntX
0aQBxtdRbKizd+k6g1thdX8XARQNHAtdBh6RZnbWiDVXBl6iQge9fR/ajvm2B2ZBKiGnwhL/iq6Q
zJZ5X+fssX9/dwu9odaJfE8eEgUv4PhPIhtjIF0vRMR+MHZ9vzdvgYpiSNyRdk90OvaAMi462zdS
7+yfbqj/fNJr7hwIebO0bhNVzT14fwRmtlVguFyLgR9+MGYpcczdskB45Lm6BwvnSxW043eKhbnQ
3rppCEym4pZn/bxnU4/jxdzw/FkDKzjEfA6aKFn7W2rJLBScnkj0QxQQq/G7FRtn0G8RcnMdude4
UnH4DChOwvYADVODCx8o4KU4hU1Tqw7LucTfIoZf3xAwkStN5yFANYg0T12hlxqMMSyxXW3L58OL
/TAaweeRUCopGyH+Kbg5m2m+NJmIATh3rh/K6OKJF0HhjsdFOhQN4zYlXfdt30xhHZYJHhKfkmnQ
DocvCaEm2QyEzJ4U0JZYS18NhdM0bHVgUTb+pnNMnS1NA7WrEtQwkftFQq+QQFqIgUzqlXfjKBRr
d50aLL3D17B05jHXt8N7rAiRuxzg3pu0xOOgi9pqTozizH/SuP0Zs82lmiCXRHYfI1fzUYwHebL1
DMxcy2qpa62kQ9W7fwUJPIuBJs3IBz1RszegCPW24dSHCEm43wMd2vijB0agw+ElNmt9qJ8zFsDS
dEg85L9x/8kCnzYPxJLV/BTlyaMphPG7hQeGJxo+7nidQAQqg8rjj5IS6vhJKWG8ZQJJRIrRzhig
GPbHaB5h8YBt/99rDaR66Z1n+rwtGz3ERWHKhStoiSiFUoZfA+5nEGqHdviOFowGdHqS3zz8/yHd
EtxlEz8aU+EXppCGk4Tfio0xw8yTLvSXrgZpj9N9Imj20T+R+ZDoa/1kFMGG/pfJ753fO5p+li6b
a0z2hw12BKivVTIMwh/mMZZaeXTEtjIg+RKCDfna5ly/R8fZg6m9quCKq6eGZu3PR1JaZzRTFZvu
M4MmVAcnjsCH5BoRHy9Zi8c5xnPUBcOs5dEmWZGCvzBLz8IkGl6s4KMtq0TqMe7mz7vMzujFwFdr
2J8Tmv32Q+gr8y0A6uWzjaIhBzqFuYsVW5LGiLdZw3HVgDLQBUK6x6w0YaRnUBpUKn2USkTVJ3K0
E9uPpaykgEm4+qt6kngr/CfmdMzKml98BlfDgPo2+VKqg1TGDSbPlOoR5Rz/z0MoUfEzlV8QnZn4
sDVoQKRNL3QYDp+ZnWhua9AVW6vlyo+IZ11aFbzYtfOWckjowxgW5737LR83pfYo/5akUBnXpDzh
+b6nVIR/L73jQ8W8goWAoyjpiqv8sQnS07D/Cjras14oeHqamDphkLSHJ8I904LP9DMEnq6tNm9T
ocFoBjCjGOw8yIcowO3/QZIIoM0kcjSlOA1PZjxc318T7bKHlHX8KB38cPhT93a8oyPP1bBDBluF
923kiNa/6PARmfqxQE4bBpsLLnq6lbKsaviOYqGDOx6HDk4t6yyfHAioRuackoSI+YQD8hhbacTY
zoqi27YaiHNd1vQcZDsw+wbOwUm+jekl2guuYj/uYNrVHoLNMock0dy8GEy0jBRBX7r01UgGGCl2
fqOCvSgtAWif4PnRqL9J4ycxLlHXLKZ3FVdFXwTQRyA44EudqFASIo9/DZRciQeRm6dhhbFYmeuq
CsTBbdOePa/9fvFyIWJIR+nGQqZ5Z2pM0HirKM1G2U1iRKbGrMZYz1cpT7lmwjUZmzFq0m7bePeL
F0dsqEQ4aUIaUAtik+Zyj5i6WLCJ9Dcb2N6+NJqsMYIWyoegQo2z66bncImdyLMXlyU6bM/4uQnR
0IONsop84WrPZPKir8kDsH6LasrxDdEopIs124QedmzwLgqMC+vqJNPmgZjmeYHQUIL/hA67ESTl
rQzHGCKeclccZhIpaHxfxXz1JOg/53znqV5mRUyPLdVXR4UsLdnV2VZjTR1yc6lUu3K/+nhgh6fe
dF2W55RsGaiMAQyP/ZojS6PO+mM87ob48OiukieO3l4N8BduTY48i53zcMLJdNc/whLUnWqaUono
WfaVsT4fIgesqV0bTD/YuL/JEYMSFOwG0H5SF4SrzX8KStSvVBZPoOaijrexealXMP/jMdg2qzth
f1Ipc0OpFYF88EUMlT5cFzcRntVAUbnuR75vs3StztlOIQhZNA7lXHIeNJ0OfjPXG0mTDURCHSP/
2yit+QYSV5lu5Pb0W6nX6C13LpZaL25ahVIM0bkmzuJlhQL6xIgk3uydOMKim612k2WFRaToajDp
pG08UX/vNeqsOm0QCj+ytPr9iQUzfTWBZcPZbHJjNqpwInHkMSsMLSk3rUgNwrDOkV3fjX/2cIE4
Wcr7tyU6o+jK1Xc6Bj/jj0YlTOQ34Dhv2UsYPgCafmeslkvqmI+L0ATHW/xwqtYbVxzlbJ6PsRMg
9gbXnqAz7ERPlbQ/Y4Zfvu14bL56sl2kOe+hAlHbnSj3a5S3GvLKBjaU1xcw1xjPyRI+CsZLBVqU
cqK6h8RxqkxNP5gnUy/p+Er9FxYGnNmPVAhtoB8zZ+5U6XWiNnF9aB0yJez7Yhkbsk+4z7+kFxQJ
AS3f1WFwKvLNV5FpwGGCCK6Jw3z4MzLwGZBE3IoowyfbeFrOwxjCkTR6mKIxJfk5S6r05/jqQHeC
iP9+FDNIUIG6zivstntpZ/OMghVD1HM7iCz34rvk3WnfIFH1WKczQLN19+cu8DPGnFpk0d2k02Qe
68JXkBH5pkyuSXCeVX1fzokhSAShIM1ch7+xAKXQMBDvulcA1+GK+N1nygsnyHA+4wo+ZaFiYAuf
fO2fKHLKlcVdrlEX+eiJbLVelblD8apMQ4Pm8zHkG02oVLG9xfoD9VvPrv3j9VMCinzKKPJ+ud3T
lnsy7BIwXVwP/MtB0nEyf8sQZxlP8X0BWAwErQNwGTfsf7HA3I/AFd3DcFEyi7N0nlm8K6NXPo+N
uRhOixVqi5TlJNJ5xFN955MVgs9GZKPPh8VoCV4ySRsHLvZD78ebTSQdWhCFQJkEh+/qS/7XBhmt
0ckuR1pMsczIzTY4JKnoLbfCyv3mvW2auDNs3lLemsEPz4/T+Rj7fM8J0vzughCv6UtUNrtN2wkc
dwANJtinSxCZDFgzakc1pKsndmI/8Elm/W/Hko0zgf5qC1bNQ4fBW7xCZhXY55p06XAEwH3n0rdj
Ydv6jg0hkeW/RLM9U4JhFtAgkhD2lydrBIzK/9LJw4WkgeRH8GvSrDdfO35Dk+a/RvaKrBsJlcZW
MbCTyCW3CSx6Zmb+W7LHktJnn7eLQZuM4Huac0Gl0IgHh368X8kn7ClzUpjTODLVQiz+WTB8llAF
zecDaqbAHy8o0YykbxTZi+5Ge3MXst5BjC2wUGLb4VTBruE+7/OjapG7l2YZHgmL3PMehlMWKU8F
qestIGigVwcygKHmFyThI3uwNEgZ21JmG1dAmh8BOBuGRnEEMUHnvn/iHCxn/h/yUGZY0ufsuMDW
sCKoLqvK6nQlSAGG1x7ESCV/vBaHsVwCU1o6+oQyajcXwuQ4ThKBcy4JhbN6SUyhqXZ9rgiVZYDa
fTmnSDFvxps8R7/jyp/ZfwHJwaUjAF5cnPJfeULPtZ6UTV1RG66O6RHFXlMEz6iR0AHRnEUu3UzS
tlphiSXeYUZFosITGy2N0CrkjtlbU1DpR2Wkckkj8HXEbl/7qW26z0+YUA9k+7XGnAyQNPqKDsNj
l5m62+m0Wafoiymgw4LySqFhuNlzbhfWaRUAYfE8rf8K4VREECOuBZOcRD3HvDUG/uSjxYraYDVP
Lc3XBfC/v2wKgNUlzbXyqTm+HoRYF2zktYTnJ0hacEbazrRO3XO2Yo9zzIq9la49Kb4XsR7RV1+X
fVZZwvpJ+Lzk1YsUrAWHYBEHsOB1sWhhgn+hpCU+ASUyhM8zQPvVouCp3OO0OPwcYioZfpuJ+a2B
hE5AhcQXHS2TV9dMrDdweMq9Uf5YAzcipmvh/0XxTjFVNB8lT0CXs6BSwfKbEHaMqVRmHtP73Eqj
B+B803euBg0CEX/CjVjq2i4dmwQc09FyTnP+tdAE5eV6PUY983p5s+ifpzACoGD7/6BUFFpet2Rt
oeF8QtccbS76pJ8yfJbZsKU7XbOM7zWZkh3JphNHg37k2+Qn1OcWYn698r56lTdpU257b3TM24a+
9rUUpU/XC3CZOZtwV9tOX7YtJDu+l7uyUW39zZfGw+gXbnGOT1xJ48z9HVTgfliowoNNChTq/NL/
j+LzOmdsJdYpWueM6EcNXIp6V/JP1RN4hL5OzyvQuKIMQiJwHcsC2H0+fcmbvFzSdmlTpZPdae5x
0KBbCEYK+s2ngXbfMjlo+p7eAQvSh5xISqbhKJGxZh8nAtakn3t6FotrHaT2Y42RltO4UaW6rZ4A
f037zbsiRSB65UHqODP+fZd854AzvZWTpcr1lVt3f6gKA9xsfVTlGvP357iI07QvEhqIfIHKujl6
lMtLuxy0EGw1Bk/pmJ4ZGoZlh4ZSlivn4uFMKmX/x1jk2E97xX6P7jBkXjXSrSTDQrKIXj54p74F
FOWaP5nlx9Q3RVLcaNJt7PN2a2F2Hw4CbiFr80Zc4Q3XTs/V0RdPy3rBVCFO2LIykI21Uvc7+GsQ
2H0oRnj4jBQIFSp7ipPGQLQBqGba15EWLMaI2uVwz9BWV8ZcgGYQe03g/uNXru0DSbe+PiIVhY+R
E5/IPYYqYytuhvnNkzJ+WFu+SLk12iWBZZECx3OgfhDwjdvLULgczCZjUhxnMT41/4eOE4Z0iYpC
ux0WFPTHgzblXXJF79A6Od3f8+BY7eeKu8yrIvdxnE5TMBc4WzrMnSyyvXjujVB07q2rSTSPA46r
BQeJDMa6WS9QQ0Z4yt4XwhZtShlx71co30XbmNitc+77WETMviXO8XqQ8bBhNGNCrYUseNIP4IFd
RQWUDnshulmR8nhFDPNkUl+jaTI/7vzDiHwlhbtV73E7klizcBK6oGmjOUqAoFo8BxQcjAPBRj7V
42tiLyhmTgvx7C9O4aa4b7wEzJvYuR4CVyc5kQJRmh9xXkGYUUzqADq5W0pTvDcx7DNR5odsY9fZ
Lvxov7RzJJ8OnByZ1M8q12hT7zuvGcnEHmgNNI2sfY4Ks9eSVcwnNTN0jwr4qyIMTEbvFoiBu5WF
7rHqbFuEWoKwOm/6Q/sUM44kV+hA3Rj6s12cvMcq8/SnsNl4cni/qKWPBpuKwPxRa/RKJngR8HDZ
Sns3bVa/8Dyl8kqS8i3inGdzXvBW3G5k9rUc1Y5Nj/MML2s4yezaywm3whEtMD8XUJdcfXY+sfYu
9hjwNJC1oFJ5KsK3BzWy/8NKhZaNsj2Of3ldnnUW77cH4j/UcE944naT4l+IkmTkOvY91MJMx3ps
ONZAB1VpmKOgIJ3lAhsZdzBSL42IHkUXYwVrmok6kKaBoIY8RJ50mE0QT1nVAWFGAeDpTi1PEsVy
l7vsk/IroqyI8P9FK/i9PqCuKaPzHIIW71d60Gc5SW009V2NwMCn16EE7i3pjcARzaoFP7O5yda+
fEIBqNNnvhNtdN3D+16drkC/bnxVyxrmTuXZaMJN0bSwtZv6hGAADP3hPbFKOuicxj49HvEG9KxI
gqbb3dEllnvAXWbZzZPtwYmlcFA58IzVe3P7Bc32ikpUma5c/eh6DunAtyls5Syf9YOoALMoZGQq
DOg8NJbVJvZ2s0pYaiFSf9XsCkS9pCCSYm7BLYeVoq6tLRDUi53xRjuRYYgmRX/tKe94UCtMTbEG
CNQcGae8gRpsff1QMBKr1OPjvsdOHN5SDzF/zuxn4/vdxsJH0vF1X1Kth6n53PPiUCbCpy6ivLhY
4ybS5ju/V36yI2FUomFCqqJ5k5nFlTBBgWv+97Gkhz/30Zjlcn3u5mr3lnRaZVqYJ7tgidckKTvc
WLv0r/7cmXCZaGUjdm5Wmnpfjy6bOTRggu/kWR3Hgyvwq0VEeihrQi0Y5PjRkNsQAnnhuK1R9BeH
r920FCIKTehV7p0VJdqoK1HgAdZUfjtZuHWcGqHprzLlHTFoUna9uIoBiVFIY5oAL+y+dhPISaZV
Sz1bOqbmYX3Pi4BLlusXUmUbqGALa9X4lrtIo1IludrYHeeti38XuTEYtIz/lSwUdB7lSvRepk+y
grMqLRYHbYhv5gslTCdZtxKwyouU/wqxGpgf7bhKQaNAULZFZ/vfXbNrM3m6qqj6EWlPSd5ZsxXg
3On0VTTLCCZAvXnYVgdtBq0hVpL31QOd2W7lnNqtPLrQVIlgvapVEKoDYEEJsbvFTozn1PG4fz+0
K4Bc0ueJpdC8OFddR4JmGI7eCZr8ZimucFWIAbbj6xcjQEAjM6gMDHDq5zME46I8SSr0H1FPm+mP
qoyPWvk1vFetJmqHC+K+H9Ygu13Nmg35qIpZa2+905GQ5WC43MYh0V2TXaEKJIad1+kSskEJSW6Q
ff1A3T5QN8MWqKPTT7a9V8a38gOD1f6ic1N9ud9P4MbcxNe2LOTs+f7ZIR80clpe0HulIZwaXxp1
eG8VbubcX1Chr+/h9Dkpvw5ejy+GANcjtpGeVx61kkF+9syoU0Qkq1ND3Ikxx3miidpmxsunXrEq
+uD+U4LGgRBB/MwMj0DlH37GgKCvFj+7Fz07RlKjLITAlcQjUs5qmGFQ35kJpLn8VsNZ/j/FEG5N
6oBPXUGXgLMNfuDTta8RM9aGuMDSytYdQ4wYWQWVrszT1vEd4zDE6Lk5YAteyuqsEmDEJGVD5EAE
2NCddnguLVy5VbunSUSE+vfnPzK3gCXFAl6+ksv4qmUMGiCKe6/IiKh1hx/SX+ykZ+iaso0BuJDh
oWRXmbSFnuulBmITPJ1QghlmgQj4SuyiS0iJvOF3jBDYH7DhAR0KFRPBwVvFgHCGl9xFxddnerlB
SPVImcAbfPFuwN9vKNT1fm6nERa9usGfJiLT0feNhYQo0OEs/E3h9aCqDt0GcQqSsOcsO9YAjoxA
kSZHf3noT7mOjGy2FNahqKDc4Ns8bYQem1VyoX0B6+/d3Nftr3rbjUgpKV3oFMg7DUfbCLD4VRZI
Lxjg/eKFkRpJlyAh7eozeAYsIs56zF5QPhf7ymBEk/JyKio5y/+88Blco3TQREXKRAmt9d7GhXVH
Y2BN4qjK5LmTZcPZJuO2TW3xw9EbmJPStMrOH1ZJVhnXklJm+N3qogsVKIn78R9ivoO+/+wo5ANX
HpBdvb6TdPugRQTU/heFUDfoy+DZMF+48BomEO4j49oQ8cHKjq8QDIt4xINeZzvjO2vRmAGWb4y2
gC38CDZP5q+mDOoCPAnZVMv9V4gn0fHeGslJueeGm8QB+p8g4hpt7wpnL7NCqMtOjWkt++V3MN76
nrXawGO6z2JVc1YuN2D+YfdK36LnMptDkvaP6MkPlFexsplmruxsQeetPye8lle75xF2RGQVWRRS
1CTIXtxnQ/Tw4QqVFmIiF1ISq+wI6ywMpdq02VWP6Ltycr7LVRpYvJ4Dusk+lDTBp7jrXLnh2V+q
8+Yt6v07iXPnIIvS7u2mDYFy5VFd7a2nSH4+jrNK+HBWp7kCbdSZfQocWkyAFXVRhHzOOptP/oDq
m9yTXUErSuf33aXoTjggFo85AasEkLZ2cax5UB02jZcolusP5l0qMT6cwh0676xDNyGxmjMj0+Tg
Tv2/W96cn9qSZQ3MZVycoFOC2PWPp3zVH6S+mN+n+fyYyRupyUs88cl74rzX/fxjkbz1TjeIDkzl
ibWvnhN4ta/ivsSGnmQiM22n8WxMEJNyXlI7jiBjDd6lLe+IbK8MnuaeIgWzxPIshxmayR0/hkum
+38Tz+amVfvAb2ijsBrYWwdLPWNSK/NQpWdRrdBSAyRvils2dV7SoXQA8UIrN10pT4GWeb/Tagz6
Wxk2ufxl2nccvFKwK16/jmGU4PW8SWuKX4WLk0Xh1zS2V/5M1AtFYHK7CztdaItxs944AMkc53IU
f+jt+HkXAeOEQYqdLHxquEePZmUlevRYsnBFyuxwh4M+GMfSSMdVLj4QrkgZ3tasvoLj0nezPOZD
mF/R4ZB16dW1XrcF/QlkNQNlz1hvk88jIEKzxrGCBoXv4VpM62azaxL4Iizw4cn2QclfsPnqYMnN
yzOAWMf2G+k/uqW+h3Ocut5UKP/uuBJbzO47A2V4kBKTalSKpul1biUNWN70+UMnrDY9gIrt+nQv
V/Zd6brsnuWKpCwHau7/7FFcQ3GNXcIQSbIscVGnktvyhjqbwb7yCz5omyksAich+M/QukTiuzJX
eTRoQNKXx64zVf7f/9NZDhv3G3lrO12I+gGepBcJ4KLtiHpLXP05E/LLNGO04KmpFhsOXZ+A+e2Q
26jPscIbcrwlsR6wiNELs99a+Qqi9Cc0nCTzQ7l24apkCvTVg2Ny7qaONzjdivQ2bXN1CcOaTKWE
iOW2erxsMZop6N+C6ecMpScm4eRyLtZNL4bYA0ELKo/ER93BVo2Vn4lPr3M3XbB9UQbRGhrC09bK
v6B5QPefrxTdTeVmWroA2+Fty5AMwn2Bm+Ev3OCanmmZybRvRqa41hMXwWbnyXUmI50xkZeS5RR7
fR1PszoXRQM6LPLHQsR3iN/dtat7l3DK3oAaDhyOLHoYbE+UUsX7n23o+cB1Wk9IgKeWQ+dk0lEY
HHc2pKD0Rb3HP0sUN9SrGdxA1/CzwfcAlIQsyoTVxQ6YFN2xu8u317JBg5iAo1usps3vb6GBgzzn
Ukt9FjMNvhv1hec9U26+bGTuGG6/UtIRG/0Asdli3+eRiXF/RB6NkTnV0nv9/INSfvTd5+OXDTR4
U6FpKOgFvlgpgKu8fIfEVrfOAzcdbXHPoqw6mZ7EQtB+5/1ETlXOGiL0WMnpOlc2GsWtOujchO9+
RPX100Wg6Iv6oeAFnu3YhlIMsAS3B4jzxWjj0Mr7/8wXqMFn1EZPwliQ/uUj1tWg9/SUhuAiM27t
zR04f46fk+FCPmEexryWl89FABBFd9QPFt54ClnEmbqsrvGWvrvPBYkx8bNYSqyI2xxYgNVDLhHY
rhxCwVKaYcJS6H731/Nf3aEpZy4Wy+JOC4H2rspgAEevwRbwCaRpidts1Kzusjkgbk5P82k/8hW/
CV761t2Y3ymQ9K5SnQh8NU8cb8tR4FsX0alurWxl3lzSgc7FuucAizdpLEFHPmBbqAjomwJh4GfM
dNJRYsmopxxGJW8bjRT6lBYdTd28ytPMLH0isZTuE7lmqlTsVhY5727Ryk9Sp5OqZFg1oe3MN2zw
c7a3yBvTtyXnxMCcREaLXBjmI3DNFJeuTGb7tO5OIxvAv69UCc7dP4KcfVMnPa3Eezn/KgeSzekU
nVmEIbogbeq3wodmCsyXvt9+I3bgg/pA2psrquVVbSLGXBikp1lzuz41kdh0gjOZ+dXjdID2ij9O
20JswurdzOMJ/od9NoLz77WUXOLbD5Zn7OwsPyrbVdl4qvH3UC42+bWFkRs0eVyFbYsYV+azeJqL
d9/hDfp5+UGMQpNLzPCguuHHfZIFUNZRhqEJ4Q6RG4UIK7o7lHZulsiyrEpHu9WYRZQfaJcJrwC9
VEStDhqLLwVxWecIV6mrjjApCLRjxh48Iv1aNajl7Eq2PSlR+vk4L8J2bHORQJnuNn2HcGz8rheW
qCzCzv/7iAOVxtHPM6hLJFP0Iq44045s2stF4ngXRcsPA0bzaFA3jz/V6/SSYCiuglV/82P5w2FB
f5NZIsTNBfAjHKauPwq8z2DLosvAQT3EvwP+98cuUnKKjcd1+7X/c9V4Q2cQtujBXGP2WQG+umhm
i8/hhvR7Av7vkOHjOqwcNNE4ZlDd+zqTSvWE/L6vjF2Y102LVTTD8GckYp5uTegDux6X13m9kJLE
hCldEgj/oneqpA1QxuDcURrx3RHBXo3chvI3h96+CUwZ5T760u76LYalOzq3Wd+6CYT7jci2Qzsr
dypjy875dbXZK4CEPMghf/Pzzj96OCIxEQsp8BQ787zoueSM9k59k/VZnMeafjCE9bzg2aqVif4t
ClLLht9Ej0xY2J2QDFvmGnSfgztdJ/n2todwMbYLn0+VQAqpIfci7sdQpsNacjtp09Pg+FRbXseU
OryV3QKPRzwN+JqGpqfthmED2Vu87sHduwTOObKUSVgEV6y3na/2v1eLphfj8N1/24eKnDmj9EaG
cO6v9wmc6xHtHt6HdL+DSoO8oy9dudv/Z0+NOi7lW1pkjHnBzY1BBiaG8lipwH+ShJsXZSkxjG3g
ejeAQ3UxJSPxmcnbho+kYZEiaByUwC+eJC0R9J9BV8NFjR0GsH1zMOX/kujLjExATbt+rCtdI4CD
u5W9BueWh38EIdMv40ezuPxjad9U6P64pdP/i3qzqpgveXdJRFV94AaSLZQG6UYS6F8N1RUghW0w
3UXTg/6X6SElkqzpi7GHUUdR/fl41VwkzoU7CGsdb0v4KxnGC0Mg9iHlG0j71uJAJo1CD3ajYgOy
IAawypuqcJqVWTJu/UiXVtZSPva6TsBibmFU30KUMWLb1Law06cXC8c+EV2titIwzD9uYkzzVCMm
xWpGLrmyLm2rg9g2gZHBesOg4UteT1FeNb/0k8Mza7RwbpcTAULMm8PbIopw5LicS/5hMQK97jeR
8u43gok4ZoQlBwYmmlHoxkvZy1xg5QC123ONysDqbMuywpBHyrL/068NRTk19F1Gj4tz7Q9Pi3NP
4K8I4gKf0TYozMTpkc4bD/OsV0WDvuibcBC7oSKDZfbfOnpkNpJs8LHRmHRMEeAUESQspbTtxrA2
+jZGV4YNOx8x77LQXiZgPHIEdAPVn8USD4vKpncErX9cquTwXSAZGzswyZu7JAs1VZgMleYcXjCX
A0WuLrQdgjTbKgYzdcPBR79PJgyRshdhW79CwR356FKhdLtifR6s9eHMWwfDaht86cibJSUbMhyR
uceyqSmzjmQFC8IAbxTGr00rGjNiUVjDjg2be4TdNr3j8NMxz+LP+SgwrA707Qfi9Z3KAva0DJbz
alWUPRvKMB+tLq8SIvxgksewFoHE/7Eb+IPCTTeUlPKqaUCvwCPsPBMtgVobFYTmG0rL4CmpV8b3
to8rUrq3HDk12VZ/IB/bwvPrOWVoxuKVGVLDKghjXnENwh7lpOB9jSfISYlkVxBMClx4N4Inwlgz
VXXCUJfWchRMaQELarPoXXtXVxlLcTdWQGlUYQFaDoiz3ycS7lSaJq9v3PK9Z7QWR5UaLh0ctOx4
NgSwI4pWVWZUooPSt1T5/Wh2097/A/rrccvCMrDWWUHEUPa2+k2/rqzeDbdiN9dXDpssrUc/2moq
cWeGJ9E8laiwTpBrRhRXxs0J86t3clKLAdY9M9ZYmx11aBnnSoFWd/grNMBxcR8Gw31ODKqFxekq
cX2hEKV5maW6/MUH8vm64vVCU4aRls+DoSBaMQwWImVET7QCVmf2ObW6094lxTvmqt1flvZUHNwZ
ewL/zUWztGyk3qU23o3IKEk8WXC0Ug+HLZQr/Ipdv23QyPceeA/WtdgCkLshCbi/XsS1meHSkMHO
tF7VoXur/BbO/16lIMNECHcHVykboLkadKn7SUw0zEGBCkTKJiTJ1Wu1fMwVOGZXiQe1TLXPJjw0
quqmtuf7JZrqU2HLDTuHaMonquEmye+9imaMctGNyj6rWiRTx4TYT/9CjIyUZ3vOtQ0uc5uulniV
jY9V0p4LVs39THl6ftL3c3H46pzgtLqdzgKuMFw1aYpOQ3mBQzOFVuytgnwwREB97cjuuo8patI4
Oz0+ts2UkGfY5aG1qu3pjXgbfC7rlLtWsaSVBaPOX75IJHz8nZ9CdM6dCVf9Hlce09SgHjJgVb7y
Qp7+40waGACzWCYSpZiWHUCvSBSycSUxIWY8cfW9k2x1oEnCxJ70DzoPvxqEFt6bX8OquUGLzdDl
BSI0C0uH8sWrK45r4i7F4agv1kmEMUFDEYTPlGXmuw2bIDnwBagdxbIXMiM0zaCEuHmvWG0rmEpo
Iq3fpRRW0IV4xqRR31rCVPLYQS9tjcMH8Xf/Xg6LwpIlZ08AtZPDK8a9G+hbzx26NAgiHR1P98X/
NT61499KgwWeLhzl5y9BJX57jDbA1LDIlBItq+r/vCT1Pl/pKk/j7E0AXYzVELDDSVuAhaEMqlPV
ORGTGIstHolW/WyH48gj0azQqjmHty5VCxxhRK5FiLw4CvQQvAIV9xMxjlsI5bqQIR6DtunieYYC
6cLR+UWZ7hBuYbVRlEMEzQyciTNCMi14L61iEc2nm6WFrU8ajJ+QS+1QFVh+oW/BpCR9xZUQRfTN
MEVTLh/tOzcuSIeRH5Agfqp8P2cBw30nFI4PaT7LarxmubDMcn38E5z9KSV3vrPG+JAIjwpUwVBO
zaepbN8KzlxPFWolb2IqLGcMoN28FQ0bCkc0q9r4JpO+MQ2FcMI5Gs2j6M6RPmZry6g6P/jQ3URN
Vi0NbHbTm/DzoA5yYHLpZbPfF9fFA9XwBI2yCODDgkDeodv7X0ybzg+guKQSZdwbE0ad2Qsyk9KT
AqGLY7bn6cNb0eLuxuYB/8pYg+hERl7n9CGEESIXqFktWE4WyGQPhf6dt7DKGL4CjoxbXpF2Ut+C
ucg8auHSgg0z7+15WaItnohEmxFEw5wdsypzJDpPf+3dFB5N/cw8UJOhZ+4LAVZTWC/dp8heY1vB
21m/SgsLJuZV38T7RJYNOUhFcbwEfGmOCUvJog3ImXxaYHw7r8INPOOJhXyLt5CB3LEK/X1WzQf4
a2wswhCYDDw1tc5+DPA1GCkC0fx3jBduZPj394Sf1HF02GBE7HAsO6wL7kEH241oR6WGjrltNiYk
qaBOpEuJ7Zy8J+HEydEkFDDOhP2F/TKvnj+MEYzADOjk6nhoTrl7t6VNAPrdHKTzi8DpICcqgPAr
BNHqqo2Q57zho5kurRM0V2v/ij1uFCL1iXEe+ziVvskjP8JD8zg1mm3cBIwK6EwlpyUvMbn92ICe
39vznvS37JafSh0fyHOVMX/aEpJ7rafz9AHCZU280wzCjYZPcGfIkWFNyG6SiLQcEB3BCLzQ0Jjb
DL4mDsaoQsSO+z1whmKv41eKmZM+ldm3uAsgS57GK1NDcf5KhDKHbh/clhCKq2TOR7Ibr6DZsWwE
eUke2XhWacqChSD4TbXQVDLPY0PpK/UQrYEfN3xoVwMUgmlc7EZI/ged0TWihBdhkHe8Rn3DIO22
ZjmxhX8RRWRV+g5njPHRqH6h8TzISBwR+hhbF3WnF2FuyqVddsuDR4bQg5b53kfKtgcfGCGqbr+i
wTWC3GuAuqVhikE74WKp+nAvVjb/5IOxdhMql0YpNyeSJ+f2PVm9RNBirSgTnNXXqUjHzjz7a2W3
fyi4uwSJ977y+AW/kx2OrD7w5w+s7zsQTYwhrz8xeXTVu87BOREgTDTP5mxBlYbubbpRT0t50FSN
8K5OtYfbXrQNY+Irdo3M4cRMg5hMBehqmdrl+sRDEELUHGQfSAXGZuvVRTfnHmBVx74uiGQ6dRhz
oV70VBnZoIypP9M1Xki482U8ZP3MU1KCshqsuIOsTRpWnvB5HM00fWwBxQ2hW21dmX00K9E9Tn7Q
BpErrUgMqWitmJYomysCyZ2Z3+OOIcBYm3h89hV8bUM012yu0Dczg8ti17whX9EgqR0aVxdC+ZS0
VjLzMudrUrgIVFVDxgabd3XabjrpkgllCZLZ/e2oQ0NwOcI7/Rqg/7E6fjTfBCmOLyiamAZ9VOT3
c7iQQHaiDRPwtK3QxXr8SGq0C4n3UWFC/roy4x6eAw4DnmuMKcPLz8LSsxO+zD+XGtzeuI1UU5ny
V0PmFzAmx1Wk7eB/VVKBiLkAyNHTYrFOHZ0vtKfe3x05KmFrgwCaOzehsMl+LIFKpMWaxonUXigZ
jRk7guISs4ZH6Vm2CwfzXDw8jUYKQ76Qqy8ifjBYePmqSm5jrNga5zqiFdMFmPAXfBpbuX5Ai0sN
4jlVpqryToRbFC0B9+Yys9fZTHunyAKJ0sovXSkB4t/79/jveM0g5WLwdFr5iDCvZVAZZ8pVlv98
Op9dymzLGEXfXUml0Z0qLOqdLP7ZjLXLoBPivKUfh0es8w+qrvRGDIjzKlgzIfET7mfBNxODLxE1
o0kFBTuQRTsy5ZgYtzC8FukSz1Macwrq1Re+sbgmYZneUbVfIYRNkMmPblhCwrF0/L8LyV2TqbIw
kcUx9kOkxq7yL5bJR8yLJCvXKatdlgFPFlL+/aNAyMrt7dWbFOOo/L4W2rTKl+O4nJk+RM4eZE95
3QtwJoHbqh/qJaJKSBk00CKXJVayBzgVfqqaHa59cAZngQMHiPNYCOSkUaPu92LQpk4fe9o9ifY9
PAful/TJU71AAZaStaiG8TqnMzriHy/+TrOwMqdopBwztpUIerZFFWQFUIUMngeTRKWqmL40O6r3
89Xmm6w7AGVmByDZ4g5pysgmrJQMUgVE2nzACUvOp5sD6FR8xU4/g8Ml/whkMH7VyXuWyHvwFW5G
LKC0kjeyxCzcTIhvTj9LVCq75kat4JvjcrMAtPhKKbryZYkhv4eZ4SFVxN3ukJhQ86MTT2RVYULc
S4zsuGLnSRX4/O0VXpmW4r5N5E+1oLvKBZt5tO1u7kuOoTMsVb7n4OzRXN/dccQYtxNRS82SHqUD
rf/eKiZ93AXmh5zNHYB9vo0nmoiDrcuyEtof1e+CoCsxgUOGD2IKfeArFFD88aVOtnIRGexfXuaw
wernnCG1c7YEk64lsrDpvI1RM9AatqzPrY+wasTsClqMEWBoIh18BA4xOTt2yBg2fOzkZQl4nLsT
9TRMqcDw6ak4u2VnPOZGF14Qg+kMlezq+vnk5o/Q3ecpfiu5PWC7Ek/JPPeGEKShmXxxER0sQn6+
P2auI6bDqYKh5mMunj/gBuuNpDJCAG8jQnTN5+KV8Is9Fu6EjIVZlv/yMvwGgvDvZfTAYqd+CTKM
CdIRNIkxFdK/nj83goX0UrDGjpid1p6xMz+oVBXSWPXf6unHgXX1bJoQHPXfNl7RWE958iJC8ts1
4l5O908RuvyKj3YIi2zmjU7aIqv1RLtIKFR8PJTpostODzmKIyWxT0Ucc5+MXvi1eQg6vK+NCAby
2O7kNQhZwzpDW6w2Lros15OLPkhKWOS+6Q0sYqfeItEnRDpGByTs6lAWHTvEMkTkbGAajF+NvXao
jQEwyIUyKF0Bk85F0rJygZG+Rr/ZJakQDyyXXpPqP0u44/MQt7cSlfU56my2EVB19Dj5IcdqLdtt
nHgGkbhskFjJ0pjwGE+TTJB6Y9NydR8+/zJmsGdLxf4jl+420OAUB+EgEjTUdb7mbXGnAdDRyTXC
FDh+NNg6iU7n4jFW5gvuL7F0VbCC/axvcFwgb6tYjkscHEzaHrP9+oNcl+eII+om8Afc/YF7pwrS
63f8b51PyKFIFCY6plz1LGkW0OeX+OgAxXVOwYCNRsWcb4ZgZlyOAMmmy3k9rhBIlZ5woiWsVDwk
pafXYwi4n/pyEaAt3krsj3imV2OOu8zXswo8Aj+p4+LjWceJFYxI01Y34XFEnREvbFWmqdwwQeMK
N85vrRjIyvMXGdEryE6dqWbgrvOr4iA9NPPIbNhOCdtZ8lubSW8eZZSKJ3ApUTOAyyhcpWigJfvm
rHbEWxi9dfNlLIF0JOe2EBDpdv9jK2iG3UKjlDP8BSHW6OuLPmbEizbrldOnuvD8K44Hrn5URATx
c5sS6YVCRxJr/bHEkRuceCCXxSlHEzBb83z4CyWyQw3dGlzOganqKppIdR4jecx+uXDXeI8Q8HcE
0tfXasOgzx6O5srs3kt/AfoN0lrhuRNTbxWd5bH2MX+Gi+lye1spduXdawCXKzIgu52K2yUUweCd
nwsF3FOiHEQGnMSwO4pe5wK3VBHDE8MLey2OKMTcJK8484r/XaqRJVH4ruxOhbH23GmDg9blKqVP
p3fSU5sv5ZNT09/uVnpx23G49/xbfuyuM6ck6qTlMkRGdR1rlwOwPhYSdCtvlOg+6lCPx0i7xue6
ClWQkC49ijdimVJEF7ThSgbJWPLDRgDN5geNfEPHhnZON+ohD32cg2kPwKgMc+Xm8+9t2r9yAB/j
08XJcrLWBFnZtdi4EHJPpOiXgIDTQw0wd+h/QlkOPg1rq0m0zVHqQe1j69i61CXKk5zcAmMPdgt9
7zgcaHwWJprIuHUeo/fuzi/DO3qDh68ltiVlW6xYrEmKnokS4sHiSSqM6geXWjdhP5OkgLXpUxjS
YH/MO8q0jK0RMpJzbf9nC/+J8EpgDfRji1RJMaqPm/U0l/8Dh4r7GjYrzUKkP2WOtqSNnPHxZbgg
SeNLR7tFDjCbys1E0mPqkY/cxrtIFxNdZOIMsdtDXFYbE6USl0sfGy2lAHsI4A1+gi9YqfDvD5by
nFoV28XnXN+/9H6zJodIMBRfXeslMNF/FhsaMFcPuWU/uQvjwccVcWuqVQKy6asf3kCECPOPf7GW
JJ3T+J1x9EKr7N4cUAFyzfZKmB/ofLEKLfjLpvF/6VyCGmw5jFG8kEAAzWQFiepJwXk/t9vpzjH4
xeolE6fnJpisuCIBO14OP6Oct9BOMm+sJL/a5jOUET0FXEhtcdgGZOTubGsggcky5AzfKIaa3vz1
h8vrWsWi2H2i/05bE3x9I6GpwP0tJpk1ixY3/2Dk0u3Ky207ul1MmsgXlLviRa/5393j4EJDyOtC
q+F9sv2ieSPpZShvN7dDzKXEkCUa7JYacvKPHWP8yMLNwjAW7CW/8IR6rtp1ZsHQJR4WMKpAlMho
U6eYB/LJvLVtFpA7ncswLJoHWW/bcuehsafn0ZiaT0P/aU6ZjiaanoNaBf8z+yuSoOL/fb3EdsRI
+8nDGVSXEjHBE/DFYO2Bk+GMwPSMg+sRqRcG25B0t4hXyn5DtYNvvzbK3KmC1ap1BDo5VO6Zaq04
LeJo+Q6njk2JRg3UK8pC7uARuW638N9IcS6netl0kDmekwKu6Kbgza57p7h2+i1N8uB0OLzyeub+
pqR77I+xu6EN730AN4F9i5Ld+UDLMRX54erYqczEyOpym/04g3ooreNg/gHEjz2FujN+xnU4kdU5
XQXEf1mxsQIWabvvexUAeTjSKlGcZnEVmBiE94prqqLqWc7/PawIB58JtvIc3P4S22FRfMkOjShN
ZHo09RECMzONEX7mKQ+eEKCtMJr6fS62EtPYophK24YYerSxy3wOrTUV8gp5uEGjJDgim5WbI1J3
7NFqu11sTB/zyqqFWDY3sarGabuLSAQOP8ajiZ5cl82GyeJlqfjb79u8aifQwOi1smQ7bI5Dxeg7
M+4aZKLkA8plXb50FZOCTRysiapz/Ebh4TCklMiww9hTpt45Hnemh/JB+RRQp+9rXwV41p0c0HtZ
77/W94/iV4x08HCfawGcK8aLMMz591lTF/dBvdax0DhfyTcd2TPQb9OBxPneHbeuHWDOGuMAffKH
YY7wxeXI35B+LxC/N9hlDG2Rgmejoe1MsOcJPPnMMMGvzAc4gPrUaVyNKSg2jlrvgHyqQrgOeOH7
VWNpV4lqdyAdt1JikcrODzExPF6EvhV5vzuDrN7jnLRs13N3+YPgpJBuSdJda2bdPO++3dFwz6HY
LpsEE+q5qvr/9gPBxnBrI78e/CYoh96VgmT5xu/20LBiycpHkO0KSkymirtrbNlZJ7isw56IXV1b
o1XoQhaCOvxBGZRg+IRUzBh9UqysB/HM5hY15H3gWORcKlE8j8JfmSBcQsxDaKFSEiE745a/RcoT
JouvoUlaAEbkMH/jIyTpGxOyM07SemnB7e3T0lDvpx7vIEF1qrX3G5S+dp+sr5vDVjBpFe0p4UrH
bPFq8GN2F8EjUSBrVEHp4Fns/pMQmIEX9h9sMnHfFoXAkIs5nl0YDrYIdb8nFOdOtX7KkPv+U9Lh
y1jCVLfDlt9En4+6b4Oib7yK+4siPh6YuHiGNlb34xkGuAXnP1GLVGoJjLRHsDNd8j7hXNOnk2y9
fr+GAi++xtqUUXQC7s+N4U66WkMRhL+eTsTlCdLwHlmV0vufq34qLPw/bqHGzT9gfO+qdI/xpITp
+DgSzwW5DFVRU64oGlNJZtOnpfy4RToMHvthqMIE6KrKqRKBeGcUnAReIcp+XV2dESH77/LxDqY3
CtOeiSKV2geCQEg6tRp3zu+M25AFiOxDn4RLvAlJu2H48fhAoxifoSLwajaC2l1FMLGv8798FGlV
YrTmF8YDMKRb1T9KX6dMoP7vd5j9/ktUUKmVB8kRY58UZngFj4QhJDxtXU3aFIWrAJtzvwiyVEKz
S17tZK6NTWrg89rPdJZfdvqOatpFqN0Q0Dk9qcm7EA52TE/21JYns+zZxJDLENXtZRAREAo1pYtb
ckZz1bh/ZoTVLmtsmOcnOhPKk7Rz4LkBe9XJHHmmd1+IgbFgysxsbKyWDT4rKnCIsVv+HjJ++kun
l7hF67+RjCoNf1D1AhZzfAxiYn3u5/T8SYCcfYEYnbakx+jBNXtaMCXiwHQO0UnDWGMLLjxT/5f2
GCGfCrRE+q3Bt2/p4JW45ek+DqPs0n1lsIvBCPw6S1xT8g3YJmNmAchMJKz9xjbdVYh+l/6E3nJF
hTRE1vXgqRzSIXhXQLjTd/iwnUpAMP8DkAdQrsNOLRD52mZNB8yTOZjv3glrRnkj+ZIOfYhZJDdQ
vfR34/nJLvOEY4tauh134MWyxdAW5EFqo6ZnLdrekCGS3uo4+yFZa1zIGFaWHxYR44yaZ1BJgj7r
+HPD6HRjLbTDAHYyIMVQmA9Fydu/1zfCFSyxKduK6mxWz2bmpuEcfgDKrOblm/bztZc6VO5W50Rq
eKB6UkPfqJH3KNcyjwj+YKIY8j0jDBClBapEjEPEpV02PIq+DRzyH7SOqP1Z3emtQdiW336k954h
juJnz4HkVQuC0D8xca96MJR9yWUX6zp+bCxQcvoxzmGYBkhFq/ppaERZMdhLJ0KSfIbUe2DpJJhr
tCdXzzC1RS6YDZS/YVWIxkGG8YPiMRSl/sav5GNoQED3V5xyQq59tf6xthqS9dgoLugD48F86TVm
nXP5DS6r6fGNbnjayu5F4ovDlcBHEkgcduXpl2a4pvfURQD8YrHoYxq7GyuQVCVE/aLCLxpWES/e
5d82+E1dbb9rjGhYziVBia9v8JzJsUyNOUCtO673boU3tQ+uB6vAGIPubhhUSJ09GzMEDnaXGcrL
2KP/wqiZYb0W5EJUpmvlwPBToSDPJmEfg3/mEyAiZADnrQrW4XXBI2anVy948nyuRiQd8wPxefns
ceX99Y/4zBvSdp41rhM1WZns0xcJ0/JsHUgPeqT9bPNt6pMlsJOdAH+Izydj9PUvZwHNVURw8OVC
5UE0VUbHkH5ZdZMasJFcL4p3LLJN/LtvnRE/ewkRInJJKyEpl288Bv4iKbH/06rYn+SOPUgvuXFd
FIU26rHkC2Co7mb7gQ2Uwykq5mYrZpsGagtxRuONkthEkZ6p7YlWnpg6uhd9YnoO3xpgrvk+jl5R
mozO52XOQYK9K3K6VK0uw7HTYE9TYxC4IpPwbc4wSyaBtQiis9zYcTKlFnx3Es1Qw8fGWsWbjpOu
Bc0KspJ7khN/sRnOdumnkqskmDT46ejgYxPXOh289T6i9Yn7qT3K49wxOW87RN1CJQAwvTP895Wu
Oelx4q7ceLLo2bzqpf62TKRBX3Q51xkjfaGtMdac5CO+NIyaU+bgxvMvKjQW2fMyrcygE6ITt9Y3
QXgiQbEtNqwN8xNIPZ9Hwjcq6W1K0L2VQiZFtk1060lEttJjLm/mrzBN/oHy6eKk7zxQt6FeNnP3
qFgGNRDpWhvQYN7i7luhOU60yKE5FIJgOMUGXrlohCa1pRi9q0KHHqU4dIcvtC84fjAdA/j+YxyJ
2Haf6HlWYRPNU8QWXqtvJVQrVQOQAcCRtkcmuE5j05pKBlcx5F9cVlif2+ifYyKm8q4HKgbkGTjl
qjomJhpfexXfoBxEJ10M/pp3kuPEqVJYEbbvIcDgPGTjnm1NYoeCriIeE1D+H/s+oGT94rAdhnzI
NtDkv4pyB16c3/OK2ko9iFDxexDjOJ48IBIt7caU9Mv/RCSy+AYUyvL9ie67FLr9qAcR74KTkLk/
CcjHNuguAAQRnzo/GErD2XZRvw64Ux9LBCHZszn3gUQXwiKARZMHhIAS/q0DmrdZEsMno6uROMqi
/eUmG+Bl6bUPjUlXMekc4USi/Ee18h1vbXWNKpZeOMaPdJxxiGV0bLy/ogHpi9fCr0nTceV8ue8S
zOm7tvfvgwDzUmiELUpuRPfjNxLlcri66LD1DYa5AS5C4ck9LFFK9tDtNBa3XKIkQG+Sfn3ETIvp
4GysGVyYTORhPqGfsQXMRxAM7wTiGyxbCuY1taF93zQVDvl2S5ZpLTK+ruNz6Q4AyW5jGyFNU9Wp
RZVjMyt3BJPdaFbTdrR/7LAYxFyYy6G1OWkDS+izhQG+tBSCfKL4hYFkC0+zr+Yt08nHZdl0kOWa
3RSwBzIeua1MSo+bkzoRfSBpPHLc/mJ1EcChwhF4UxdHVDSTNc4hNFDZq9pFOvrNvSgyf1DPWSea
/igReRAS8oqNPAMwdFskAWPH908gvzm6XU0BBh0i90V02DTx4sOCsOeafsFflOda1I4zRZxRQktm
e2sN5f0pjd5sRGzu+9YhaBm6841NYBvfq8berK8LnWqK9OTVhMUDpIWwYM26yRXi3Q8UBS4TFeAJ
v4KD0vFm2UjXw3UMQZNI+02Mqil8BGE2g67QMsV1p/P4IvYgQjM3RLEo7r7j6fwM4d6/uG3szZhb
rVB2CeGZ7HjiDUBcJ7QAfeCEwTK+hRW0lQ9/fmEaQo2fwI5ncnrb5WVWOEeAHKkqi9GXlKe4deHY
WmDbGo9flKw0gMdjN8Di3w3O53EDKbLMYrrGjFZF0zruzSRIqy5VjGhnGxWGZwJH/KtlhrNKitKA
mezfTpsSettp0btEjHUTNfVDl9vEKcP5ILbYbcxKezLCzyfZzUyUnfSvNtRJ3p34L4HoTvUHpTXD
pNDCUri+2wbyOgfnv4jyPqTrxLynUxdEcpB08mQwWTxzTywdDRAo/EqbCTPH272PxSKfyL3QVEm0
JU8X5kkl2K1c4Q1hZ41580zG+IcSd8dCh51v3ik5gXwQvJEKb69r9LsUGsBJ8rHxzf57I2r9Bqvb
3RybTSbeEt/Hbn+F6b1BKUD6QWUF28uJ9OeaZFuP+ZfJRA3IztD5rc6JDzRfWir4vjB2znA/tHZt
gkyHDmqyN32zfqTXBalhSmwVYAInmCyAlPijCyOjxh3UQVhda80l5xcVX3b5PYoS/pDApwtSHcSp
hv+fJozLOwI1GDkRBne9m3+cHSiVHeG9YLPTiPHRTMXbGtlTJZzjqphidias/6oxLIsKXj3B1K8K
w0xMJFVXe5HnTfVHT15uW71ij7gNf/n5cHL0d5YTjW3GSGX7aEHNesuH1uyUaed52ag2J6rmeSjc
sOB36UAnrbmwQWHiJ0wjUGI9UOD+9jW/+I76Q3XSW1TLKZo8tRa4nyc1mbKViXoCwd6ZgD3AR8HK
gkzgkOvYz/Mpc3Ah6kGUWk05RRgTGNdtuFxpw7lOTEYfbTINTrj/0U4Jll8JNpICdNFIiA3wDH7V
2sIhRuiVoK7GMnc9nq2cLpDbtx1nhsqQpMiwoUKoatRLN0teBign5MnQ4sf03dMfVJVdzdV9hN+7
Qx7+dP8iHCQlNzxzFOMitx1qcuqAiJP4Oi6XZKA6rn4mBJfKd3Qq/UXU9Bay5FRNG92OiUwhOGWk
1UIZHcPp3Hhr35tGhwqyNLiU/tS8SHkKR1ZKbuyzSFAEbdM6mCoIiOMeclUWpMKCJUheoll3zEkj
L8tsmoLf036ggKyYJ+ibSZYFSMVDdqDXLBMMy0Cg0HZEh1xBQL5Tpes63AR+x+iG5pXlD2LJuj2l
D0LBiw6mZwe5x1wnqofR4VE5IKLNjSBT6zuX6ehfIU6zziBetXS0fV8lJJ+SCBN1j82e+Cmo15QG
SaXNMk0+naVGwez71+ZQ+DouADDkOQZij3HP4KOXz8j9bjwLagrQUFeASdTiplM08JAmYSFHrq9A
uIj8Mu7TdhSdYsfwxtIYgMuvU0POiCcoHzUAW9KYCcH56KdN0rSzs4q8HF1cXuFxxUhxcjeoECVa
gvF9X0t3lHhANvjgMiXUf4/fCXSQLPB7Y1GWmJAhsKJev3gMNxZL4DCbZUuZ91flvxFriwX32gFj
UmmNXCaSq5bbbTIK5HMw2xRYTSlo05OaJR1EscZFfqm3v0BImBr3nrnAQD1PYjpc4EKWxxW4N2jn
LW9cUu5XsSqQZHA6OI1R1gbmO6m4ZKReiEaNRTsTna+qrM+UZbd8yQv5NP3W5K/wkJrjCfSdVuMF
Xjy15OurJgbz3C878b2U+a8TkIbTHoo51SXNW0AAywdLSeBJN6UXnqwbjmfItaANovwzwNae0Wyv
/6+djbMaW/wQcYb0TY8a0Dp88qtdBUMrR2+ocKLFG3doxaNxUdLXXna1oZsn9kDukr85D2dkJ7Qs
1ot1D/eGwsi+FRS+8jZdQ61wvQGDP1dWInlrWOS9QRPjdNRyyjf9z803fpuGVNBQlAZ2S6oTCGxC
SMoHqm2GlAuIqYJr0OzlAw/pLd/idLo+My+RRmjcuYLkQOfoLeV5u/N0Bd4PlxcqSrPigAoXz9oY
JMlvZQ5Te74iGJS5mNncVto483Y2ng0hjPcjkV0ybdSSdO7zT2oeulorOsizyanWBzuwn3KFveCy
IpMLoX4MNmAMTxeZS60eLpLmUw0P7ghic70EPRLqKgRlRIcuHo1Ol9YfN1qrk/N5kXFNRKdfoW21
Qmpn+cD/TF7tm1QY8CpVKozSAhH6buAfz0aKMOfCjSTmmnoNe+CLP60Y2FwMVS6a9Hq3IEGKWL4t
J4KLiGrq895c/TbuwJDwxneq1Gim6kV73pcYnLV5SYJm1oLtps3kSXP5UluCtSBtOBaiNG07zweh
o9A3YDXLkkzu4GXFnDS3IOJRSjIEQnI1Xhe7hKoM3Ucz9S35DTqboI2KjmyIQ1ZT5iw26IHQ42lT
Q7Q0wfnuFwtWE/v2AGvX4X2GMEI2mfX20SX9GokPJCl14AP0fOVhYUC4jm81T7G4hgWo5nCAX4oO
jJfM2Spd9MU54gPKDrgp/lcecLpCS1LxOB0kRNUbC7X1ntEzgawmHSwsr/czj70fURTNb0PdZTyx
/RGc/ZnWNEOdrSRND7RHfjvDXo9k+k0G6BBggZ5wrKAUnRu1BVh9c32cm5J3hqH5QXIP64IKblMG
5z6PT+xctUKk71w5Ph3Zo1uUKedhNgrGIZzBvfp569oqf2RUVWDnXueVavA3AdAVZ+Km3yQWs7xG
Acr7Z/eRmRDVBOti0Oa8aUZAcu4EO6l26+5v7WYsFZ0KTGL9FuNxGsryY9sGpEcIS8LIQ/lp/ex0
xjZ60xDpFlp07gHzWID1EMMQXZWnF2aUlWSbHsLTOYtzceBjYTRa+aEHyG68eGSFE6dUY+HuNY1w
V8XD0K0W9Iodswv95I7sBzpPPHGd6AL26Pzc0e1A+OFtKRmlydT8PwUF6l6WrtoUV88WZS1fC9HE
H2R4QaHAePYAgvQ6WftJrSi2gxIaO0jyWk9rrMZ4/l/HUEZg4G9qmjsaACkxZEKo0zedn3Q+PKej
R3gKYzRl39g9uDsGdGKT7vxhEVfT3xMnf3BEp/2k1b/gdEbPRXUtwioMfmP8sfsIfHZq/ka2sNu7
3nAf/HXHXERNuXuNxnusphBKhKSQ0OilLkLd7QPGeCm05PFMTXKCg0DQYxnDLR+esFt7Tw5Zp9FS
juBiHbPIEGcJnNzdIA9V2WUiLux7fxJ1qA/wwbrhkDv7pQ3JF+9H5ac2KO9TrbhLrwY6GGWA1xmU
DPTriOn5quOYiyJj5xNF2wIt76/gFstptsQF19MvVREWs0wkdBzXSw+8Vj4OiV7U2JsRLyX1FBXN
BaK7AxGcTi0n4cNIxRBegJEmOzS4vA5fDcaTLFP1NQlih4zzvQ8m/wgQiL5gUumJIuzDVeQNErxH
4ShrkxNe1snvTkJOuSmI3xRw1qlQXAWDnOprmm72I+TuWnF6683JJOh1dMQZjrXjyyOeW757EzDi
2fMjudYoBTczVCuwyiwnz7W8Q+Xcu2QoyYJDOntvpAcbOP/N9Nae7LJbzBbiQZ1lxVLCWj/DSEV5
7Do9WkE5BEVjJLjbstOEQE7lFzJ9BWnBD6ojwfo1L70iU+O8/nEwIgUZRK/7nPh0EYt5vCMlLqpP
pHre3MATiFjjelmlI8bH7DwT/H3YxxX27FwtaTww+MrELjdSj5TotRyPVtVt82SJPqRRCYgGgDbP
K8g9ZD2GpLRrj8q7ZHcAG+ytXBGNiCuwU3CesllqadtZY/OM/3CcBJh7gKyfSoTfIRf7phUu6W5h
pn3HNYeuQqSR1clp4GRurQFKxgML35Ec9uRN8m2SMhjAamiDu70W1BZ9V4TEd2YLLk7+mfaDxpgo
gWiOm3CkvxNRCMmn4LBYALGu5fHNAXBIvYUhRz7uayFyP5D4sLCDz7toyDVeBERdFmLxFdnS6Z0f
B+cX6jSZCNClMdhPxGHgknee/nghYtSzQK98pI0Sk0WeFwvT9ZZLoHB7Mk5Hwvpb/TvD2aKIawdj
/6XuHiNm8F8qG0qveCOa5XcLGR6sR6vTDW+ZO1O+CBi4RPFeXSG8nWvBtF9r0Y4Ii7/QBaq4vEzG
NBV6y7GnEe9Igtj84uZBzjdIarYy5etiyZILqxHIeKoY9FC36Lkgxr+uXTDkGhV+f1MhYtQk+Nbg
uCv+OZF37PAh3hGo5X5CyPPoq09yBBMF0WR3nsJ1Ab8mbWdjGIQZmHexH+QrFvbY/8qm/GB51IS0
A53IwMFWPHper63xvAO50iBJGMOVNsed3De5jFat9UREJ2Y6bEDg3To8LQa41ezEEu3d2bTQN4as
OhB1zm1/wNWUUOu83Xd36N+mY1kUteikfcSSMIVl2n7uNGhgFreZcczF7dvGLeGsRVDb6vFl248M
xR3UNA+j/3tv34c6DkjJlqtUSM7Y36RWRUiki/QOwUDXIdlHv1ySplZbojDHpkI6zFyguToS7W7T
rL4gILT/nUv8nzWHPJ08cB7lMGM3NMDoTAt5WFj9uMX5QIvmlnYQfA0bWlhsyKOcG6VL2JpmpvBq
+VUIUhPSM0nZBw1Ev0/TOgW1nM2JFkUZN6KjPIMnoQLDyN3dHSmTRphXcKKyem76QuMUjKkELGt2
QRK9xK7PLlhy4cAMMrRGxwkIZg7Qv1JKMUoAZgYYJPvzzkXNqO+xe9nJy9iQUZUry7o+dD0zVzt/
rDOJpAzf4ZjMTDyLN7vKhGD1rp2KSYh7GS0w0Rq9ig7roFZNKeTh0lDbMgGh3DdJRYJz3mh1eKZc
ei12vB1MTvsY9byKGToFaSo2wFFe5fuTKGtznB1QNf9dz+bWVp+sYlH3w4auZrPxmxPf1oyxW6h0
rT9GM5Dc6AjAYbCWnTOhYGvBw85S4TZug//Ef9co7RgRQve22RO7TbPOZEnliMnr3+LwA03zWxY9
1AXxqi6+Aqu8OGVbuTlXyvrUy0Ee9xASWHMmmYWhR4jt3HOhnEV94jFuEo27Lr/oQqmKIW4EgbdH
jyQ9/m30ifmcqK66c0PGcC+1d+98wlQk54LsM8idJoiUdS+vNRS56DzORL5GDhUwfYx+zM5qPW5s
NjOBETEeLFmn+qnHXYBmyudCEmx+dn49ctCFYhQlStjvus8yl+5vB+bpyfb1g6NDv7CKdBDxBpmW
XQxg6UGNDKkN9KTR1JwlMagPesTKHoSgUbVRVwfazjSrQL0KC/6LvLjweqEgCOJ/HUVgkX+k8PFH
2+w8n7XgNgqUNyBSLBxSlUpFWmtrTN8gYWo8o1CbPNH6MxuEoVvejOZiStQYA+HxvnM37QB02kuq
2JLywoJaTEgCWqXq0s+6kHCwn2494pKNokudzCIiDEHCbZYWOsWZ4zxUUoK14Ufl2i4LYX0MHjTi
y08SnfOMZ72L/Hqt9Pf6QzzygmcsUq1G6Tl8/vFCBWbcKNOy/PPc8gXazXlMM7DIPEStZJdpWCtT
TdgOluES5wP7fbgVfuyGlNnd2VmcpnFUxsXqskVFIUztkNxRunuE6Ssu1Bf6eyv9kU5KrT/vMhqB
Ve5TOv6UFXj0p39pFLZpbg6y0oNl0uR8Ogcp3W3ceNusR1EXRdoDSiTKIxx8pGfkcxCnJH0HDB97
AwQbjB9nb/Yh56/vqPsGrC1NBoZwLRuw3TCjvtq7MhqBCuL1R7WjqmNrWkcxXehTpCFFEIie1mrU
Zwklkw48bK7I1Aao3mLsvwNK3lpxS9bjSQ8pIaZyPN0Xai1Am9JTyLpOOdD8kbt9quN7B423DsoR
WyIwyMxlwj2N1mBbIZGdpQx4nDAbIsepJKQMxZqRtP24JHlOOq4EDIKyBCxKp+wuz1QW/eqyvw64
T5mX+JxTO5plmxSeae2iGCbzHKgNc6GKMACCitI4lbHJuyFf/66Ab6Q8jShfA2JRfIa7UsnlUu8F
BlMHJMhr58YvGI3SbttonRH6V82GOYzAnB46GsAIvEXSimYNpSPWcadixxSWmjpDIDXCd4mK4V5D
0f9TcdKeVmOHCw6MWJOHRVKsjqNO3g761AEs0lxEgv9VCKD0aSsCDX7nQYQZLjRZ7BCb+HEn5vHN
fLJI/krNGvdGe5vjzmeKBdGhyjBbzUL/taGbNMeOfoYCUXdnz7w80VHVthVkh+ehy/mDMpWy5rdA
z0wj3CmhWUXbAtsZdygSAlcdod6myQFwCnqg+9AJ0UzoOqSZdpSZ4cqM73ts7/G9EpGz1jRtE3cC
JuFrr6RWie2VMiKphftDQlA61WT2X004kfWvNS4JpvT6AhuIw2XTm1jfw94pfuO8QRVSNVgcSa1X
xlLu1yqqbvMyf3VMrmSjs+7VSKmPfJAQJhS9cw94UCPYIwhKoaY8DxjEV8TQ9juhXGLXIJyy5FgU
2tSJDxyvsF7PQ5BYsIfouGZ4Jl1hIOp4lMcJCwmf9P8s+x5Va5Vx2ZkbL229cRPS3PL3Zw7nX+KA
Vu9GRjimxypBNjo7S4yyRf9u+NkHt4mV3K3YjQ3K92rxWXpyIYl5YQRNuMAux1hqRvS8vnKlgm/m
SCtpTXFoy0Ivre7b3R22LM9PkNNBb7dGD9zqCBbejFWsyqGytQdWIRIttEnV0p8LyeJ0zvCH6zF4
Jets8BtmRn36OPl9UdIuFYEExKcy3xLl4m4byN5xqDyMQQVruGwl30Jn+eJ9o8RDkUQ6jxtoS9i9
1jK44C8Mf3HMFV/AudS1dPb3jL9Bu8jm1hMG30hlCphDqFzJjQPFeq3KOUXXf3N7iZ+DjnmL98/0
7IWzZ4yiKY5l99f8xOGPlprp0EpowCdcy5yRy1dW9KijvDdrUN+HPxVEd3GSUitFpDrO42Gvlq7f
gPsc1ynqU/BuCbdpXFcztuW3+0IApbaYFEejmaeMTIsJ0+c169776GtKFglII/+tVO+xAXfa10Sz
/xOwoBtq84ZFyhjN7DR/k+UWw20MC3PLKKeucLkdMUekFsxqp+nSadx2RpA+HiwNACp52VVISsja
em6rCi2ju/9EEQSvJhG0YLW/R9wdgFTJFqo3NOgWhUy++x/S+5VVldUVVclQFMJpBx5Q5YohavZV
6f/vKBUYqtCINa/St9bhEIkJyU81qtvCFzurFpU0tGGH+Bp7binLctHlsLlhtjVMUg6QXr7sH1Zm
WanVhdk3vKXRBIbj/F5VvgI0Cl8xr5TfvMmKqXfnNRysI6dh5FZgX6sZx856VXLomDCNf8SnhZVh
2uAYqJpVOQohagdD1ubhE2njAocN/7GYqvMAQug77S79LXT7B2WgJUwcXZpMexkkBRBLeM+rFBIF
bjjV+Dk4Nio1S6uzngpGwQQa6j/gg+n42cMFNAgJxkfwtW4D8jkX3aqt8ipXsLma0sMyxsS4GnrS
2Fc0DGcGRcDaE6usOZnPW6c4UQzsLgHHR6ahfeclpRUHt0s6Ta3EkXdJUdAss4Dqlkqzk/nolpD3
ONDly/ALXZqM/uT9PiDjg+YRTWKWOECdWW29wRnWhVqEL2Ctu8iQI0gqY1AC4dWJbFBkQxWss1HZ
2/XA8NKWcIvlzI6anIS1kXckFVuhztlGjIMW44F+KK9iH2OvY2jR1+AR2da+2soeQk6mI0FMFdPo
MO7GfHCue+nArbWTrxupT+U2KZI3TfNF12jH8lnkTC/1x27qWkkFMlb/rdI6HjhJkWAIcWpR9WZ9
bbE2NCrtqHBlHpmotrJaFhfsKHpD4LZH9iTTRHYXr3l/gdteELpb2gdg5afZz1Nf//kugFDAbPyV
hLvYmKt5fHbsnsU0O1L1fI1t1kyGH75lbw5VUXSOgWfD8iuWgPExwB4hLrSIcKZQtWEyN3iUO5WN
5mB89UGQNffDfo1dg3Xz3Yj4bDmHKmMQFHZBhD02ATIPoWn9aupP1J4idWl0mbpDDVVz7uJuBhtQ
rT3rp0gdNZYGbXTlqoIHyFJWp75GFZikQnMkIWRZ4/A6DiMzgCjVK/rciIgrXhwqs1USD8nLYcrV
RuMBPaIi2sbr1Ha9zdDqv3E5IYNsgtot6XWucqi5uPh/IwOPNzKNXxO2G9Y16hQLj2BWGmD0Kzq/
lVYdz+oXZtVBtsjjktKNOdg5F3BMPFcdJrBbCAktrfp1YN4owcC0m3TIIg39Ofeim22KzPAJmTE2
Ktemw1jCaZvvoY3o65T3cr8I+k2URfnXe8eKTT4YyzU6huu093wtCZCc4zEXQF0jhtHQF2Wl5sc+
lnDzJGowpNGibnaycReMjscER34BAJbh79MIXc0uCKq1JSuWisn3fC9USPrw2Ot5MPYkzAs0w1hE
XaCrr4h/NSN/JJlXeHYByqGt5Rou8G2PG8+Pt6brbvB3/2uscV/V7bWcVjyQijs8wQQ+JXRUphO2
8xazsZck+IjMiBWy+zwe9MiP24CvkEG+BlB26ObSmxQ1Kzi3BH9kjFqrOC1wM16+rQaRhe9glG6Z
8TLJ9FtnQ3rXnQQxhi8sdIis4k+0W8y4IaItPyGvBT9yMuDh64DNyacKI3ELUerulykc3PFSzN20
OlD8dbFLlulQ7T7v8M3R4M4r+TeXW7m60wAceAWB8tGua3FD56zYxZvyCNI3zA8awKcEJR6Ey0HU
s9b2ij5fvpCEWZbbbZWqYkhxlk+psOGgFLHQGcseZJ/lzcr4+uFdGNjB539uLQUh8OCvxp2N0TW3
V93/BVZU7LP1GkgZWCno4s1gegcsXak7XKZxZgDKkEcY9D3wzW6GX0wXdRhIO6L8fbI7jArU9GWK
73nJ7pOCxc/Kk9ydxru0XiXDrFvWeUNo7+OLhG8yLV6e9qYtjW6RCiwSH3qkLxtNJt5qg849NydE
lq3Ty2RSU2DFyDVRVQqqkqDig/C1x0owsYIyJ4vEMPqAl/AgPhcF77dwGtgNd3nrTkSNQwj47inI
O9/BcZPjnRfqS2EeOf+wItMq8oYK54uzNhUKhEwTcnJGcoC8J3igSGBf2tcnntGg6IfnWWwhX6LG
e3d6OQ3OLrkCwNYDU4KQWzBbQxvAWSHRIPWy+DS5iauT6KGo9p8iCvrg+D9JxGKaN0JOiq1mNvcl
IKmn5vFZQ3bG/pqxg2W831sALosLCJehpgMZ35q71qFexZk22ej9I2YxJPdTxgMk+VDzQzvxwsSd
7ROcuHDKTO5WynlLlLcPR62CFIgpjL7DrMrrQ8FxxFqK6QSKxzV6jXKSbF799eEEH5vN8R8B4K9W
mh5NpF43/S2+xiSBBzM92HkgNbI6iPIJGyqlCupQCsWmn5X/GsIxu0vnfIetyohBg1FxkHWUe84U
UgEfGbx1Q6VyZd/5BdcdgB5uX7YA6m8vRqnuX8HMPolSNB0r27PrYwzMoTEC+mX1l3iPqCL9ejt8
9oT8tQZb7f2HZfg7dXFlpB4pyEd9U6s7aqb+smfd0WgwdhEog7AlL2gl4mTFZBKo/BoYHYNIHkcB
Gv+IgOesulTf+YDvi3dGO+d9yrqq5yp410HKsa/aLKCmrEXMTm1RrWts5o7cB9RClbEj1rxP44mM
x0UDI2spaxqOltAu11kaKRE06Vke+HDTwxYQEAZaDO2eufGf+4ekXCXWVn1FlZsx2mt+zKrYEfuH
coxqH+Tw0rHeeiCNAggUg/VnOf+g5gkmaM9n6jVlJmpwXZwtsjVokb+oFfFSkiBYZWGbYPv6lI4T
pnkz10Q+3d0LQ9B+wBXaUtNVWKkm7IuOY6OyoP5YRJMhvqbumkPMpMBhWcjWpDiLfV6AJ5st0JgS
zFUWQl59Rw9VrCw64TWkaJYXdtIe5/Ow9PAWBc40U8r1bwuRkr0KeiMimWcIt6Ca5RJKZx9Yl2Qa
Wys9n3HBeybLEBvMOe8rBArYxeLsCxZMdEIYNGINlHZGHgyUoRf0klawZEMnTsofw2vqu5lx7W+R
wJrgMh2hQNaSmE3klhaP7EcAYr3Ok6VHDh+bVfJvX7/gsvhaLwzZ0okJKbXixCbuS3Qn077Py5Yx
u+3RcgiSRfzaZZrZGoof6WezcFDYFickjxyO+bUFRQ/XBd4k0JERcYLccPniJLK/7CIXxf+f6mS+
YZVfhWsAGGCq6wYlHTE1iN8ZxhUa+StSqXI4ADQoYe9Xj/ZgDWqkU0h8lpcpjOGuQvJCqhfYV9bo
MBah4YiLK+5gVu5YAe4hxTHJEBeKxXZGK/dgp9wj351iNWONOCY1HMRWt5IUnV9pwENkvtlYZLAc
2eQj300wXGqplZy4xcQhJXfXtC6wzt3hGyVPGezHOp5CX2jfUs/V1n+H33RnB6+5PzAJ1YNqDECA
A21g3tGgTd1L+dQISJsD6DxD65zzEkXsngzj/PE0yLLnm6l78fhxFxNJgpdy0vvzreMP6rfAPiZ5
aN+fAIFA7KfVc60nF3f08bGnj8qZ14Cp6uaWi0tqqvgL8IQGZOJYGuUKTnN0NF2EjRN0Cy1endbO
NIHlEghJG3Zmg5JQIoqfppspO9YzxRJHYPcoK0myso1cBoGYmhv1GuVFQD6IZtBCbmpgm4yjh2cH
NPyZrvQVPsuoB4lvVNOoK2wECwuC0JSrNYiJrsMIsI6rFTVmZiE+Sn3QoaXsQePBuLIDm3HaqvT3
tpHXhryJ2MHSRGNMCzxG2hTeEfVgQnrCo68mqHyW8IpqC8js7q4MjVVPzLdFx0icXbcMoMrPB1n5
St1MM6grohIV8sb9FErhdmrtmFZorBe609zr1viJcVFTGY+wuSv3vnasZ7kmPGnmPpF+H3psYQFv
ogFwlQTrFc7Ly9eIbuJeOF+xe6dT2zd5wgDYMo7azSlxpOumbT3NC9Zwo1hyj8H0b42VXqTmTA9G
rJhKQ94pHgBN6BgqcGfCKe39vUV/7iWlUDi2ua/YLmkP/Bp+FG+2YwPSaSR0tkpbwvWG67C4LtDo
vs3WjWrwHWw0+VJLl795kqL9rQld90M9C6KPardGxVFQyCO6otWxG8XiFzY0sQji38/m8rvak5CY
twal0cJUX8Jq5qZ4K2D6kw34Fb6RKqC6CAbkFVrR4jV0QhWIVeGEWIKR62nYIDjrwGvphv5+AZPq
mHqZxx/ne0U40xMwA4bRxFIIYp97BhMrNxrGWQXKGnqiOhDffmXfrjA/JyzAvuJgonMz63sbpMv2
ldee0naY+wki0cZn3NmtFqj/giZJmb2sFZjKde7MmOyH4KT4gldaNkmdinVyZrOHKF7234G8ePAa
Y47xr5tRCWbiIdu/bOkpniZb33lmSV9HtfP1h1NaqGZ6L35Ols4O0DmDyU9Zy+3zCBor4K+RVHJI
hIsLClkm9iju87IY/uaJXcFdOv/MsJwo79VJ0Qo0sivQj8/jUyJMTOOmPa0mSvoKUPS18KOPhWU7
CflXp/N1B3KYmvQqXC5ON7jE4t20rsz9tXxC2okOZF2pYurDOoogSgR+6vLEzM+Gu08iCiovRrs0
DHrFXPEuxcPWoSPNN+YUygoLfl2KTSjNdG7zbJlPVYwO1jwhyY91weReL3q9XlIkE7yk8t3exPWF
32ib7vZuW+yYwczId+C+F+stV20lXjNJ0ErmHkfwuLnQG+StfIlpk179y82Gyw4Js3lddUffNYrL
lPe15/cYVlPhfdq5HELjz3O7l96EJmG0ZMKgsMfQ95s8vhK0d0mIRoBEoqGYmAtN4vKXotaScF0H
Z9y4+CBuHBbDMjgydWNX+CYreFib9ifCPLdkv+EFoMwYhPjtf6gvyzUO7XT6PHRNltOTP3MK4n3k
rXDwRBnx0gE2uNaKGfH6EtcSlcpf9kN4mTrTsYnMr29NS8ghl+5JfFo+fWdYpBJnliP0kH/S3K/Q
XDZ5SJbJwTMP0m1qSyCW/7kg1qb4TnLTydnNvVeLQAuvquQpAMRSwH97dPpcjhtCocY0AszS5V98
1JbJyToUOoSRNRcj0dVN94hX9VItbV6sxCcovikB6bYnTUF6T/mtnAM328RTW1j4sWyf13KHVTmi
XmCRQEgSAYUULfvfuSPUlqt/M21qv2EGDWSegHcQpcFOILGdOcmuv9ehgSUBj40Go9gvHid8Q2XN
7S0BxbxRnRdjQscS9EJrEakWN04hVWeOJcIgQFE5Bwg5QGL6B45Q99h8nhgpyVdSuokFEaXswmuM
xDGjcZzN9w96S9mW9NcKWeQV3OujQgtRQyM3Nd4Pv9Uy5vTPps1/Jf64E43kUbNqjsbuk84hWvm5
7/zmf6MdfxuB1TnVojls+hUp+dgKa0JJntzG1iXQiVcZ+ABBIwZmEFGKuegDNRXmz/iZAAPZkLo+
GhAFSYDJEQ46syWAEPzQF2WsWLupjREDlampnu281JNXHeJeAywhQRDDiZMsiJoFQ9b478hehckQ
1gd/6omhK6U39zngexEtR2F6Lx9K44i9FcyTw+/MQxMxcOrSk1Vb32Xd5KRLjiN/a5nBA246OSFp
5XgA9EiMl9YCSwHdLfXGcCeI+9OzXsujXYrQTjRvYRA6Scd7IlgQN6BcxUYy2Qx00IH63Evpj9lJ
i0ZJbUUEDzxgLwurQ/pBL8OQLgr2eNallBxm5kz7BJ79CkUB1R1+VIuMnWFBm2SNypRpoVdMdZ1t
ggum1Y0R5aRc0mRI01TMQEJVdI47VevfpTiDgSRVIoBn3QY4Lc2uDm3FKTRKNN0Yv2DsZA+OPhOf
6Let26E8wCZNkQdHvCxeqmrHTDsD6eB6dicrO4ZKyDmx5hN8HkEXnE85WgFxYg5cB79190IKo0zg
6SQWKz4jICx6eX+Dq4hLN0IfU4am22uBidXWWVFIFhpCG1K5cg2KgL1WtMhL65uGn4mLwe1/93yn
LTS2z+/GHQRbUxfVkWARZY9DWXDLL2LIFQeV7hIDsP7Sx8M1533jsxsnTbg5K26ybIPfq6o/PjuL
3JX7Qn294aXn4IqSLsTjVuStqHNZigrIi3BXipyrYCOY5OiYebGMCwnaXdc/O3P7KVOmaQ3BxVm7
Qdk8tv6NbZ76YPbPMu02thQqFv5JJesuFu4KfKXzHU1OqNnzosLS81sQqh8db7svltHxKbkkXqMS
M3iiZVKG6m0OA0ZuYjOp3uUpQv/ZvaloEc2Xuq/wo9QK+QB9A6xCeAvHDtQZUW9KSAe6l+i8/ziV
IpOUYeF/wJafBU3WOUusc7NDttfaV0csD7yAuWzHfmtmtfDH94Q9sWlXHsqtIkKgBuMmXAtlY+ZB
bBwqb3+yjxsRthGUl7Hs1kXvydBX7euyUwer1OwN3I7zxuTiztiBqy9VVirbsMt4qrgBpWKbEfkr
cgH2FhxxsdK+m92embe4GdSYGO5zcD5I6ZkluFg/lUhom/p4MgTB9KJm13jfG5BOw006R2o/TFIO
4EWg0I4cGNQ+ogQCPSbeNnlOAGHAS4Gm7mwSZXUucSnIn0ICxch2fL60S0eTgvLIitbhXRMXkl1d
IGgCewCnRobqQxDlNPP81ZW3BMCPg6YoJyHlj5Asx/mYuiAXw1Yb2WjSXBYsGkDHbGWYFQlKerCI
NeQKydauAM0jatv6NgIoeszOwCnUJaJ2q3U4BgQgc5zsGdxHqGt/wl9cTvd3u3Sv5YXZRnkpNNA1
F4U+NxjVT8+Qj24By+AZFKDQJd3+908UvsFAdn+OQRtPcKS6qKTP4+xA0U4UzVkLTYKxInWCjq7v
GuwbM4NL6qGrWAYC5FK1ei1RuMFe/jnu1QibsmYcWqtZ88qc7KRWrnO5iniar6ESHiTyNYD56la6
AsJhfNKv+pSmGHWy4gfKWPlTpTNCw1IzSbsXyWL+MjFd+dPQ9Vmmxi9aF/LK7wQOxWv6bg69DAJX
xRc5gfiNh8PmrkCnNi7LUi/TKeHMWECzC4bod394OHJMouvMSMdCfWL6upmARoH/4ssJGmFGZAPw
bCh8pcOH6zBjgTjci4PPYr1dCy7619Dskf2CpPospRIReLyWfX43uD/KaYHmOaAv1bGDhXrURyRO
NXn2xkPh4dMFfrdK1L/IgC59lrYQC1C3GZIpbj+vJ988hUTNkGc6wJkV4FXSuWMtWycx3njkq5Am
Vjb/8NmAdbhZQ4ec87iekJfsyzH2uiy+ucxnAc41RmA8wvEhB/QClvPzZLDVTD7datOtIBE0cTGe
Z0FYIaljULXN/8OPfGLi2lPVefXgwH4B8wguuiZbjTPziYuWAmdWLEnn4GcZQvvhtfDoxQcVmxp7
y8fLVozE7HRHvJcsCQg+e8ahl3M2axdu3wgUlYgJB4oBmVoZrZUu2t5A+17JaND1b2zBI0djOYR/
M382RXOun3UBylMz709DKwt2itAIzenvM4VXJnRyTzckgcGlcgj4QFG9G1kiXC4GcfQrRfk7X6jL
dEMqmH92+EhAWYRAam9ShHvEsD4FWhKAhbYu0zauPnYzQF0qLabhcemy9bgkXpTdJ+9NxaFK3lSJ
Gb53GGtL/RIBDQYELZE6iiYC05SgJiDNtoHf7orZHnK5YBDTYfJfci+PGsrIyvGzaTwSiuyZHeXw
GTbY//Ludwya1AJyFNHUZW9keGF16GFbLczftEoz9k8L53SMtu2JZPimGxquzFnNRw8F++3CVIZ0
r0fuuAWUphPqKTwMaSTs4zRzfvXOM3mLbcYYJKGK3RZBsETtEopVwz6/qyCFXQ277uXfXD+yfk+N
pqzSYT2TKqBauupWE1MWAUkCuuo9xC3809QAfX35/6IxnQXorc6l6fr1EP5n8moep4rAESUNPgU3
0seQXQFUaSmXU2w5NYlKkdqs4DIagU+ObKw2t4flcxJoVtrFB0JDiD2C3uwrzvWZsVCakp59GypT
9Kq0NLSHMTsrPmLB8lP4RoYDJSkEoWr2OOp9j6DlVcl0CbK1mdaGGhs1SBo2QbZOeYZ1mvviq71E
/3wcx44rIXo2jv8PQgfHyyodVAUbH/3jemU+1XFiIAGf8DNJkXr3glk/wnL3g8HTImGhbX/vdkBo
yeQrF4JnZG0nlJ7Zav7N4h5SCuDQeViCMvRI9KJuqvCrpAj72/s0+SBQUeVKZpdMrou3ugRMWvvh
UiX1dhwlpbI85rfEb4r1xQAotLZeaajxWdbC1xVria/26P11tRuGUIOnm8Bz4eKkEw/LZS5onSQQ
jB7ZaXxIuC6YKqmbvvoYaw6cdlubPs0T2ocE5cghmMra4nLsV1nG8DlK0MFTxOhZB6XZ0ez4+piO
st7y0N4kRlgdMwM6pMlI0Y23R8vmCMvZZ7fmRLgjnzKhrn9q4wrrEYp8dAy7+xwMVsSLxF6Twibn
l4xgcuPMhA+d1G16kCKqyWhpQTmLMkXEowT4ICjIOO/Vx+HNfOqgZSpJmup+UC8VX40WhdKMtKu5
mY+NmRpjNeoRXW/NmJiNHsLJb7+o0+WkaWfdcLWYcX1N/JSxoCwltDkyIdvtCDskdaJ3hCZ0mduf
6D1l/DZr0ERHvchuGhY8yBG6V/zc9xjb/FD7peRAWzuvMIWYLmay/Xj/Ox+AIk1dQDy02/XvCZYz
kfEpGv3KA3020S1RIc/RKVlclneSvSdiQTl5BV1bMKV0f60IZ91zCTrkt1VHQfHPvV3sUaZkcxaK
tY/OUXXwdffP/DwifIFmv8Pkfn9hvtMIWbsTAycqgnqz06tBwCy2neMndHSO/z71BF/ztZx/zfiw
ufT+IaZAfzXjJ/SNpWCQLDTAeSQNI7sqghEUlh4AVq6wCc8YVyfuC8+ySDQK58cwtlLzQOW97GGw
yyS9IrgR0CebYeJfG/eP/lX8xVWy+Su5FXYzr1AIu5Y3WaI0hvQUII8HHfCwQYm1cGNfBkWd+p+K
WjIul9Qjzf+BzwIyvsnzIFSJkViTMg5sOlqRHBCX/MX45E4KRMHsr+qM4ZAbn6/8IselKQbidKao
p/ewzvQ5SbC2btMv+88SCDjwG+K+GlW8yPCreMWZE9KICQMkHQiM0QomdZlDt9/Wbst6mM/iOqZi
H0cGLEgr5eHkNJ9UoWNmSzO+ONVfDeqN1BEleQS5NASh4rDLilT40c05C9GmA2iUWY6R+lilhrid
SjvN2CsV5daFO69Hhm+K+hTj+QgFzDavnPMpc4GtOHNOovJO+U8fOvdeT46+ODg1YD/jDmRYsCSw
+A9TGRtIEsw05uORg2GC3yUsJqnAxVjSaXxM5Kij8HTk6KV76b3crxPDsxwf9dJ4ccuUdwCgWLUF
cNIiEu+x+bh2OUxNwvMjqYRpb/S+L3Wi2keTbYshXoURkqjk5ks6ERRtr9EybKoxLocNOs1KgZQU
ojuHcLTVFqjIocYizs2BwVes6SWgAjEYtb3VEjZ1jFnSSeATJe2dK6I5NwGiHCSyMSF/H+I+V/R6
8ygmxwu6MIZRYsKQtF0cCrCf5lWGHIuueDaSpTPD2W5w/SLgySsUFtsK/p0+VR39Y4s7kZYvU6Yj
IcfdvGIwvxNHIloR3ufZeqq3BIyRmVfCq+4bjzDqbHYI5Z9GTWo/g//SsDmWSAw37nFUnJL4+/NC
3w+XjYI8P1jJ+KPPcBE7RmRP1NO5zpHojSoCjASWqdaaflFTf20+mOk2klY8Q18bX2G7+VfIn8uF
HjKAbNotSjnKg1XNN+5XR35E3OprElLKKMi3R2TtB/nDS0K1Ol+fdn0GKFoTDaJG1SZd5SAlERGn
JUlIfvUJGUVBoKhF0WINK3IOJQUC7PiJm9ZmQX0mh0TNjyD2iJOOoxgiFb7zpM54TIMliG7T6F0y
F45XSMBCuAU6mWXeo1W8N9yLDIN1iIHE7AyVQ42qK+a21eniZNVMZbqmDa0hD50J6IWO05E5Yo38
dr0iN62JyRf6YWobWVN6WM+Nkf+FoQ/eBKkQBTJYJ2HOS5m1YjiMIvuJxL+zQM+y8ZSr6Lh2wjD1
EtUuNaPkepapOzTI9o3TBy5eAaKbDVGTFHUFRNYxKt/eiDQ4MAHsVyyDkfHpyIXeUcN+diCWeDd0
EunmcLZ9/TJPD3jGxLUUVz80Wq8wX3J52YQgryRKTwOAGJYFKm1Ecf0OXyed8KZzf4vrjnBah7cw
kZGOChgNr+De4mCVBszehSl/zkCtIVx78Ycwakoy3cEO1Y6hASIhQ9MFDm3lFVcwMRQ5A6MmOGHS
xGbQ5mOQU70LS7GpuCyDmc05WYqgMX6QYLxX8g2vXvXHT9lZG/gMAojQXzyVe7swNK+nZ8/bLtq1
7cnwoFrF2evKhDiMY6PaPDp+9ZWuSZ8ziKvn8tAodcznQ8jqbk1XrxXUlPgJT21ba5H7UjBWNT3A
aai4PCXMp/6RkPdVpPE7vVno+FlgjpTa/c7/yj9dHayytrc5ffx3R2ZIjEqVmSl3VEdWaBbtGlmL
KWnMTBi4j782PiZ6oD17KaMDcPwsY7vRTCbjr7HghAcGD060ZHVgNdnEMKRYVCCqCxr+RQ49gebI
1qxZSefXbQTp9BSGFRs3N/tc9WC8pLY808Sn+TnJ9yRQ8HRcs4jVwAH+ogXr4KLqphHPrWNGZKM1
0qAcEUJ8W86nbDlmmb5B0tW4g/yUoGikjI+yrwPpdvlAGTjSEJXW1O3idswLF/XXZL2oOzhJoHKv
cQ5SDzzxW7v6Cv5tQUBK7SNjsb/Y+23cfvEbrAWUPhbgo+S7Wm4Cx+lfAd35NFUTwH2twfM3V7t3
gBtWgt39jMuQs7bxrHXLX0UyYxRgkQ2l8PYLpIisnA8rjWA78d8dH/eoC6HhZxyKtTH0gHfzCo66
BB4mo0GQ5o0NigFy6qrQsVM7nJa/GqpRroeePQZQ+7ybnGzJCHISivtOtKISK0NTfjK6Xlq5by14
zsSdx0jHdSWtOIxvxTES3A2D2X6f8ScCxUw/3cp87CMXwbuaso4i/pX4hB6yLGnBHz4560H9QJUA
wIVHHGvJFd73RMOxAcpZiuhCj2hWBhJXhCEJ5kzZSqKjyhMAMaTD8fzuKvpvMIMXYrfWl68quldj
PfFya0SQp2EUDPpswlykRKI/EEdOObZVeXf0W4xitWB5RYn+B2c6Mo/Hntze0sj9ogRM5foUXRHS
EcdtQH2Or7LpTp9o4a1oytEXJPWMO7ITD4URcI7sfUFL87gbr4+9dN+9TU5jSGHN+UlG73JdrRCv
QVUjfE9pjFb01dYsDU89imh6x2VpfcXyuhjRwfHl6IcCqDVntz2/+3JVFyoY2Q1Hw1RfSHXFt02B
DkDSqAtuATP0RjdCIMPZDVR+JbpBowPH4CXBlGz38q42R/LAlEKKKC9GWUyh9MtR9uK+Aymirdj9
tZFWXCsFymYWuNWUKeeqmk0/GqbPH/D+18CJeB5VB47Lq4S1mIAHgWlZV7ngmosndUGReoP+RDuQ
GJDNiNbGtOxyoWrklG6duId4L1MJ+8Nbq0zc952izDOwoZ1o6sEAmN30Rj/6o173EYBzzy081As/
YPzHgQXPlrvs3pLAjYa5vZVmAXxzKqKZCtCYdKFcVZBc0vpYfwCB5BkKfJ6N0ZALbeR+QMHYDvTS
nxKqKOyyZPoHEuHl41ArLKJsXVt5EQK9LZ3uUOKEPqzVf6Eo5K6KbbUpKIUHtKSYVOuO2Qwwqv5e
xxQfi+zVL9vKCGeCADxROx88BGvyQVA3XkOyB22DwHaEYNfkEycybcJQFPOctseKI+7KOy9vnLuR
svTf0HXGqKLhOPq16oulxYwi+h2b69TAHWfHt2BrbNX2FVgj9OMxE47qks4yySB0P+Ru4TA/UBAy
unV47BaICNAt26FnVZD7uIO3LfdZXyUoh9IAVRYZ85IGq4Pd4UtKG7o5OqCYav6Po6lZ6Ze/ulSf
ObaW/YvHzlICuFOLLCA31WoKL77a1fqGpEQlCwHzD/YfieOAOkrn5KSwyyUXUTi604VBYWOyJA+J
SB1mSmVKIQmdrJu0iOFCZlMBA/PDeCw55xLs3zDl6c7OKcm7N7ja2b21+a7MhQ+hiCR783fVXm09
FqG9+1UMvy6JkET5aIDt7/RF70uh4YcKqipeXKut9jidFl1cr7uYqS6Cz6UcsGjWJJ67tcMhN7YN
91Mjj9w/+vU02mudbj4Up8Iu6TvFngdXc+61+OwQFMI7Zi9PEP0voP8aN6XVm59QOabrq0yOEJDa
xD9ZRfoS4I8ibevTCzs1Lo294KAx+03nx0V04OGjerN6pcXRCdFoim/wC+kj76j30XbexZylPz2o
mjQEouosgXFG5GbvoCMiOfFgkwyzQTe82zym0gbDOxJJiekMv2jUJIkx47xDHDVgfqn+wSxeLnHh
S2JnbwcBTLfkfDZOGoZ5QiefImnU7w4/MNDtTjqsZIL8XhGwJHq2HdwVwrTFz/P4J05FwEbnMEDq
IJ5GM7bElwYUirx6L6YmewVLEpISMDtiyjkME53bsBn/Xwe8jzTVZtCJufbM3D2M8faYwyiY5RkD
gb7eWGkYXoKYiFv6bE/9H9cBNijy1Uqvmc3aaB3MEW2cGha8ucZ4vWw7U9zlvQ9rleDPPV/K4aAW
ruVlxKImbxAaGqB1aO50hTN1SWSGq9u4iVEG3XJnw8bMeOYWGKFZfbR7Y/EU8tvTC+rv+XkBjv/n
FQzA+FfJieDug7v0hVHZnCjtzKxrFwfSP4ytntWFlfXOHAHTc609FstJWCeG5Qyx6gZ8fKQvf/Ev
ljtFz3JMf1q0q9tMh4dXHim2PK7Rdkj4PH/nWqjoH3g+yjdEFlHsYxlqiu+yWHxIgOkGc5lBmcKF
uTKEKgNsoGhY2ZuXWWpoXFck31gl57ewZZplLVs9n/PWRQTLyG5Uluqfjf5TD5eadNQ0ROcelFBL
QIw38QLpZfVynvLxWtC5/4XX6YeGjlxfqaZfWbwVUEwMgSWaY0AG85DYNJ1r0LaSlDP2e5U7RTb7
2FuWkg2BVxKd7zNNJBm+tbn3sOl+OvUf7noEk6c5P9h3BqRneh8y3R9L3WcepEZqNrg/9ljTUJiN
6qRLNUCLAxz6qqCC3WdOru2LlYYAaLo+gLYZwy9qML/bBAaD4QAnSqF+Sje5p9nPbmS+EyqGb/gz
EHvJQkcTMUL62/hOsaGt7Yb+xkY24Y52paf8UUTt+ZxgwXoHcKqsdbhU+vi/G/lL6sacSHla+mya
RDxasyvh0zbxLb+wf5itewW9Uf13qY6W/TPKlb/Wa+hFCg5D6W/JODp49Z/KMkuftIm9GB949scB
odOWxcWNZc5ixkIbwkBrsGoY4EVOzmg5RuqQB59P6cX8FWRKbt6qgJn6V4ULhBmV1iukmPGsT+tH
NfUofSZ3MXxWb/QY9oBZEXzL9hc0XpNR4rrwqDx3XMC3RlgP3Kv5vBl5w6V4+ZQorw+YP/STy2zS
M4Ftmqh48TNEa6MsmcUJ0pomfdZPRfWJumc2ku7D8G3H87Bm7wdrdja2sfbV2awfTScQPcXlSpvM
DYgVX0ZwDecHweLRGPgEBkuevkVLO9VAh5hKAxZb/A5IneGM3xU0Fo1toEJRJAcjV+zIy792lrrb
rulxqZEzUZxaqH/zJrYIo+jZnhxgIikigjic9za3HU88LDAm0OSJhm/uE33e7nWwMQQvVXCbXT/U
nCCe8skLf5XgK17ZyA6wr3a0xZgxVT6/77WfekxNs0Wgqach1GoEkB+DmFvuByckLwaro0y5xs99
qkUvLwK2mwayi8iPccCO637PwSppnLHdDg3Qos/0wjjv575QTSltwfuqcrhj/XEKidsXXP5ejjFk
Q+ZK0X+cWWgUWY2Td9gGr4orX2YSsR+muZJSHzkPUUwQqRX84dyVi0HioF8nIdvnQUcoPy3tQGHL
lNngf0W/2Pqy/QPNabxvVOSTbYOaSl0pxSk50uSBDSqpk3NRH9M3BfSqRmbN9GsjnaI1ww2GlyJK
ILNzPkNdgrq0DQbJzY2dciYbGHTjGSaS1520DIcH+vRk0DbrONeTq9BA0P3q36dwHNQjyu/qJEZ2
06EavU49eKEuYxiLnSdvQDddnyj5vZRM3e/ulx4BDst/YHf/YfkeKKeMmvVD5LfjY4BRaHg2niFR
/vFMDpITvmSaLCYYZEfr3t04j/O5rKsWU5Elpvc7sTfxKTS20Awf7WBTSUaibCv9hXuoiyepSS6t
TuSiELyna3wX8rps8hV2rdCqrb02/pQtRUaFt5ZTeY6L3itvrkKkyYZ+1tLTJDVfKnpmKXhPa1IO
vcjvqQ/8dB9IdikySPhBvp8Mi0pYWtupnSwPwayzA9MeDB8+1UdcbqFGWddTu42+7aSKaUPmlPF2
P+BV75iiHnPZv4jSNkDdYRknYUcfHoRCmjptzLg/+wPyOCs/UhEDUP4xDB5pJj+gmkzYGMUYL+zR
xlR0z4lWw/dSnMc16IFFUFhcPBz/Tj66IZXKQWWpfpO4C6KZrgyQ3pOXDqwt53fOEYkuRTtIYoH7
2udmi9EZll6DoSlHi+jO6uSUyubHku1Zwl+Yixq10IZYdK2H47gegNFWaxJqM+eUK0UBCgSgDFUX
GhVwVFwOpPz4fCHTVTJ1epJG8FsH6dJHSRgoF7jmnadaAzV62tT6A2lYYRWmkf7bEUzjV0oAyADb
Yjc0NPhG30Z/fucKyc9J4d7zUmgfBPpdHTs758Wy3eiRdrMO7+R4DcqSpOQhZ+o7CJdi/FCjIZ3+
ty2H5/g1fRAMmay0oEZuB+lV67DIDUO9LiaYCQi8U7bLTf3g0dccZQX3CrLzVo/gXN2Pe1AtsPIU
FVWbyiyyKrKtkZMNwFMVJq9JMNEbgGBXxs8gEsuKfx5twINjigsYMFco8cNeb5CKHxJtzsA81B4y
ZrgKQKGN8jfN9KFKA+zeltm2Cd7894F5j+EktQEotVxVARxqOOVSTuFgXp8GVbGdmHUuzz10Ke+1
geMdH2c6h+uqKijkEWseaHapNVYXRzTbKej5ZilFn0ridJthjhlKgL69g0fMUhMKaT4qSZSzXnHV
NxF5qHWshyO6CXrV+jgZ36KhRJmK79FxdYW4DpJjdFwA3atkn/y523hvF2iBOHzIOMHPrSMjLknK
tUG5Lxz/FdoG+AJDRpMhksH06WwHGvHugpvxJmVT/55702uipcuj19S61Hd7ysk/j6ms/nVbqXgc
pJFp/Ld59kG8GxniA6S6wLX9+ojh0Rg/NjlRyVt2JTQI6obeGbfU0hxGbAMlXzipaKhzYwRfqq3i
ISD2mbnEePKJgGAQQCjRqp2ZX+eBrzBmoIpHssYre1q6zqFWNQqCQfI+9DQPWgGz1tLWAVAhJq99
3IVkbcRMU9p8l8UJTwVtNGrZ7MzTfMbjIE2M2+QzWZVr1aRoH2smcP//TJJVfb//JvRC9VyFBab+
vdnD7lUfuzEczFI69qnVe4h+DmHBC8+dcpLwHPqLUXUVUgcNgy+NoJTPLJE/cAqO1U3uL1Da60Ou
1iW3nGsCsIQF9DxDB9YPsYwKj7uH3WpfKOu5CwLhVN1GK6tMx0s/l+nWoN5zuEpkpuT6fTg/RSns
w2v9yIjYiVv3+NVRXaB+eKLQuXc2OnZ203ZMcxQn3TlG++ppUw9FsWwS3f9tCAkzUPhfogQKGJYC
oibuYQsu8ok4hok7OZZ1xkl2VwLB1GRgPXs+XorB1yrmZvlEntUY59wEHpCcArrU+SZ60qID9Exa
DFz+OedRZFJyTW0gDtg+NJEQpfrNmSrZFg3vUnPEClrl6q5HTAPaaa8zwCc+j0Xkq27h/pTrJYwO
pYob5WoY/SO7zDrovW9ZAFWe/XxVqjUIOyLOmFrtv+Q/MWXopY8UNk+q4MJ+yLvWa2L5gEDmeEHX
VBdj4IPqTpFI0dz526gaBxtWyztlj3AJ0wNC5JMxISvuq9tM+D4u6J8U0PXoKtDzsV/jzzpb52Cj
d+zrFjW4jI0cTAHcdW1w+73co4/eSjZmyJdnhdx6tXIbIoQa5CaDA+J/aHwVybamkckAB4hf7Jko
XAQgIZsccsW20InlgAO66I6bdY/e5cIPZ3VWsZd+tozqgFii36FeQ8yIsneOKbEIsshr47owt48n
elvodnuixPZosDXa7P/F/hBBGz7ppq36IwwCVDOjx4h9BxKQR6BRN+8+mFrAIegV9qdy1tV1an3r
EYwU/HKnQgT8chF/DZbYPGRR4kguSIBoQSWTMdad3r5zaIhPg80s502n9yxdO46g2jOXBYoH0OEv
L4PFnaiy7CdJLiogr2dxTI1WL7on4rO1qe/v3l2yttCjfMxB588z3h4rdvCRm5sxK6RJlFztSohA
WgW2ZRvpYkoqH39FeEKRUhBLmu6g46xXXeyWAXQBvD/RYXm43WdS/+KR9VAmmfznYURsup5ZyLsX
KXCNKFwzqNwPosHXL1bhmZNY/PxnnrZK2Dg+pl1UdTUyRfH+cmAAscsIP3GQ7oVG9etHRVI6frZd
KYlzwb8QCCpXh/WGSIP4bpk2aydf/xbch3pRVCn9EFKwgtqO0JivWYEopzAyjXwuHg8spC9aKHrG
otXLH5eTZNFerhG1p0W/ABMeASz9ETYYiP1n/sHTms9V4sZCZGP4pN4eQIvNedUZK5mQ3SLIvfIK
KNYLU9NJswWTh5aDL6JuaxkOJaDuZsNQQSLQKvDiOdTCOwSiWhnqKsxlkQL0+uGyIjsSASLtTZVE
HZqjqqOJeBzhwh+FAvzHM6xALBQEcoTy/Q3NLu2K0mSCENFKbaLU3ImsTpW/RKUy8MmyeEybOOwP
85Wn/7XhP9n3u1yRaWV1NZFLCZcw5dZ4RznT0AnT7ZWS6VU9/FrNMttM8j2fXLrPIVtcf9LFlEle
ovtWrezQgKv25hl4qKStl+VZiHrkRhFD4GFFRaUZ45jTq1ZOA8OVRUHFEftX+Ata5rNQYxiATujS
qcjABY4lVt2eS3vwyFaYPrQtjTIrbcwG4ChutqnQfd4Fi9NlRuZdkd8h1ktrTyLw7kS+MHVFndIN
12/cx+Cxw+l60+lhERqZx5hgPbmHBiK3Mzr+5dsNQXQFPUgAVq89sNOI756CpZlH6zp89ql8ut+7
S+g9pv+j+BFbHmOVkPEoe6hHbW+buSEI3jHgp3ZRUF5vjc7QpzyzU4Vm00/386ZpPIYM+qh6ZZOy
7kENU5dec+oe5Lwu2VmFmuf0+BLvQ6l+AZzYIaDyEHhMKdl7cXCJX0+h8MQWTE0fkjY6wUuOMi8I
J7vW+c/1cL8ZE/7dviWCpVG/sxFCDdUzgXjFArlqzPBlH20DNB9pnWgksCzrvkVDdUJW19KAGpRK
4G7B+ZfJtx12qWPeqtBDBpgvHvEHl/QKzMGHDH1vfVc8v9AL1+YxUi2ffAYrI7t2TPnht3kvgDKA
tf1BI0GYpXxlWzRor8k91gpemz4jL2Ud9oZw4QrBIhJ82+a19XARkDthhSrHpi/pPSXPoyLXwrO6
QwGAVuEga3SUGH8zDVkp7o8jA4+fj99I44tWfd+xQpMSK7uHYuZxIVPt6pO1LThhADn7As1jVOw9
7kG3ufKEcMz2XgzYKDyWdyU2K521Y8QjzRTSw1p2nmNEBTQ9UQy3OYbK/PZxM7zJ5mQsY+772Cn5
eeACnGlfu8cQuFJ+bTttwAM8zWzsEeM+H4BR0uOGES14YhzaEfa8DON+0EhIfZIqZkRy3vGZe5Yq
zpN+vO0+Bz04FPbx2CY2/ANCPKMG/fBiFt3dvcH9aWcsLIQJtKkgbTC2T/tQjRScI7M1bx5D+vMH
FilTd6dfLyJEDCclNw+6PyP0eo9FPj2hf9uAaX3cy/MrMXjZhPPEkBbEikQrKMDVfiV7Sy+DY+Th
nsZtZSkqnreV79h9kEUvpAFLuqu5MtIW4fZZtV89UnqYJtM1G3FKuP+YO+1UnN1Xj1p9nKeDNvoo
6A6XL4pAgrXe7GORhXH67ouxIfLPL6YiaDaFyN1N+APVDl0g/2KZUtqi7OmGcSvdiJohA327QA7n
P8cKpFAv0v0k2TNhbS8rxemj18OIWqE9Xb6q4Iak9I+VeXitqD6Y08iODfsx2rek5EvwGAfXn5/L
HiJEGz9vApXDxl1mjdOETmOD/wk8TdICGGbsBQKbxgZauE2fgkkRtgTgDrBLSjH30KO4CnaCgJrP
EPAl9YiW6kWFQ1z2G8SndHTOyRMR/P5z/s6+M1gp+6UvVb7pbdr42kYG+cqroz05wNV2rAKzW/dv
Hw5/2r1QWvoKkOgN1YM/c0W4k2X7LUMw1/ojfrjp9klDwlO4NSDYvNAw04BHk4f/x19tYennBrG7
KNZqdU1kWKNqqtsB1tpFB+K8nvh+GH6JyGxEjPx229iB0aTUZzOZsed+5C44Fyx68Vwzj6Qy3DjM
e3Ul7iztvaGv2NT47mYqTuRiTcMRXUyVkpS/8OdhvYm5GWYGv8c40R3TUdFbI12UrP8Llfez7qmi
1FAiWZzsVDIsixcArAlLhB+L8oYP904SqbDd0Tq8nP4nn01R1ktCZIEclPhguEaxNJDdOaum/CUc
1PjJAR+4mtOuTiL6faMbbrpIiU2tVlQ3UOR99qRJswlmvrBerBqIEu14hLNjglVi+N39Fi7ullWT
C0U/nRaSoeAlSQURAnOFRs9+MKwZtZ2j/HO1nXAyyaj4RqHCwZ/SG6yYd9amE6Zz+rHn+qM4gnBL
UtDXwQ1KxtBqG4lsjBDy8XFZc1WbHKilpN0NI+Zop4lnY/L3glD51ME/8Z19h9OYPuHoMHiVAAid
IWDtTu0i5Ksas4ZEQZKBBm46211ySQ37DFddrgW29nE+3KzfZgQJTKR+IHGTvObs+cIwFZ5rX5Di
zYUfMCWkYzdmZrFChXRO/GvaFf91DlY1pz4o7pNjKOrP6v4JUTwodbF2lGGR+GHsQeKX6sjuGD2b
pxQFQn6YZbul2jY/YheM3mn/vQJu/w9XFmffgl2uh44guXdeQcVD6dkCKlATuGkSJ6Cw/jHMziZf
JEPCjIWa6fdsU3GSa2nESHwUEuaM5hAvIaQfo7WGZnPbGmr+JgFaWH9cRvX+RlVmcxn6pjSvJs8d
AYDPM7lLot6cbRWxwB2ZbC9/tqg55frmNrtpyyzqZ/R7eceJ0W8y4cqZc68dQ96/XZOS0sBIPzA8
K9gFJvgEa0xUonXPjYI9JNExyjFTkz86Eh4priGxtbCxtAYurUqnA6uLqMqFI9DaxQrzs5x8osu+
FU2JY99ZJ5NuKOSPxLWzNQXdWblYrVIpxXwQPX+sZlFe8+dTq8o2Ecx3iCaE0AuOscKQSm3n6WDa
v0C6g6CyFWHvJoyGhQOKf0Xidw0Az52hiK7zkis/IsWVCH58D4uwi2ghoxhGbpANFnU7vCYSAVD7
h1+EKx2gLPyvMU2wv2C6ztImIqXOvYrRzTpBq20TRKwz4yxAB+DQqHn63CkVOCZTFE4DyluhQLYr
W2mnHuKEr+qkbx/5ombrGK4M7+ftRN8Ow9KvIN3MdzNqlw7RN0qJe5HsdY1YwvHFmtls6nU5AIc2
0FnHCLCPUxpM9dPaq0WswKhkaFh4BraWB+380s153HqJ36px/XXvP0ZGR7vt0f7RI1N9IYntKHIr
xBnwE8Rmw/kos8RUaNPvps1A0LQhdjaSnAl+/gieOjOKiWVV2YH4CfQL33d+ScojwvAtZMSE0Eyy
rjVXFVb8r217ic6yM9mfCdCC78AObBmTimCtSpmURR4QYr2Ehd4fOeXt+0TaP1qXxFhdUBt8vOVb
CxA0Ag6dhMXd5wdzBAVH9P0zyHgUveToaTInyRYbq4sw61AOLPa6Bly2c819hPKaV1tvyYNnJORz
odiqsN3S+9GwoyNXp4KzcJhG0m9Tknap0EOS54NupIPL2PZqkjhmfqvY5cU9zvivzxuznZLVdLmy
kaTEK7NyJ17LmDdOZZZ7siCbFyA/eHABqzXX70iHkOT2phfoXmzk6dvVWMOa89qDTcPUYNuDxjhe
iDagvh5yVxng5E23oTDNem+IGJCjSyEp71iWN4FL4vhfGyPuXoXPki/mNy7eapstVatW5TnaYH3L
lfsE1yvzEcjAPdYwp4GkcdXN/q+ihNV/of9g7pSUBu+2Rum0XU91HzyBGm1BFQuPSIaLfHCgtExu
4xPY8k4+Aj8AvcsKPeyBNm2GbzGu9rtJ+5fCSFgmBp1qTuETLbJPXOmkiugAmFzEPSrFiB6wm8Y3
/a7Dx8gLyEOKAVE36NyxAVnk3g2NSNkn8U3LFljnF6XWS+XqlFUD0F0KRp/Hg0rsvUppa+nE70Q2
nqtvh/jd0MUof3zWiRH4bxakxFtm4q+D38QoxxEYpfkm39S6OEjxHqUC7f/SKQ+ddfuIm+GM6fnw
C9X/DHEnry2R880ygKAS06TbkvS57CAf1LdJsZEB0hQmU0t/QzfTrotl3luo+lwZi9uA4Hm3c1av
QbNlpvdzhSKjfDpSfV+U9DOsgXwu53yDp2jP4XSeefq3Tkwbw5lCsd8qylAGkysxXsMvXb6arboB
V8jBVv3sZwkX4ULQTYaDgR/Q+sWpgddLc0qFdqQbp/BAenf2n1ne0iIofXWclF4ViJjtuLnc4wCu
GaZnw7pzqokwh8FTsN0q1o8LTKri5z/wfRBvPDrEe5+MslGzRpcfPIjDfK1svAMOoC+I+bshlt89
DW4ARuJiXjVbkkyukQArgzn91lQZYPj3Vxm+wMh6NK0eOnibdpAmH0AVu296LcsDmshRXa1IQIIa
2/4jCzHXx92BpauXn94oIB6ano09Yw/AJsOxR/o16VRUGysIUJp498H98zsLCO+VyZwNqmwpBnq1
1nFCM6WdmRLnPsuO0AdGQdDJYdxAd1X5kUSVR7DsllkPj7p1Jv+ttEQ9W0ApUfq40VtWFI+tXNq7
49VMy1CNIykgq8ZMLC2muKhsgYt9qQC1hHRwNIMuSfvE9nzSkFZeWK0RasiCouYa+Gl9icVgLuiK
vqu8pmHnCzGrLKfYW0IDWzNRlF+t9GqSPzEQoIXMerUYarAvtZMxLTOFVD3gSS0vw3xfkGG1PdaR
mR7M5qxuv2nOBY2ZlQiVBRTBsXHJ1zNzzOU8hMvV8CeTIeBo8C3Iz0yNYFJ8RzNaKp5akXCE58Oc
969IXtnA1IfhRw9/Nbo8loZQTcXMiqG2ka4Ck/FdlM3dTuzZDoNO5j2Xh9/XqQyGs/hKY6KAwi+4
6OT88xXi4+Z8/A1S5LlDgxsEXY2KvrfF7xn5chmoCWnNkRH3EGNBxvhl1VoCoyG9FK0LBeWp1zFe
xrMazUYdYs+8irOKHndiwEjukUF9Pj9TOj9T1aNWfOg5NBqC2qvWxtqnU8oo16pTz3qxx7eloIbV
21BzmpAnXCRjVeh/Hmlsz4INw5PCRLOlzy6TRWJoCHYSpMVW8VwUW3/7PoL8Rm3j32jSbwcGUndJ
bpqoCnkhjieI+PWVvh4TG0BrZSySS3xQqDYYD6PLGG5AMLrkvaYRNDQyMbiHmPX4RqSYEo5vbv0o
F1otEbYOZ1M9bNGzpfwexe4dgYKuFIsa2ASVfIHLKG3Y7b4iHxGKO50PXULQ+hcGi5eB1okRa/nM
3ZyU2v6NYimzjixXDJVE+dbdQSpbZenB/mHGJR00yOQtGlq/kQ/w5l8SSv0EhoDhUpsaRSLJjFFn
YWgWHuZCmzJWCzGzotRwfBeC3dAPZEIvdVOTHVnBhBkKlOTB0n2uZYwz7I0f+k9RWpQoNmzPq4cl
VENnc9g87xU4qJTtUiQvLvjdE6liFEjMBUe7bcrpJEhMi4inIEyFWYMgljKCLa+X0+5gRg0737pQ
oyowe48tOse+/pgEmxkbQWmRA9ea4ba+qVU9bm85f+VMHjnwsEJQkfAdLuUTJIcCthO2psfhA52f
dVtX/T8yfuw8ASl42qw8RvA6ZLnNollscEVO9Td3vE4tPSWIk7qbLl9viKmlZ7dZmMVDxT3BvQx0
Eeej2Lb7wGHSUOzef9N8jkQRG7ft1A+IPNYslQ+MECpoY2QC/2Ab9w1zBz4Tem8+hd8AmG4WFkAo
kiXmN6y2n6eU9nUf7ifFxV7H5GBnxbb8vn0DAp4AK4StPgulgPQGNiD8jC44BANIhk4vCZE8N5zJ
uL4jmKs5EQ1aqduA4LKXWm1jduwjiHWAI7KD/lRhb4MkGRX6CsH6yITIEVXb4xlVXQjF4Lpfmqeb
B1Ofs5qRqNLjugrf1nJ9yb2bENk8500n3BmCfrGRq500Obq5WoJ169xyjoODntDWagOo1fwDyYGo
anj3Bvt8RdS4I6/znZRdNhTBEgqMjsZH6YQaSsR70pDqxCNsIukwwx9LwFpmFhxSHlJaKuQbEB+w
ZMPhhdowOrShYUERmJRWW76ycp0WkPQAktYE9qGv1+clGheskh9nfTiWL18JaCYhb1ovPR2Ksb/v
R1dcSApmbRkTQoQaDZQryYsuAFRmctkSe8quX9e5PtRiKjKuUlcEykC5G82xU8eI6pIyNXbOxHIc
nfkWAjMBSjDq+LPYbEMhqZzolv88LhBpOpRlIqjOTwZtmYT82bovhNnd0uU5V8bLFpapN3oKf6zv
m2/bbiFBLAdkJeOAkS2pK9h/N7R6vvChlxo06QC8eDnPT5xcbSgFQ1olhLLswc6mGMY/8Bup4Sxh
DH8S7T2ZBDaUg+mhxPJvmqWSw/rN39taSWqjTOVY1UKl8uic1QQeylwIp19QbYXgkTIOCdNH7kll
4XBJg3E5+FjL5+oxCW5g8t/HfR3mE9UdDUoAy6ZFykibAR20dHUbQWXXauEu94ecsMQmB+Lj2k1V
REDiXpVP4fLWSIs+lJUKf2Y5rLQbowJKVm3wyJeD4LmokDRZnoCa3f+6saLVmBuKjSmQwDTXcSNu
X7Ax2qLp72HQrAUyiKcYT2DUO/V5wRukCl/Jv3d3DzhvYJHWGn6K3lMTj+szMmEdlwXqNqbVfxlc
Ul9o58hNU+N0XMv3UUJJzh86omI0H04LPkUCaZxhUix0ZS6062i4mrGs81EO7X8P7t79vMZV+aaA
sx4vewUnwnhXDWQRp6D8vmJWm/sUaGMoUdBihyw9DaEa8LB+/e7La+QtuMYvl1M48TyK5TiTvJmF
7YruLp4O7K8WVn5Hweb+Z+XK67EHtPSAuS0csyNF1UtjzTbXNtgyXHWytSTo9uOfHGON+adB7I6q
LDRchUtr0iYR7XcEdPuXQDQji6MMrwbsSLmduhAKHY54dJW+NLYERP2LO6V2xE7nY1PzF7XKAmlq
X+PIFzR4V8ijQgOD+KvPZ8XnysfRIXZfT6K8Hwc26Ic1B7S11EktHyTQGNDEs9RnVoqwt1iq31tN
lI3xWQm9ZUaHkKi+DjeYKl5R65prF5yN/QWjpHG5VrJ5U/mxp+Y43qPVWMn8iSCYzqLUnFO6n9Sc
8S+QxYR6G/VCz2hPNhNjpr1CJcy6fvM1SjObva4sl9G3Jn7CMbTvrElNdnEMw9zkut827fGxapMd
QUeYNeLQHZDEIkNgLVvSlzGU6LlTjAC1eE7UyOuq+D8DfrwG+3d3CvbRQAbqtZXiXjzqLpIjNhif
7K41wgo+rdse8ng/mRJ6MKOe+X1TpTzhb2sxtwpx8ZpB9U2y0dws+N2LjdmndtCvkx3GNWx1AwDi
i/zfTKxjIPslzEwOQJ+Tl9OCtn95L4gxPpdr27ocLunpv/nEB41sOADmVpF5jpFzohtUa0KcC5r8
FSHxyRaWhCbjxAqYniCdB1739sdAETbSDxeKEZZ/qKAYw0dFswLH3Q4jbATKGAK+5YIelugGQEK8
536RnWOpcCzKLS3J1TH+Zh1woaZh59K17+i7/gjy3iM2G46iDM8j7VSpgiXLpyG5V/93x3TLi6uw
wP48OlYOYE1y1XBLoWqpwPcyfUesiZBHpaEomMCzIHPZB82SFC3KGTJJruRdFpKxbMqvVWE1Scyd
8XZUZv4RdyME5Eq0avKi/3PVg40FZot4QSv2QgLGutkyLMsIIpIklsZOjLfIOeZB82N3cvxQyhCO
6++ZYPmZlC/BJU9WAnMFxMsectxtXoL2GyxMI7oqnq+sXU5paXvgGWZGu1NVNMrYKuzg1X4d088K
eOWWrJrTWqQdG7rAdGCQ4EhCqFM+8PY+0zvvnC8MwPwdgUZaKCBJoUjp/lUl7p0mFF6MxsRxxVvj
lNNcRV/X43oW4mhV8WE4D33DwSMtvnLMAXReuJ45w8kP0IT3ubp8xOTfjq/hcHz8Yngo7UQ0/Z1m
5qhgeL1Krsg4LX/gWjAXVGz499lo9t3uTEQ8B8crxZFIJPSAAV1ei/zon4J3jkshq3jZOGDRGPBw
Azkvjq7XsGhsMdB00qD8bhhrsLciJXDK61w0dUAGQpg36gn4Pw2pIk9OpKLkRdtVYwvi44Pw46T3
kzAoCYoKijA0oEYga66R8Y9YJ0l2p7uU4EYBJaC3LacGQHPHcpSI4XFkwk5Rz/h6N6Y+vxyOFeEm
mBFFGuWBf2SR6Ffe7wIoF80T3cRKgiAVtpvBtLIH1vHmYFoANv9b3dq2RFe+ynrzdNliTzk51O2O
8/4ojR2+4ZpRubD9U3Vonb+g9QdA0YB4TpMUfPMZfrxNKmbs1GJbio77omyoegj5aYzveOO0NoPR
3zxxE8KRTfI9xhFC5CxfS99xVcA7QUmIVYsbOHpVDpx8nsXvYM/md/gbv3dGFSYoUlYyelqP6++X
dQ6ee9pTDuqaNa/SB23GZELCdhCRUPfRV+w+Rpc1rtn0peA51Cnz0yjLCLixL5gACU2K/0XpXaEi
K8cT5gDXghijGtFwcv+S8OtGrw/Ul8zhjwa2fj2rv+Lao6kbEPp9R4f+q9ViADiwWw09wFqkakbV
B2xPwwSEEZ8GGJTCE/Umm1z9YiOUp+IO1wz6dEFt2lY0BaXxEdH2AbtWzHPyjtzepzEvj3O5247Z
fD5+HreMQ9wDO6akKG+A0BX11u13b80rm6cxiCTTIfszNnlp1F0gEgSDsZcPYG65VQ7XPZCCDRQh
IZ4Z5sGVIvrTFPWhJYS/AUBsNWllgpBR8WzwBIfhTC6q771ObVeL+CKiQ0O6Dc/LFIKEgKVKWtmW
Nd9GQX6sT2qVGhxC+WYagyKVN6D8zqQqzl/ikxSZM8VvI8OspK8j+0LOFBMIl36Vdy6wVLhL1e/V
qX84tCCi4w297QiW+QmnkSduWMEzOli3/kY6ihgHEERG7h/sLYUGhQ1IXshAE0jnWIaxdB/MlwXn
6FeRBmnYUQzotNzoASLqLBCOxVZESKEmPg7JpQv4DvSCffthHJlVFS4UGVeznW5OQ5ypWiKeB1P9
1Mi+x1OPpR3ZObXwSBf66iqe4ODV1paT+kckl6XSY6Flxp8B4i/cnrg1licPYvgjcwKl2I80hBAL
pRjeLqH8P99B6Dr4FDd/onD5GXjZnycfYSMhd+tlEqeeG/Onym/ZWE/rWWISf3ARi0dIUdhPA34t
OmQYWetEZsHeU+c9cFa8VGmw9V7eHl+4k1eM/8Yx0mnXQJNnHBL7dcECsBoNkAO8zq0JFtC0EC3v
KKW3gGm09gGCal+Ar9t2OOsLStBSBT62OkfWfW8HHRAVKc+JDukJI3tUuoN6p9fpuroBqeyz+1jn
JGXPbDDQbnFDw4pMCNb12732lDNbtcd/xBsJjcrtmpxwX7nxqI7Ct3m1vJFh+5Da3wZ4oB+t2kOJ
1tm24ThNNLnCOCg9cU3zCxHxhRBdOMhmdcxAZVS5hMgXoprQM7hv3Yusv/Nv8L354ahM23Mptz7i
deD/YoJzTlfP0MYvvBQccfEPbdHttORjwcg6C2zzA5yPFjaX/utPZjDjiB0O6uCCy2Rt8rnX0VbL
8qUl21wf9W/NRRG309ayT/5qIol1eegePtsCcxe7jBVa/XDEC+0vDT6JAz6ebAH9wixxlgW79wz5
hjZZ0XUAailYDcAcFEjNAE78Ea8iSbwgJBjrgsaYgnamLltObuQs+njDSEmEL9L5NhhwloDRG+F/
0rC6EKDgHk0WI+SfmNpeYDfAA2mPnZ2RfWIt2w1iGjl5LGct/yRkgSwC3+UE4pi0pfe+Tp6EdMml
uB+GBLrSvjC3guGjCugX8u+m0iFjY/dfQLE2xVMwXjnbgwfAz6Gpsg6+ebJcyrT7PjxN8krlny86
WRpua0zhQSz0x9HY5pk4haub6naeryDR7AMVdJuPTnXp+AQPklaR7+qVHoP0jbfg4rl4u2sGZ1a9
qYj+Wxz5E4wRVxr3s4RJeRAUW8aUsuDW4HeA29MKyiiBHHTKu85/Vh/89P9dyI3C5RbR/CGDH5Vq
bqRG1WM6UW0oY72Wdpbs6r33AjcdV3LgYlh8lBWhNWTbffUFvRGiUU6S0DYZvGqqkIUwt/4o+ZHn
3RN1AjjuXR8HT4nbe1iKy+z6sDdK/muidqorDVT9WOCd297kR97ihUqMV9T4TSsqhwpVUKbvbwrT
zyA9uKtmG1ICJOyjn7xvN3qAeBk/+/dNt0hcqJs45De0kFgVU9skdOgxKiqCVIELJw4829hl92FI
sU0D/sdTrjP7zIWGL/x5vVV9wU+uW33jM6alWj21DT5TBFURnK6E16Grq9yf4POFwEABvC23CMJn
f41+zQd1zo9u2+AJfSlGZziEjr2MbkH8AhMwWsEMjesuW1GMJUY0doCZSVr7YT1+HfdwP1pGjX6A
pLJmy65ZPZFJP57mcDxKvAESuBzedMHSsKfymhF/TUMziGhGOU9NemOMoymcD0c3uWwWFV7/zxiz
9h7nmIMCS9Lu/phwOC2UuKqD6wgyDJw23cJ0VKutd3D2VpbNLfWX2tYOImlX1b7SMQ7rpd8NLxex
93RX7auu6ejNrgQS10za/w1P2Ab5jlfgBWI+rIMkgq4/VKwKmpBN6gg9jHqiqKO4mymRxngZ1Z+z
ddIbFN1n70qg75WUZ4DWFG7j806BIsywOFjVseXleN84xYqD/eG+gPWdkeYP1akxsO7W1wbyqjgc
FlDXVYrRl0IRoARF0IlLgFk8Z5xHr5S8/zEwvzhSKoiowpZM0/LsKPqAUoRF+8T5+vqT3nre7gOC
tCLuvb1QiVReahuv/+EdTAHRQoQYhbCveNT81IFtNFnWl+GC7iislEU6pQtHZ0yKcMjF1//p0mc5
/kYkKtYGYGqMZONdskWlLPfYDwVruGGb+f1hJM54wFxbWLe9CRoemLEnyCiXtW62nh932XYyqXLQ
7IXI0lQSF+zfKl7lniAYhFj/ToqZ+fkMJhwpdyGXHuCJDltqYnffBTWhSgS8GVcULkOLhHNvrGwG
Ok/it7idSbENXDgCNYn+2qOuoBUIXqJEww8klgSJ4LGNGJgstiZ1n5PUyxE9S0wJiz3K4ATfi61T
6vlAg3QWWQCJ0L1q3cc7O46OLXj+9Hqy7T+AIlpastWE69rzq9hTNBd4pFp0boSr1qbq4HGEfUho
0Pc9HkBeeQyJbbY2leDeeSaN0HGhv4zzpd7ppJ5xK7NOiKF5YTHMCzd1VTn8kScidWxGOOB3Q1Of
ilYzM6W3TXCwy9S4yQYvYAmGnxDv1VoM1XhOp66sYa3k7tkGdrFytKaj1lFYpt4k6nKLtfDo1XSH
P+qJ3U7Oi09iXCzQl2aRaXFTgAgtaOcMAU7+a33w6PBgzPFCGgMFaxTQj0KVvopV9wzp2Ue6yCZ/
IS/4jQIO6Fg8yO6G4zS8ZHIJKd6Rh4kssUad5okV+ecaZcKHLdTZnca1ICnYQdX1iNr7NTjQEYJ1
FvmtGWFszXdklwc1XZ8DTBz2AMXaDsyEETxRLEkae1mgVmsl94B0nKp8zQUaRe5PE9WsGNCDZ6Zk
4m4MRz6e75B5J+9NViCarMweneCV0YpMIkFaGjBEomdn/OMSRZ7Bjf/zkkIrwlV7eK1qTcwk+NVQ
QDtPcPYsedF+bJi4hZxQgv7TtYdXn/orpqLJCeYZA+OJ6peTmhGOY6Pb9aOQgvwLpwRcUnZZ9oHq
f7INUSc3/xRhfXpJCVRMCtFPPgI/n7J69Dk6PCbBFPkpK9TysYfUyWSbF6mvbLpl/vv5JFFK2DyS
Bsgrf9cBTBnKin5EfgS3Fhw5WUInvI+Hbq5zfVK7ZYOWys0es60R6tmjms9HA5EDXeZjKJrC9mBJ
Aj/Wl/PTSzLUQxv9YMIz805rx1+zvQXMftkVRSwYNzzWr0CD34u53kpi91fRy/EMJF9VB1tiaOfl
9UOYDu7ALdc4lY6r72DJmQl62Mv2UW3FLlLWRqdL/1Ffc9gaFHVNl6olaFZkEC4Hq9UMEx3lfNrw
tf+zhlJV0DFaKKYfO5AnYOm8EpfOKqM0nvcqlzjhNY6wNScFdP8ekP4akIj0Kg6+49RghtZAccWN
7GUUw/SbIRC1xxMqELzQimLubsuqPKh8ncJrn38N1olS8SE5QN4zcK4EIab+Zvh4szfjvbJOHp1y
76c3Q0EXwYTogAKIiHskaCB/fMVLtCUkL0DzkPAxhmxb1XCet1FYYzAjU81j2rwRHqD/H4AGZb1J
U9lPAl2+Nn9NJ/kYcmzR1V6eQd4mYV7x4PJmdB0ukE11cYHvwi1H7a6jbuTPO5ILZlZ4aSovjzE/
dw4fZXOoe1gZciYSAXmSjp2Y2EfCBIXxXeYtrDXSEzNTitX2lCcAC0AogqRC56PSdfh2rLPVFuJo
eVskugq6XQv862s/mXrIIYsdLwu0tidCeK5buf3byU7ism4/mI32ctRyUy9r+YBPofFbcZGiDEuy
trv2D7bx8lVt1o9Z2Vio/zLDaCSW62q/sqEmQb0LVIQb3mBKayHpiyM5RUiLSmdNobLYPy/Jn2W3
8PDNBcVA5j8Qo/2Y2l6O1U8xshPeY/97YvUPQ247oWZUONL+jdVouksLfT+DTeM6u0bgPVxsgcaL
F8v1k6uUjRgUiN4p1KcFhUDGEy8J849BYx2JW5k/S1lCC2hwD2ZcXjlocsc7CP51yN1KlR4uv6V7
dJMsFnnNVX5g6VEBiONeDfKOoaDqkcLqT435WSUDPy1xJnpein2C7HyZf5hXSOm6mfQNEZJnMpuF
7z/PEssF3yr31XpAF+EFbsl5mkQF5qsKBzaAK+oLVvXVvxEfid7CuwM96Z6TPro3beNlTHIXdf5n
qT8TaNkBeIYzJaWMv/c5H5Gcj/EsNorv6s9uSiKf1B/htRnOVz6yoFYPOpQaprWvkOHVZ8lkwCN9
bdEZk6B9YnZ6FKXKyrf9FvGLRW8w4yhCu15fLQZMeyxIhuNbclSb7XFh79fDjrExMsHOsze+5xsz
OMWoDpZjkfryXpLjIu0ifEAvrZRsR/Awuk5ZfLzNNXIxU/KegBlomGEjrdlyl3SPjhh/7wk2YS8l
fyxn+37eihKec7Qd4HLWaFYlF3asP6KbiEPxUcVYZ94MSWhdgPT+QqFeNOJ9pqqjlpxNUzxjXu+c
NwhkeyiO0cFxknvQY6cED9cj4aU3sq9NhiuAeSzbHfyYAH7CgTT84XXumuVo+BwcMuM6mgVQ01LR
cLCIBjX59YVeIUO3ovL5RtU99C5J69cC4/dOe1f0YHVFQKibwOshZuh26eo7H2KTKC4GbOl0X1dk
du6By5B+EQMpH07N7NcMmaDbBbP6NrtYsRPMAlzIk5Hqk4gmLFtfCaFQWqgCmtv2g7zSUnDJsjVS
LDdJGbz3fFTBUmIXcj1yN3wz8Gt4koCpM39awUshHzEyHPh08/11wWGReQ9FK+XfmYcPdJOwEieU
JNaiAy6AEOt+XYhAWVTtjmU9vfB9dqeX8HMrFOvNMJUtinBwRFtk+6TpEEjzCtTpUii4uiH7LEI3
jeojYiKKLD4gsSY1BiC5jZ7wzNn9gmsoVs9ZrsBM5u3sqcEVo+aflyRA8tK7u1YTh8asntZxa6QI
oDzTHDnUe7WqFZ0szRIXxGfjRgUSygESZ7nHQK+7sVfH+gxfrDvV1j7L1Kk9coZ5qUXQfNI2Gv8W
4d6TfGAPueWB7FEpJxiuBB+BtqXwtIO08IJ3yLI4o4RZU4pEKjfy84JrAcYKx+qHoGSUSnbCA/Kp
24AVRTU71aAftOHCLyPMqLmIUsWxF7hg+nFbTD+Jyo60O8NGvpcm8Dl2orlV4Ikyrb6Ws35aFEgf
1MPgccjJ1Zdq0p4khclfq+pu0SSQFjx0bEL7nommH1eQUN4cqDXEN98ERs436/JJJYDkUA2/Fddz
x95O+BYL/ygU90eK8BZ3YI+FGF+oI4bjsMy46X6MX+BSnrtD5wX/75wztWZ0bNWoeaQnw5zlZrWY
TXTgdLqnTEAZGdLfKncu257dBSbL+UWwPEQAZOk/GqLQwwNb3mrs7841YzMIeUVQ6oGBEylYliUy
O2Er9nbiuLnosvM2BLS0qbYyhufYKN0jH+yrY4/hbsTzCK0+fWV7SeyQ5mFaS3ut2DMylJpL2MDs
N7ZZfBpBZPqka0Z102efuVWDADS3oQ3f9wxjbDjdDgV7NrYl2yv47FYAza/8kIPNUJVAzP4DGZIB
Z5qmTGQbQ7RFEVx5/Xl9+7YL9A1Ltyr0hPJ/HSC/tr8/Fp53qocd+XIBIqbGWJ1u68zZ8glvBoma
gL3lYh3SIwVB/48hPalBwVQa3CgLljobOOeKkuEfecOyNrFv+HXNgU97ddG4skbJXlSKYncUwEe0
ddO0MMjYytaiKXABpKH2Dh5vGy1P4JDDC9UrUKsHvqWdfmBQHNsXxwWZVsuPNmbIyOUOnLEiqitC
DgWh94kAHs62bCpa1UCDB3E5Wu8jmWOBcc4bV0PVbaRLI+rpwQgPWixrJw7B0pb5vcaZIclGoDVI
tWS96Px9G54kyWZIKUBXt6QtBHBU3q9k+ZFekzcAUKjakyBuel8OtSGWt/UYVzszWKUPpJ38AUar
rXLJx4clZXLPSOYvplHsIR/WmNJ54Dk54dGZH69O3yzIdS28b0s7hOftqG8IjwvwE6HNXzZh34iR
qqW1h8ZlRhUdIdFfptRJp9zDIeSkaFUMkTYB267r5krNjmnga8471F4lTUBXCObSWEgtcsfNIPPW
IDgujWrwKDt9z/LZHKz8kkxIIbjo3Ivj2fKh47djuhOsxPUJHaYZnBod9UTiMjStg31DlxEuCKPX
TuMewNuQJH9YTA/tqtSSF4TJHIaBGWSHyf9p+Q5upfsvAe+7JeO8ei2oHAdJcCcaDumAQTIUnKyh
JnIEVWG4HiDlHpUyUrZ2Q9DxZIEqUQQC6oD387afAEe6g0+mQ7LlpOfmjUFTqk+/AScPXvT3WRpU
ON66Ga8b3BB2+/c9mkHB5ZhNAVba4saqOzv6ik0CFywLx6xq3FEmH+8aGNMuX8dJN5+j5b4L4K9O
Qsw1bfqj9Zzc5h4TudmhAggat3x+1LxRapRe+VWxnA/ZS3MmgkbnQrVJ+zX1Yq/8PV1VzRmxk9pe
ywo37pqwjETharja238RG1KIhiBpDgZjMU0lkuJhNgUtZJUmuen27awN6Uo2vf6UyvYOHfSQUYCR
xxv808XpbNhxy/5QC66574iLvdorDQaRz9ifx9Ne14bbHL8XmAU0pF0VoOVkGitLkAMgdONfnIUs
3G2LV+JtoPH+cZrWhWjD51Rmsj2aXb6/hh7PQ41Kj3zcjhsV+RvgGOl1dEeWSsh39bK+A4wewyDm
XrI0HucwzVF78rbw8pnFhdKlxHsZBjRKkD9PeuFOAI/BC3BqFBXEmF5YaG9Ddoh4PNN42kZzMEhG
RciJjVEhRulI/yopGdE5gJe6PiGE+9XwaJjW3GBJSLvmS/mkXEcsXAlNBRnqQeDXM1df8vK4U95d
gmlckvjE7pRJWyLAYqGcomQ1x8A7tZh1fJIzGvGRWQQVwdUEWN4vQvL5vak7jagah5dmZ0JUDuOo
UJQFgO7qrbVftpF+PR4Zpjl8W21390wJgz4AU5aKpFgfzQa4qCzT9+O2vWt/Etqtqx9mi6wKJE8L
Ew2YGRlJT4LUVzYvxcff5OSeuKMD6LRwgRAD56Bmxg5XhXSyah2pquUcFLQKagRRNSvxZIjJjVME
MUxxgYnDMtxGijHSZgEG13ufH4LqkopXj8sGCml8EfjjLnViWfS+7Yxibmw6x2XqjAb6mLiwACUt
FnBVvbYataDTzOQ1J8hqWKVT7NDKhagSVuAQQcm2Oa0q7gSniMDU5PQJV9j+e0etGGvKrcTH6GNU
oce7KOThRQ8y1MPfnEmrkCy3ukAzQoBlixjz5TjO7nfpq20p+E5zwp0Kd4Bh5CdZOVnwWlAVIYsR
CEwKwHbsSbi8cXT31OHDqC6+oD/jS+fhgIGsNMS5hFwj9TrsPSMHQHPn2shJifhKlRrbBOT+MtQ7
OEf27siNSEzrfexz8cg00RZXKSmXmNriDa5d78R0VCJhHa8Mt/VGK7jbSOsGsKellxF2pj6jLdHR
QtrTVYHYZPNgGtmHfEsm1u5nYeZzD5omnUhJXwj7wMT0U/Wpcr0L1suGRI8GxMx2Gy6Bc6EjCUAl
p9VpUchWfEbPRynNRnGoPeEeW68iQNVKah1jnoLGGVTMk15V7Uz7GDSCfw7oEfBaHmSjEy80fGlL
ujSSwa6QuJYpRRgWDEJ+diqYQ13J9SQ3AyR+UwMr95Mc3SZaQie+j7OhxV2qJyEPSdqe8BO5MvBe
9Af2xluckXLJ61QjCpnpS8setBHbtrAJWifwx7oFA2UEz7890F3G7w2yU2pUqj4eSfZWBjEm5Lpw
YwGXEcTcsiMe8n03PQkprpEqkRm5vjWXhREc56W80aPqFq95hOqsJwZQQJEzoL76dCmfXlJ4ASQO
nFzYsM9OzW5O62pM0MszFCWYw9endnrNfkK4jOxckotFu6LWUmoiTjfy6HYQ2s+aig41OCQqJMvS
Ftq74lub/2fn65LJetUn8TkRjnAUdw3u54ja0xVMC//JXgSEdUu+QN+faK8tUR4+xUzx/mCu1DrI
tKpC8v8GrsriNmshk4MWhsVv4G/ht33YMOaoaNVI6Gl1dVS0R/85F+3i3BmW2rxiFwUr6kZGbnDU
9h3SyoI1C1oGEkzI+Lf+8JvAxWY+cjHJI3tuYIqGPyGgLbdmqjTv0N+n4cbEYxWTspCekXkFpp93
ickgSL9f/03xwEMEIixF0HcYrMik5XzN89k+o/ivzJ7g8SfENC5fAErv4O/2inosdVOgaBKKEG2c
ErnIoUG4Oly3z0ySimDa+oC8rJzrn81+B9ZMS/LouNp8Rq3KR8qZCLyHUAvMQQFRb3I/JPAIMEX1
RllH9SNk6yP9hppHVJ9cwaLejpRkq3kRiTEGjbUAR7f2359NfBQk0mMv5YonC7SGby2K3Q4VdYCE
RpxrnCKuRGQsqrpOH49l60rsSvfOudle+CWmIHwrNLCfLXRaOiCcGcanfiJQRcjg+QOf1oRDTUW7
seaFWNJD++1VYtQbT9S8z4zD6yOOEMId0bMMByHYGbWWUOPeps1evRrlUXX3nQ09DVqIR0DkRlQN
7FqCZiAKWl/A2Md0qcNUryc0cmxTFPWU5a9+9UYGcGRfDAz+QIe/Wysv5WRuUYM66Mdrgcj6+U4b
tKgVOEFXkaB3PWNFklXzEbvfiSOlkf3FymYmsVugcw4N7ZVJRQF62sU++aQ3uF+MmG6Vu3yNyhLn
03bYFWQo7dtnXQWdEk5nbEp88u2pAQs6oGCem3p67y2ctMXxC5DiRZGc6Q29OMSUF5NEOBBDAed7
bl5VTfUZ8XATnkZJol9ejLn3VAYk6LjFw+XQ+V+wPjhWEuRz1KZkApgAnTEIkqcyR/xFAeslqgMC
tJACto6BBHSlHTtdgtd36ih9Pu6GAa2li6XIrhK3u4YZ08LaU5uLzloFY4ZPxl3kPIF+GmSYExFC
/48sJLqcl0hLrG1Q1PfvbV00t9be0rRWeo7SIXzyxBnmdUrGZDdFR4LHHYeReezUqC+KnRycCE/l
ZLpM797WHFYq6dvK5THrnD2Ifu1HHRjzQzlSPZ67u6UCA5RMrb6O5gtzRxlg2iIsEsyslVR0yuBv
H3R4IRbsPNUGTXPp3S8mVF0UnNXGHWK4Y4UzYversBZoW6Wtd7BsSR35Z2/kud1ca/7Cm+nwGMLy
B6Q48SecAvkNfS93rJ7cGTMvVYhc7jfqEwSAPneNRGaXaI0HR3s2Wa+6qAQotdAYD6nypEjRY5gp
J47NWNWDuVpY1gX4xvlAurW35TzQsbpi+fRrjW1/ApdR1aTMs+1GQ+3vOwdU1hrd+I1MYhCvLbcJ
+fwl5S9JkFPyWk2q0EqpdeDbEB6tnVI+0DeOGrgUkVmO8j9LA8DWTG7U5oj7/O1TUG2ahE6pUnT2
4dIcOap9wzezmgIYkeiMSFiCnlT7KerLi3g4dY0Z8HVIcQ8YGM4vw5HOlihIeCKXQs1JnMgF0Rch
+Fkl7kOYrNyWDY984xh0nnugn+1FvLnBp5FF0bi3D/69Wl5qsaXO2hhNuCN2GnrAz69MyqRpNmj3
y0A7Z8x4WqTzYW7eaG97I7t50lw4amL/gXBmniuswLsm8Qwpeahw1j7ZsG2APpFIGrMF7yRMLuHE
/hK7sWQMKdGd8au3d3PKTD5KcvWn8YsY2uJQmQmLJ1J8hn9uHhC+Ayxd/uLUf6CnWevlC7LrCyy4
fx1SUNneZiYlclDiVAw9RkbJpKv5x7SlrPEXKdYPro2bQfy2O/sOwIqu8nfkhq13ceOLfzxqC9v5
OUVNos/oMwezVcOyCowWRz5dg4sMxAB0P5S/wcGe8LAa8DXITkLtxdd82Sb554tvbTJ9wK9X/GY4
FpyQ10OBWERvz+tkxiO1gIyqsOFOPoNib7UDA9ljWPt1URnGaGHcKyV01N8lYhgA/if2/TgCRXs3
jKHrj86Cu53rCycdt8OS7lZJoQZwFbVwvYGibg7HLbijDUuVy12tkZeoB1HObGYW04E4h2PkrHhF
TCGTPtmAQhTbAp97otA2wRIcw+6qGxONemoLRBFLaZcFHDyDWg6DwhVJwc+Z0EyyOiHcKyAUCMYg
7nPgRiA6ayRGhKWOGhzd9ZJVpyQROMXZYjZ7C39YTNewRNFZB/0tQpOICOFNXSNAwpJe+UlA80i5
cdRqnvhGV64E+o1f4Wl1dg4dotMELsOg1hXJ5xsSm2cPxIlwPt2314xJlZoVedYlWaqbpWxWUN2a
k4oXTALnyxCwlPGd7IaAujw0GrlUnuJ9ArP0uAIQlMIME2DZNT8aA821yRWJMbss3PvAV+LbEGjk
ULWy/S4SoqEP65MApFEthQ2Jc8l97LMMtOqx+y7gw2mos8IT2oiFwJ/Ao6WbWuxBDRm/xe3+S6N6
jB4SMfi3cXr014xPQWI1EyjwmCbfJwxir+2TLkaTm2RhF48r95jfPrDU3X2pxqTMNDuZms7Mdj5P
qpGiaHU0NyFxGNfRqeMcyRNhTeqsGsS+htBCHhrIr45VgO1q+umulmrG8a52qfvS8ODmJutrcOaW
e8gMQlzZepYCRv1N3iBJRnTmTOCdbckoO8/+1n47K4/2sAksbvBnlZrG4UaVCS4Vua5CH1a/uDmq
uDSPtOgQHsz9BHvSDH4iqCex3u2niDLck8b/G64vGWuQVV7unxdP/sJEuqyCbQBt3U6YQcQZk8on
xiw69M301Z3nF6+wnHQX3UebKr1V+71VKQ26MvCSFJ5TcbGVUzzjmJwofXmf/p1VpMiWA4caNLVN
9AXsW23e39GoyJHis/h/gICECBx33gXJpzLvDtM1goyYFRNQUdN/NnG2C6GRzxiUGIA5vQGcUtvR
LyXZejKIB4tR8Rcm4sc9SefxvQp1JnwsfVI9u87jBx/1rckg0ifb43MDoTeOFFy6lklsTiEt3s53
Mup7DPh6cgmW0t3xWpSWly3u5XujhDovUXgiX0y1+xcRWVxljKm/vQmDa9XMT17l6whfWwihdKlX
xk+gEoXlXdlt5tdgn5xQIlxDYOKtG8shujgz1znuuyuMcd4zY6R27GqIe+7wtC6g1EqcpYiOPuB+
SG57RVI/beFjlVXLvWeSClJOcenyR9qdfdtl0dUSamsUGzOIGJ0lyjkjFGTkRhY4MhGUu2nx4YS9
2AVODTzcym3vhhlt4pQmj2+udzLa8G5Vco95aLtwAO9Ik1wKPmbNxp2Vf7QI4fqjbne6C6VaXwbm
J1Nmf0YG3eFmJJx4Q5r2PMhDBZ8kGmtaru2oZyNCe2eybaiQt4AsAUsPskWmC6fMxiPVB+ltXRkW
2qpnfjwZA4kpkUdeGMY3xgtCrcvIs12VMvaH8AdAKsa7Q2Y1I1jM+FPxeeMEgqgbZ4UnJrRKUEmp
uoQn/YIfwuU/BZcmdw3Su+31nJsi0VaJTcXFH7QNHEW4Ph+CF7c5p8+t+ITadI1zj3U9pJJtnWOD
AtqItd3hwBpZkvUqE1d87Ny/k/Njyzj15TRZ5q1vdedF3kACKcjeO2KI/Wv5AZenuL+b8CBm6i01
J+m5Na6U6yUi25YN/CfJWpkWiJTvvkAbhLrUT2XGoI5z1Wk/3Ps8S3iE7X83qnhQUiLyDir4CUr0
Gxpr+YVfGm01hMpkUUwrvE3sYUTDjjTY3LJhvAvIKSR15vXaY7fcvuHBDka9W/96/mOi6SoFAT9R
AKQ2xRPSsGYyUCUyMMgCuweqfscsSzo9ziLTK3FM+quRgrk22vStAVJHkc5eLxm1GFkjjupcsBgG
aDu512UYgeZMZvXRM4nTjL7CfiH1stkT7PqgdBkrOXyUGbWavvQ7AYk3/fsLjC5GIPz3rRO3XrUW
E0Onu8K1xOwmvWsmfBVTXp7ve+WWSl8RBk+kvlo3QfFBaI61/RfKq45o/RIha1bdnrJbT0gtHwQ/
1jBkk4Q4L/lfoPaiGlkE4UB5iWtZ1yZ/D3yS8BJxClzQ+5JpR58q56WT4ni42KcTLluuXXOXFmuK
Ki3TztgFH7XOiPFaDcdCyy+PDKlXXHeviaHN280j510r+X7Egp2uGiUN/CdNRoSH34nFVLqiBHOy
/mFzrkJxCJ9ZXP4/b/nPjEpRqqy61K8AjSKAkORMSwWydM5fW+aD0iWnV88wlrXlVTzNNoli5zv0
XpcONPuQViXYbsf2IaODekl7sSdvX3nsyXHik7hQulDOcNqSrpqtQl+CGVjnxstOeyo8JuH0q5EM
cjdEmFCFdq9HD0hTMoj+xHjdiKL8u1dzVyz/hci3jwm8V5NIA9XoS0fQvlD9hA3s6w1mFjJ2e+C2
qa3Ic5qBkKRX7HESOcnUkDAxVihG6LOxSYbw5wIJgOg8HEEh8Gb4AgdeHU1kEqj7cW0WHXLgchtU
JQTTNb9WbhPvK2Ed+wlSqv/gX/IGum6PODf3fF9erf9broYK5y7xGXNQH9co5lXAbf/2lPR2CMDe
e2p2wFJjWn5GuOmkI1hRA4WaSh5aPNXxc+DG8rroQoDl9P4uanPpMqDKIHgfsMPHqjhNXNC5SIx1
MTncNqv9fIntoxL09hk0/TofvXs0NgjSLypHJdPqo6zJ8xMva/bSseZtTrk7CJj+LbAIn17uNkcO
jc8GFUNh8o1pX2XMusTYlfiSJPI99GiVnWGpVMb7Ofwp/X25SppeFCyu7Vm6kIlmDFOkjJxa20h3
rSW4Y39XDbAKiXGTO3I+SaTS5sDAgGgvr0zEuEMnWhq0YDMcA3z0XKWVod82lkgVBPiYeVn05ZMJ
7oWf/6pPAx4akLSFSM3FrOubObfPaoBZgG6YKGVmPufLTZ4nZzXbcwGjX5L/ttlEn+YDIAdzCj4S
vI18bfY6ZI7MBNrLI+0oh0ClneDyiOPd43KeCj/ykwJ2etfuPr+YBo9blrZyO0shRCiHv1D8S5Ds
b0l+GFSRs9b3Hbb1KNniVB/Q+sFz61jCr/+nTo6uWuhlqgYZhbRzif5Zz/PhfhG7G56n21NJhoBf
pKz1xNRldmJ8/EBu8SNbOxfddoi0I5vE4XpPZFG8DGdY570uLLLFV/oW5pg/umQssCl13bafUQgx
p/iUL4rocHEyTbF740EHsScMxyRcz+JBMRO/3EO1zSqlajj7c7BmqC6e+HjrNX7deEOmXqSBIGFE
BaKG2bp2SKEcJq8KVO+m4Ed5ujMdffpZz2E1e5/qO6LIaOK93YFE2yGVgnNsHZfPQjyISPg/oEuu
MT0jVZpUvRehnTr40eM3pmiCRSc6QS9mbItJBOzYtRZxOV8kBlTUkAjRpLO1s5+pl5no+429TInx
OoDVZBOIrTuobNOURDy6uMz+3gI7AezKSEIO9JBa2znLc4E4106iQyLCBIt0yq7lxUXfkQn1D7h+
nvLlFxCBU87VzlbePxMzFdgOZPFbgsLorQCshceJD3R4Pb4uT6vTbJpjGl9Q8hZTBrBnd6tBIaUC
BfFwC0ujdvWPx1zKHE1WviqUOzkB4jEvnm2NkVdonT1j5YweP6Ka4yOj4HgpsD5kWM6DvSuj9X3z
ln3htZ0xh1yFAMfpME3JBlB1LIUXp4UJU7U+QYzOCYIZlI0QbpZpkihG7wN8VWTSfSQ6Sd6pbbzz
AN3v87He7SWl52zSv6n1VgmNwQosK4kn9Oy5DAbDDBXvbbXfFx1twBSv7mCjHz7RLWqfhyuhrLHN
zMFLLm7gDnSdCcdWNoDp+UOZRgfA0L9IiNawfFU2vQUAnm6AT9D8ZWJM9Nm3H7CXVFh/rmrG7rCp
k4kIHdQCbJb8feEvWESqBn+SMo8VZwKIVlFyN5wkM7FV/8a6YXqY3Uxe8P5r32z9qIuhpULF+E7c
CbM26pk4fE0K6/kZzm1snA+0QMZgYDeN7GqqhHGYwftOHvcpOqFA8RUSGsSSCr8LEKj5KXV1Sfcl
KBwnWkHN6X71XqbGjP8zOfor6DlsTQ7lE+/1lKq9zj8B3wkpa5ul2oD9wQJhCUrXJ+sBlYytHCFt
LHCLQQI8uoAYLnqBoGzZqEGL2LjHFVuivDRqxEId2VPXpEPJuM+rxQbObLdRX99WSUED9aZLp4dD
+lKaoNslCtiAS/5jx34QW+AcXlpv47sHTAVZT6JCmOWx2ISbXdN/HTKgGnz1t0ofjmLDZPKtgAXT
gsWJ5/hJDe1oQTtbg2x9qpF9+z7m4s3uSiGv+Wi/S2iu/xwA49dOBaU5Uu5YAY30NTml9HX0bZOo
ZrEfA4alPXd9XHwdaHKWy1aEwj/e/XeXSYHLBVMJCJwCwigyWCtyh/+iZEsk82usbtSpx3+UgVKx
tJXqzVGRBGyjFSYJMBw510eQZkjNEVDCfKEcn6xoXzQkmYwzBj8xUbnuElk9Uj5U/ZImOLo2/nou
UMdtSKXVpPepg0fsgKBcZ/VMExEHFZ3GA7UAZUYHd5i3QLN0SPU/GyauSqvWqaUkbkhtG7xWLv5e
JKvRKb74WxRZyPraDOlNFURnsJEPRvIE8LXz2OwoF401b5wXdq20jRwFBMa+LLFO5CM1E0rmHxQN
yx5Lwdr33aHjydy5ubT1OAhgPi8Vf8wBq2nZ9zDh3jogphSUWan7YYiUQysEM2TiR8P+ChGpdjTi
ApRkWJ/8qNbXNP4M8a+hzF+gGaYV/w1j9n5cq8bboc1TCnq3oyJvD2v+gNvWMLYa1YTPjtLT9dWq
VMmeuDjNzjjiX4mnjGb1IFXj+jvt8KmU9S8Wb4GHRlunHBoswU06AwDy6wwzs0fCj009Vqfem3H9
4QQAURCTfg0O7kYuFBA5IDJfWyA706i7/Ee9BZjKanLMcwN5YmOn5g4AdNNXT0hz9c03S2TXyjrk
JfNOcoutD+pFV72fwBlDk6xVF6VVOEdp4cZMHxn41FBwzaFFfTidHs5TImoJX5UmCgqsvjSPDCG2
xppNNSiU/xb1iPCNUogt3hHsF5HmhSngKdUDAET7KI2nzIY8b/qw0JSNI7blHXgCmaza47GDi0CV
rC7Cfg/ZnFHfjbAQ2db7MQemv3aEE1oeKa/qLpfP9FX5a44RoWCLmzbHQ5LUgMnU14EXgDvROdxS
IEMLvnSzvXtK0FBmj4x73Hs7u8EknuEpua/EPHvWToYe36WLXA39Kqkx10zOlEiIB4MVrwWSlifs
gHAOS2uyD1ExiQjzAV5RJ1nR2HPnXR95A+Pbpsn20GmYYCSYdGvwhQCSLjf+iS2YP/vbFUJc81sb
1duK3FVg27ChOyB1aRwAjLojzUcYv0qKxl0l5gGQqc/ZcGZcalVlox0BGFw/ueR4Ojh4aEaeK0z7
Z97xcWGbsByARJe81XKVWsEZeWC4lRlvSg4IaUFXJFh4i80sSC2QUuboySXmp4chxayz6svFP2WO
Z2cfDJUWm9FUZ6iXI9RT7MwGfzUgHVAqQiOuY4kZTFGkC9xTSeL/e3ulGWmvgYNPhV2VzdKDYRgj
5S57X7NJnVuFnf+NrT2qK7rkB2/19DQBi6ieRRkzrBLFy9jAxBYmRvGNw0FLkpsv8sBcF+RBYgMj
oh8Nofa58qPQS3ayjsRpJrRUHnFzh1p5hx1NF6pmbL+DV6BbLx5wBow79CfoM2qLG49lnRckzq4U
ic/2hD3XB7iowc5VzKRtwkR/VleRQObSindXGrDMb4a877uNxU46xL/L4a2knHoZRmocWs48co/g
cSMml5JGUsDThR9a82PxpcrOQL5BlohzZ1bjIfTLZ5CZOcmwQvaf4bkXVFVUwU2FMW7uUgBcvC14
jpG17lFXIa356u2Cu1FJo0gVqLALhrnGP6cKNJAMI0KUTd/O5B0emLyzxPfhfTRmXN7yef8GY0wd
gdxlRfIvtcOdF84/IcBZTrITZeAxpkwuc2RsUjuOba8t0iSFj6tFZWX7Uwfk3OBPVnmm4niCo9oT
2folTU73xdgaPdm/TwaTP+1BgPdoji+fcZGP8rB7TTAGboigQwls1FxgISi7G272qVEEpQmQPsbs
jnbD6JllwlZQ4JV0/Tcw94aCKYG9yl6z84PjJ+AdmfZeHCc7wy9ec70Smioe6VducMZYIXxunJjS
IjZiYUyahTgewMadfHcx/tZvSyodL66evp9WymWzloJNvNDrANpzGJdo1yLEGDhG+rvQFoW5cS8U
aO0V+CwyFfUTBoSXSkT5awAyIJYBDNUdhiBuDgmyTxsimTdBeRb2FzP6v8jgAxmFaKVwasxiCjQI
IRPbM8uSOayMaNJob1U7SpXzrWnTtNXJ9r9UJ/XDPXbu5eHIFMSioU3hFOeCFaqc91OOIbJgbhU0
Oy+2PTFIMeVsR+YD4qCwiH1j0Ba3avU9cVMGmRAjhaZrfbPzbS7J6EfqWDa0DoGannbjnbm0Ucjv
IDlMDsGqXzWHBDnHZUyadLAlQQgkaAe723gzSzL+fXl2q8pdBLDdBH7/eu7yWS6xBmYQ9G02ynxS
QCW1OE8XXmfEwWJO5xu5dT7G3JEyZ+ggBCpw2bzMjLBg5XbzuBS1q1dp5WX3ulTxhdR2GoCjmRDI
m870OSGvUoWNUlVjalHrYp0sdsG5OKwBJQhOsnQ4CVtiftQnjRlJVSC646Hp06iKfh313vASjLzq
qBJxKMrFqq65vJkvpdZEG8Ieq5ppt2/hVGqUYm2LxkcAlrmz9nJFpZ0NmKKxqVZFfv41JuEFekO1
ahKkHXdISXeqqiZHCpGrzezWM1L/GJPto3h8TRumV6vKPcMRfOFsMh7m/F9seUE4BUITek2NOIyG
Ct/HLaH2dMDxBjnwVteixXVXIrSaAsCRdUMtHZg+g1aU+qiuOUl31A7uyBAma6xkWoN37lEKoXPu
8jvFB9r7jKmjbMgmS3xJgemPSJKOP3bm6wH/n1mJlR4Kt9qAYUEwVyBMz4k3JN2LGPHrARXn7wvJ
x04jq3OfQxi/pErBjvEgttDq1sln+ISxwab3SUVUxCGiCPDhF2m7RcaYoBZoEsWQxryA45F13iRb
N6lTWjrKPR0H1CtdEzFWctvqBV7ZKlTqMzfBfKlC0tX29PdFBZUaG7seioWKzqwRkU4dFtB59PLY
NHYyJhqFjWYi9TjWG6fo9+0ccFMkgqfYRCvrqE7otiXKNQpOB1rGT+cDohhGgxbZJsXtvfmgfC96
TDCRs19bHiGPfxYZOqoU8UxT0C0eFxLu8K8364Vbv3fsnm9vL35LbJ3+akravs5LyDFx762gQ2RX
RXygUUw4SaAE/oMIJTtRHts1S4nC4NX0kkXwSRxPefRvVGJmRgCBaBEoaZbeHbJO3pyqgc0Pptsd
v2qDhafYlA79PIx5iLPtBgQ4/g0TTo9JnProfP5gqDAd4b1JsTJPSCRpTUY0WP6CJgnPv/E/ACgT
8oAfymi3cP4gPIAxM97JIjcH0i5uW3wrwpgWkP20HMopGJP/fTC+YeGQotE7QlEmWyuI2qbyfzUI
Rf/315B4xM9cBY+92xZQiI9/t+TRpTk2TwUAoZWYSXdNF/AuSfhBigiHpbZ6vqeaVxHwq6duZf63
AdKO8ythurPVXB0MEt8rufVjpzoTrejGF3xWhzxoXBdPl++uyaJ3qd48YmeZtGFkgSZCtQIjLxBP
mwXUeIqrHScTWtK3OSv8zGE+LPlb/bwitiYBHnwFcqfOOcnt/WPTw5cdBytArwLra2jTYShr9xaS
rAUCEKEfIEHoH5ZdmRbFsGpsc8R5mJOz1za3eEU+pDlUiK0dIvxg6YyTty3TjO2oxe/K5VJsmt1d
hHiluI8CGoDeaHtqPgexFlnej2Og8MCSvPk6/TcZwrCwTo5nd/sSoKbTs0oopkkjbWO4fYR9DEa5
+LXfreDW8Sp+oMs5HT/4OVE2LG/8q6WciDaE2OZzQuBH3LC3PJQkNxb5h7cfS0gbWydRr4eE+lRd
8Ufaa8JwUzDi1rVSiX6Tg45ndTI3XjRQbAJMTr/8lwdTu4P8cTjXUbgItqJbfO+Y/hWwnra+16yd
BfzpFQwWkF1Oz7ZfyQSYcSF2WAjLcpr5vhSdXuhu+K6OSX9f/icsLweXdCfrXb7dhi2YZfHh/Ur+
sjJwvWVoPV7NAuR20xE0vd2ADIBFMozJchSz0bh5/txq8FbQ7fk70j8oDWB2US9thAKGn/eUSPvK
qViOlz69+usRv2nbrnb+HMezVz4rZjvQmvwVDNh4TQVSBJ1KYjKrA3f8BBZx9tcDGIBAl5DrFVZE
iaOV/9yxdayd+aQ921NEDb+nYoimARC2UrC8YcCgYqQtthybZWM6VMTM4s3sk5W+jEVqFbqHBuSq
jynscyQVwa+DLO2ZQ+Dbmtp+sTOgUOid3mE7g5hPkOf4WDtg9D9EQ9kZkEYrhjsZ0ELLsN1a4PJ3
qFO3FGax7yMiaY3xL9h01KCRmV6q9e+Tn9QQc2RRdFOHOggDwSC0zz8p8j41afhyeJ1oG2cROwRl
o+l+vHo3QQhDGv5hx01eB6VB2LuGt1O1wRL4WD6UDOU/MIc1yEdu2IdIT8HR71Vy1rihqsZ3KKr4
+pfkzy0T2NFL4X72ofPRUoBP3kHwG1GPQ1ueQ9C0gzn10F1XIEJPk6+Owle9DXgA7apE6k5Ag/Sj
RNGyc51yTBbSenvxs3S9wp2pHetI9ca+1yFyX45Z+kdKTvX1b/959vX4Euv79qq0pBYj7c1YIRcd
jBWWAAtDZ8A3fNvK6uCoo+UkF7CQW6VZZR6680KJ+4AqW6svylNgIRCXTV+gD5X+TlkgXp1S3jOx
dP0kxo6mHNia833o8waI4KB3tacE8KXft4jM26yVPiI/vGRzQu/YxuNh8a5K4cOtkXTDYu0l/7K5
1ImAqXouGTbxSKcWhkHZSuS/Rb6NNwGAQTVVamdtBU+iBQQ8iXrwfuoM5/lwg5+BakbgHkAErOJV
tXk+5xfXqgUvHovsC7Aw/0T/rEFyooiCP4tFtPw1Ex8ZVi0PMGrN978JJqL97+Jhic5x3DkvCVby
+XeQGHfSJ0sFuaK2BfHidCKo0F7ipG4wP3nCA/3x0HGOXJvPJJ5j7w3Jt7Tee8X2+kukPw+TAxrY
keZ3zbLU5xlsRUZd/K/2KC0RKqbchiyWzyJuqHjD/Rvte0eLKro9F7Uo05gWv6ifVyCCaNTl7ohr
HX4GQgQRzl/PGnd/ULH1vFg1tJ2I9R8CK2NLWN3HlEie6QZ6gqCMChY5fLSByHgjOB60odRicvLx
dksAUHbwkq7IcYkdO4O5cHZFe2hDOrQ1B424njsQVFx7veRDFucsGKXymwkhr+6yNAXIQl8mdK1o
BT3vBLemS7Buo6BnGBJW+oqdEi6B45xQGsthQZS9IlJWujy2FktvEZ4UhRjXF1qoVy/0Vxl7Byy5
T8y4deBvlCFW0UL6DVEXvXhps0Ev1E3/VHVql2xuCK0hX/MTC15eTP2rMw9EP0hNly4iQttbhDoB
PIp4KaDB25ymrhXS20YnIIOKMSoQ1YI9EnEqKszCrvI4C89g5FsVgkm7adB2Hq1+of5gLm5gb+Yi
WCOFFAvH18/1+z/kcygh2hyi+7F5w84oFxcMiSkF1YMP+2IGXhADqDkaHxAxN+0H71PhD0N8+hJT
ad0ZGPmDyQbSXPVhZujNe7ByCX+NuqWMldsVANDjf8GoBfsZDA0H0NQAEOZjK/r7yFZaVnhUhvFG
c3LZlE1a0WYw/QRshTq67q6D0sE2a8CaNojc4TZT+V1plZ4MA9A/racph3aKJZmBpfefHMZwnrtN
zIzohWhPwxbZOHyIQJTiA/aBM0vPrcubaMG+x3UrorFJdvNF7AvU/mHAeFwl0KrqfRFA+Myabli6
TYuOiqcQUSR0XA4LGMOmHqNRoB1/IgTUFIMyNFZmdqdyuC2eFrRVqIEYFjAqXPkIoUpJDEx8mgBz
5w4R3TCJhGeuoUVdkMxL19NzeZYXN9pgvcO8KeSTQ2XaoCeNslOU9q99olVEzLyjdAqqrzL2iwaX
Kv4xPpQ2HHffzOz5aRKRtn4vcDvnfQXmkHcsbPps0Xu7vxWi2sGS56KNzmHTpC7QdzzBoDF5COmz
orjmKxy5tpwSZqisPMLoILh/4hFyd+6hlHImm45TfWbyqtWdoMngHvfkRu1s24jJHU2wmiOjpBCQ
SZ9e5PA1l4dHbzmn6sz60Qqi7FDMxSkJYLy3zTB8QjpqaLX4YDR/fHo22Wg0eviN85tPS9m7sxZs
+h0rV0XQYEgi4A0rmtzHdhNVcr0Nh2v3OVsh3f8XTyV8e9mf6BYZl7gXYzoX12KBM2i3TJBJIrE3
W10ECNJkqnaBlZBviPI746UI4XX3wiib4vNJCGxshNRkpjn3S12NpGxaRhOLCW/huCzeiEq9yjtX
HSAq4d0CxPFluFdWt2j8GlVJovAqTPKo/DJXcbwcLyWZ8SqeCUO3cg2Dxk9n9SAvY1g//nfUNAV+
utLqVaOZx4LUUxkBKufvs5wjNfpV+9doQD0POyxZma889zFyfp9F+HqfP54D0ozeo0LyvaNhey5q
B9qQMurBDNb2gcaVFaXl3WkAtdFcwyct4g8Tqx4OS8rfvY5FcWpBZGEEOwy3QSXQ0dHlks69Oqko
ygy62MSA7dIZWKfbNfGdS2nk5qfVOQMgLldMpOL1DYPU0RIPtNTqOkfL2pIcT6O4QxNui1wEGlOu
aWWNsx4oBZtf+02cgayoM+ZvrLn9b+NmWL6wF7qdGoC96uqYkKyT1/ZdZ0+DlEADNoyu9k2ANtVq
XZUKqks58HjjRdWD7eTVC5CF9j65lOX0cLQO/p7pYfZCFVG2/Va45ndWXldkr9rENBuNdbKsNMuK
D3MgkNKP80Bpyx9hVOW7S6vcC/j/HTHyYvra5iDUyu5pu3d0BG9JFBplkT6BaluF/vY8Gh5F6YMT
ivZs0kp8bRk83WQf1ezkj+P/cSCv/22pLhKRN3SR8AkNF9iyPSOfAMaw1saOngDofmNLYhMB1oPa
/bZOR//JAxSFyIvxY5c6uO6VVpCFL1DuTdPXtAFgJdbI4gL5dxTBUVvJKz6ycklTL2WMx5pijldQ
6roHuUfIEqUVDvRmeVLFNn+UbvLZLV0Cff9umelWe6tAL3m7Bu+RBACox12yy5p+MBkaBV3Clxua
jEMWrLRjzHKL27TPMu9MuXjJFw5lgJOWOqI/VuTRUBiaKL8ysdZ4RzRh/8cXga10+uEHCsTZSfhF
R8OvnsyD3qr+8ZdaNvx//lHfEofeUL+16XVphKVzsopijjTry/qjfrj+u137RzKUCOvAFPo+7Uof
szJ/TA+FznsIx5h+hvedAhJlvv13bP3F1dkXYaL6jtIadqD+PzIMnHSkXj4lK1KD9Mtjm32EgjTi
S5cqaawM7GbQOT0ragFC5Be5huKZzmJXGzHcV1Hvmoe8pXFlJrfMh3a2bLurTkmUk5+LAKDTTt/7
n+1DsTpnIcCgpogECWM4iF0zOwQq9oWOadvb1NHYkmVhu/cQnQijd6KtI3ME+JRg9m6v9SRBQ7VH
rNYSngufNGD6W4qJq45kacP7Au8HJGPrMSdq/vT8U+Co7SRwceX0IP4NSFlR0tbdD8D0ODDeksml
H6HuxnrH20hI3XITr3wPYvivDiCj3S/0f8dwbIA0k2LiIFaCcvUGZkwYqePMSUq7skIeq3MKNK2D
E3ARjsDtPAwUEWh4byttIXpFQIhmNosLaPDOZ/wbRbxxy07KUyQn6TL7CMXjX5n+nk4ezDtCLWSS
EWoMhaVV/AfWpWPfd81m0e2TCOtNkM4bOC+rRoVipTyXVI4dSswuRedijhSguUJYkvFnkiw1/GPO
LteKzp3YiyU8Fe/hgb18VKBDyW/iYf70ZDCVvjPSeTcYFDqJerTJKEbB6GExYCCFwIP/nNzsS/gc
QJb060GLSiGvdhJMX4S4S4dfiZq0v56KjgingsVNtpxAMmc60eXwSEHylFxbG1CiElA76VAHrsBL
FKCEbnrOOE6w44+YW4G7WoPHAOLU/0DYxDYKY95Z7AFGhZ50oaa2xkY8v1HaTW5BP9LlxPUlIc8g
UgOxifBDXPjpX0yXtaLIMhNry4PGGh90blWQ9+c/Kofengv3BLvHmURiqMJHQxwATYLpkNz6xHvP
dDgQwTNAAL3C7RpiJjc5c8iw8opF00GC8Xs0+KBEbvEGqSFwgc3b5lUhPObbOoVQoEZcXlgDIrya
imKZ6OSKZ2PGxPeXfULNdFi7a24mjo4yXw5h0H3l18z0O7k1TVgzqpQAS9DrHDLteaUTIzIiZyoI
lXXZt9hwHOjX5vqdJSKWgsU6BcxlG6rkIloghOLoPlFSwa8Wvi9VhH7l18zFA03bwSXJ+p8kJb0G
UcxgJl1MhbQQhTrhDe5u7L0IOkPAVmdfznVLMa/koEoT8G4MDEBuySWO6BW9aIX/n+VfMfZgMMWx
khK6ThA1Ko5zba8+WPmzyfot8Z4tXQ79LUrw3QoNcoYvzP4ryYVS4z8TZ7LUutY9GXfvujrxSk1F
oGpCRni+vyEKfHroX59CKRM7F92G/H9Gdbv+tZlmHCUqSjOsuj6MjvGDWPB/8eLOUjfNf2Ep1ZzO
6y+chUrq8VETlRP/eUtiksF5iMp1auR4mQ5LkXgtGIQyODHTXb9UXw/xnUGYkcee2daI7/jrUioH
1Yq7TA6Gv0UCRvVxCIkA7S5wC4tltLOjm8TicW6p3k8MrDIVsVA/MtczX8xGp4pQ71bbQBhn2Df6
zASTQOD32VPpulhwt5DiYZ0BlSG806zPVaX03ywfqEXPTriH8uOPKAMkCec8MRXbtgNxWQ2RDk7K
zS89mpBkGlBldhAdSd17/TDJoccmmGC9/W4lZqxayJppmKiGfD3+qMqKTSlG6uTNu1eU3bLj2iop
DFbdOzOHSi3HHvY1Bb55rq/RBxcyeQllKYfvdo6UjusKtIUm8Vjcl/qluz4p6q1CRU1+p5WizdeG
OGHTTaPzpB16iyyQyn3nPWCvt+PqGvUfYXd45pYRxHe2t0ei2+Z9E3LSkBykI3/9jd8wUP7i3I2Z
b1mqlyAllz+HamuaXiDCCqdKLTj4U+uhL6hOzIox4IFrpTFzZFMcnJgjU4wqLNDloHsj3cdR4sA3
HnJepshWr0e3urOXidCEI0bnFBaE0G14/FS0JOpxRoUJOMLJIfoFb9BQwYlgAgD/G1O5NV9WUY4F
pyeQQWte6ebMyqpRWMDBL5n4fBoZwPs9ZUWmnhFEM3tHwfF6NYOm56BAaW6gW4zMDQaoAy6tlKbJ
BfzKh8Z0DDHipttKxabBK0UG58P/tstmUEgHkvmXGsbGDBnIaBMxy32iasxLmFuUkDkFs/Nh/WXi
NJzQl+WjzFHVGDj35iWA7rzdy8Rr9/CoWVWqka40gTs9N0EW6hqjTj+0/YPXBaFgixF5xm27nT4i
h59MLKASZRHF87hLYUtgB3zarZss4m90pAsqb7fgatGhlKVoDcmeUWR2R4NOx/uMhpWA1oag6Caa
DDQXslRcbd1SshlSxxqE4EYLjsZSG06kmQOszrEeC0Ky8HbbsvLS9ZEZffRjugtZUYHt2Kwsjq2d
z1Fn+JyoZg4LbNpuIVi6uooMrJ1abTLNSm6eV+A/h6OJIvBcwLB5mNS0A43CK/zhcHrEPOtlBlEE
UV9taULuS1MDO9un8u1QWkL17KD8XhAbYCa3+aiTEIK2qJWBU5/WA4whbEyy+2ngXRFpfLlL9U4a
uME6j51qIiSMx92sfWFnjTWPXp0Neikm/9y9nvycMbfcAm7t6RwrArBW+Ltif4JaxRJxqONfvJwy
ABiMPOzNMXBSXXq4jpGPss9H+Ed3Vw+Ji5Y4qd2v4pzvGzSY218cCBSsljXIkdSjEStDerlld/rr
4gt+a1OYBjRAtN3Nuomu5809VsyD63RGTzWBf2nfhzpOIFh0qBSA3J2Y/DprbR1nDTMBvWFwsQLK
EzgFZvozIQxVCV+Wz+hc2V4k/aNXRIKdoCPQ3LLFAQxPIA0sN7pysrYsDfH8oX+zFmzpCLsk0jFN
yWbVKbbBm7U2ZcCzeN+XUSKPtJZQw5dxYq52Yj9wZ9HWuaaMQQGVafGjDpHqWCgxWe4+NjV6zJda
CQigfqBMWW+8L7fwBBn4+UOtIvzNedAZ2NzFNOU2Vh/aaEuZbVEOWi7O7prnRR5HwF33UYSMGk46
gJkqOKut6BLGQekyciH0UPoYoFYJmKuok657Nmx35Y4MYm8VAbQt4pgy99Resb+HTEiOs0QgDU9n
2kw822hHZ86pu+zizF3FuyEI7M3sgHxF4W9t02WUu+48rW02OsVCgTeb0qSpsOhLTE1jhJbrBgux
q8ZmP+RHCanZq1H4tsr3K00Sck3BzqnMEJbsyd4xuZKpU1nuoOcS/qIW9ZUSBU4yxWtOlEVivLDB
DP3tidQY+sRCa8O5aNIEIvGtAzkntfkcQZEg2zE6j4+v90fhfbmp3iOnsaG92OcXBMk/XtXvPY43
+jE8b0wUneQ8spKDe3zoIYrI+3zOnn0IGtUaI0LNqZsJ0K8TMHquJ7P6nMmAEFRPdJFgQCiUqWrT
UZBVpGbh98tkCY7mVPyTaRjnGrJletZ/CcJAQxQlUaP8uUy5xp1+C5vm+9goQ9JdGD6Mz3du89S8
R2iLrzqpmtWe8Otfe06NnR6geoKI10f5MvFpGSLATVqCHB9YKRATYhunwxFjXyFrB6gyXUwH53JE
AZAvfqGXsqgt/R8tTssyvPpQB0rS0IUNS+LJ4+sMRNBGVcot92x7zbLMwRz4cLrKPdpKNjsbaVt3
vrEVMs6KlN/8ZCGCUpQPnAWtN14b4bk0V+SHLdteVXB+00ExAJSVK+KXSurwVCPMEX8mPmiJEYuU
eID6n4tWB6RG+DIJx95onHeXaUzPYKzLrarqA2fnzSlDJ/GEQYbQT9+6we9h4JzO6RGAu+jUs4J/
c4YMD8Q1UMMKbYwFSeujsFhF6jJ6odBqyWjQM8p7sSLr5QGT8r0kIK/7FbMYki2IeF+8ErXuAN2O
ifxVWD17tQ2GXi7Pf3z4iZvYAqpog+TYwF1npnRsHyySRjt54GEwnTTRZB8ZFMhMxb6azMVU8M65
///In5M4gVueZL7mmJhe7MaqWLAEiscqW8fGIO4+rD9fILWvlqy0HtQfKHX6h0bo40SfQTwzf/Wk
u0soWBvMS4CYSPrk4Kg2bOp5IxzcIT8T+ilCgkm6lIPwidS3amPCIevUW6oqAsLaZ8zHntYXrss3
MKkC+Q64gJXcaPGME09UR7oShz87lUi38Aabb2P36gTQoQ3X+q4TKntDXQgVGMGcp/bUbdbI18kP
Xxg6/WpRdgmyY3+BlcyIvH5eMtNA6EVYAFAe3w4h3+3AnXNDHeddidoTwD5+1+UyrsSoggBYe7ze
l1MtUsiEV0NbUe9+XrLtxFu9G1yUC9LKoxb4pYdrus0jNXeTpjnditGoszCh8/w1s1SJ5ciXmZeh
5g16QnjJYx4S1hM2ytjgkrTBkp3t3Ozg5gfITDv7xz+pF4c69Fxdn3wWrpLXu+H6ADLhjKrGNsrG
PoXuGi1AhWxGHvruCkTNcxw+SVYxUBgBcrHsC/r4lWW8Qx4mrusq0P9j8i3Yn0i79LQEUn8t5SXv
LOPPD9py664Ega9z/EnHSaxAzMB447otig7hyIK0ippSLg6uP0TuViTwSdTMeTeM6OxLF5nZ1XFK
2w5FdqQur1YTpjTzZIzqn3EF95ukpikYVi4xcxzPISA5uiJZDQmp33+75YeBD2ttKqUew8pjoXr/
9fHvudk9zVPKjawSdMmz2t5S329z1D0rp82or6dh+980zfUPrIojqGSBvMbXQkzDFxWy61UyMdTR
ISi1hF1xdCdn0NxOP0ZsYVpqK41Ilm/CYxRpq7fSJLIQ7TgKPK3nLTbwUXyiIREkMx6PvTGD1CZJ
411gMQlQiJzF4iXQAPjSEJq0onFZM8qBn2wUJCDb6DEMYE1vOhT2gYmRR1KXB5vVa0YN5qkDEVxx
oSv+HXLcoUx020jpfrTS+irgw/++jv7Yje68YdjEIKc0Ly7plb0xMukKQ+Oybdl1S2qpMm2I3U1O
llMKUd29VW5ZRtKPsrRcsnk2bKbPogaQE22ah6uuxY2//UWKd2gbLsxXUz4A82SxxiPJDQY+AnMR
iOxAp7ZYmOO17Gk7F4DlW8caschijmzVsUWNKvtR4i+knrxlofMMHXl+3vXq4PVLq5poDJcY/se5
VQOkNSlfJhAeWiFS4xX0jc8oBRnu/hYe8ii7UsccKuNy8YQIkQJUIewOFIX6TnjLSgjGvVmSn9K3
OyOLjI8SMw4X6oU63NAFNdNTiGx3g1l5BhCm3Wgg9QHyOrAlgV95Bfw5gVBSoX2R4S/1h5JlO4qj
FbviXRMQWgcaPzSeqo6MGsEZ4k7Y1dSlUXYdAEwcz1c9nu/hhYrT02SAwb/geUD3bHJ/hUBd56lP
e8MWmsq7YfM1DzJD3Twn4J/JL5InDbGlFX2pLTixjCOwu85Y24K/rsw7KWOw7bEa5HMOntPAzet4
rlGLt5ovNwCDQpiblTdklZ2TK0O5awePItlqiGqqMVtzUd7lGU1Y0kpKNP8JAR1aqxxODcB4KJxO
VDDzPLLz9aG+8sUS/KcEK36NLxUwScYMTfOiCJ5kWRJ2uzHrs1aEvVZKc3a1lyu3z8F3vt6v1OYz
B0KDDMkMpy+wKIvpo4dNpyle15OrpgP3s9XNHVeBg9OichxKwhXp7USrbwtJpJ2Uil1eM/5wxNvI
cEwprjTZgSffh4Wq1JxYlYvppuFbB9Ani/5qZFhpR8cUGGaHzC7xRt7sTY/hC970zG8Wtg//9zSA
mjEkqidMz56c0hCRaKmx9oTdzHagEKOz8CA0hqZ3v8h9CRkWTpKskWKSLi2Umab2OgrtpPjISNb5
A7wfqhODC3ZD/He0TmSMEufGHsiKegHqTB19SOe7xbo2tttMxrX4jgDwoBX1KnPRQZAUEI2mfJmm
ElTZF8OFmrsfFAqrRNkO5Mw8k6KZtOF+1bHbtv/l4208jLTe/zwMwVCl01mW1Yzo6N6Rq27QMHs3
K7/gnSC5lwiaTxzX0zzr6i8ic1kzEzX/fPyDNk6k3Zg1vvt99keGcDfaURqRgI3ytlinkMDsPNFK
zBqKIQ2LoplB3jqO+PlSY+OShEreaX2v7VND/B3+xgpAo4kTgl4nyAEp+iftgqq/9NCAD5pV9gNI
iuTw0hjqTXlMmRs2ajXOqtmLZbaTl/qgCHdH9tfm2dg1ltpMHhFCOJh5RsyRgeAwfq0mej1QQXhV
EB9ddxRMm/ePInXcPSEJvNSZBeTccOV7NR1KRY7UOZ3Ntq4z9KtJTq09AXXHjqr14ICyhkhpBMNz
ZZQRtxOfhTFnjjqepeFbrIMESLk+hEC21aDVi8liHHsKwRzFzECnDG6bxgZxR5d19IWzhhyHZ3Da
6/0GfpbwNK3VqWFY1hu1Pj3mSKdp7isv1/rKGzTHM4xQHrTCbjbs+oklyxkvTor5OF9b1D8I/qWV
2K2YvRrLsikuH6DuzSc8w9dSmOYX1+s8z+G+ivSSpXjXf9LB/quwGF235NVRu7O7J+SjJrx8Kxg+
BHGG1hXzAB5H4UG2KL0aB3exYCpOc58hTzblZNAFgJRLJ4nfCrYojzJ57gANMTuzZ6PaEqqkBRtB
LAvN2pgknWtNhKe2K24wxGP2L0yVN2Jgadz0O3xnm35luXidhhJfpHeftW5v2mqgs2FY5YEKcKm1
J+pH5yt7+ry+/TDUCqFu9p/Mc5gmEknGdTePkWQpyYRXr290LuHQGAwqkXRW3PxpuCGPzHQjk2Cj
w/sVbTe1ktOqo1a3k+3vfJ+5ohMFW9T9i0uaXn8fD2TvEGmowt9u9DxYS+M9/4Ra8cOi3/d47b9l
H2BHLHsLI1Dlj5/v8KXIABVDKugMxZsLMOBD29zDzMdJTazMCD+42OKtaaP80k73XsHIYy+m4GXW
BC1SEqw1I1EuYWRWsnhHS3NJX6OUVpZ9/hSe9n6/Sj7ZupR4Z2wL7JOY/El/tGaCVM57OBkFFYhT
0dvhbziGNKZRnSl2AK0pri1/QfCUbdTckrpWgTaLoFTZc6B39EkhnKQGfH4IYyKC/XKoWAYPZ6pd
WQn70WbH3rKhdFyZmuIHojwpPQy2OiprytOCTWsqJjujGrZVH5k8wcsZ81N1jHbjqIwcPSipEXhV
qMzqjsHojHB+Z9Fn4Ji5lsgocYzi+eDvCdcp0d9fI6rHmB+TDBfhSR3j+2jNck+ZZe4UXCjoFDhl
pmD5C+WWttmQfxpdwCeuyBYTz5ZpG6wxwsPhUVsv8PpBESxNUp2PhToR48PmIoa6mdvUTGKdZNQ/
npgMuRbkaoYAJ5KYkzTFN2JMNDngLVHSrlyuoWqZM5FklyoBg+8ndvAXJYVpI9JxzMZu9AgPjAJD
/IIB41whJsYKT6C2RC9oxegjmdcLf3cBpxYTTlwh9e9IBnshztwb4c/azG98WujmfK/qfSFCDFub
BasFehtbC8Ps13SrTOtWMgd69kF0EojaPMKQ+fy8hrZ/0zv7mc8+wDitOfd1mzfW+ZnYsxM5Jmj9
96bjh6N84ZORNXDOD8Cwa6CJJWmgTNXx8q1Sj13pCCr7N3S2fGg/jlcvaFW5u0f0OFKSZf5gwpc2
o7MtzPrzJ3uPMskA/nqlAh8M49jRvL6QKk0Vul3ax0lxwaAWVqqT2Ow0i7J6a/IQMQPdVTX7T56E
J2BYmxaJOqxNkGkgANQM7PJRLqkjROKYOz+wNBSZuxJS5SfMxaJptRuWK66/+s5M9VDdBPYBwTRw
Xga/LuOMrsoPF9rJwGr8vIDCe/Z50Ontn5RF/dd0ZqS9nw9TXTXXjZejgByJGdXmHUjnU0iXwbFM
R4gscANKjs1JOmqGLaSxr7Ti3kdW7kWvxz7Cv7D4zhjKDPsACNrHqRcUtMdMYMzd91ZybaD5vw47
newqFWXZ3FRTGjaPmEDgah2facaIaIF0D1gNcz1vLsa8KJPhzu/2xRdzAe3n6ptNcSmkq+GWb+LF
BL7whcI9nMT8x1eClJRY6oAuOB7oPa9+1ygOP01uZihDdGaj+BP9f8V9tYJAUO+UViRfD569cS10
OtGktHUxfMEAOpzKxqfsel6IFpg+p/OWBYX8rMl220kWs8yoUjBZ0wXCrfaJGghjPjBBpKLguXnA
68thxsvaz3eeqxTCcWflnxxhMNW1fiOcZIVI8QvJaMcKw05lVydpG+R39jDE0bAg2ICGC4M4ZfhB
chWyKCP+Z+d7WYqrFCClz3HuSZJNWB+K3GFTUseH1t6i0LgOiLX9/D0ja9kWJS6aK/6JClhI55bO
Xn2d1g67b+3tvp9ehIIGLPVAl5EHXNubFZa/FPQG4uaNA4Hz0bNHZJHqAEXd31W/jSalKbNM+MTw
2YYDoA1sU1FR//bAcxwVtxUJ6/csmvmPeTIq9/gKoC1tol7x5BSpBzBYSsCp5FkHBKWZ0Iprqi+p
7SnbzjHsRCUJYcEels82/pMt9bOQ/7q9LvGRNYSkpiaNOoGwcbE4oi/GVaw8bCb5oScudibFyff6
IK3VQiVPJCxQsIR0wWoinePOlKTFEqCAxUP1b0dgR0xLmJ80zSBmF5vLHR5upzOVCDCQqSxh041b
OZRdL+bvfs7547uqmaWAiKVojlGB9C1QNGn962uTsESB1K8/mnzx+oBbcer+eR+lSNGryJdqnRYY
4eCZwl7Xkk8r3BKHSiF7ex6huT9/0XD6xqb8gZ7biZtMGVVuNGOISdDWpXoDMPXlQBY4mVDSQuZj
5jr/SBfzK5bCJRfpl7peWErxPaS87hZhIJBQ2KmNWh0JfKVv6a7ouxHafncyQleLqjNKS1GSaKG0
a644FJYfu5zvy9GMIB+nTug5QviRbq6filGrVE0++/2Ndj50wD8TaAVINlpBnulgSwJor4ZERgaL
nTMRZn6aCyBwydkQeRm9S1/S1uwS75K3LIIRT3RYBnwPW25Rye4sSFKzXfRfpc+qSGAppKJV8lFV
S3LX6D7JxsgrkOouEbvVvxakb/xDt/OZjJUJeS3zGTsOwCo8cHnywagwceXIaVJKmH7MoO86KcCX
aBnZkv2rq+R9szkYy0jGkQThKHZOEj2bM7mUyyPXGhjAS239/LcXEB0PyVNVJyzn5fcv1JO453kk
WRniYO94dMNvxekLMAkPDBgNNOYZPrtslDl9EzpnL1a4011G7x8FVUmSrLTndObk6x3fFunsbl5I
gWMd3lTTmCAPze5Lk7I998F1MlK9pnT8nUArXdpTzwa3LlY8IRywk3m5cryc/Jkd8qi/Hn5av05D
IE4E1xoPD5d0t/xup8GwM6BTgoOfhIos9JniSJxMmnpWuLMW86etQ0w7V4OKm+CnzzFdy63nQYeJ
vU9zVwTlavjJWvAlqQSO2bKkaVegVc5UimUiUDc2NgHueEZcjg89bVgGa7B3hySXu6+XWMn/lY0S
5Dd4qIuoFoHImxmyU+RC/jPhkVEyKuyMSilrTRdiH4HuxWCqI1HkovCiem5xNRSLc8mDnxCSCada
7L+NIB3p0aMEF2H2vCdOR+sqL7tZeVGsQIs2bsMHB28y8YJ/tAYoArSiWZbMMjo/aWo9FOnaJgft
BM7bI2EkxWLXGnon2Z/Q+hOM0kkN29tqo/4NNhOO1iyECK8wbOc4rWsaPqz+HE81plHkISlXseI/
OsD1H8cOlu3dFBpV5TbjRVmQFqFvRKrtCR6VA0q1puyRZhdDj/VfL5Dfz3lgGd36AdUdNOIFoSLY
4yeI0eQDsjFFoPOxiqfaZi1/wURvsYXwsJMOXh8hzu96ZXlDeQIe8c7qkTYZNEdA8EbQart2o7A6
0ypVDHD3Xo3SNyYjZVMd7pCQBp5TUSCjD/DW2J60m1+wPg084MRFniTQGF7w2YHmYTk1ysn7Oqmd
veHPYJfxsUsIYAlPjX7cCwyqcZyrogJRJ84GZ5zBdqBfIf57buN0gS1Gppeh9KqVrU/D3qecaQQT
XnmNjkaSV+pDoa6diAC1yFoM4UAcPWQJPeC+v1zypNylNYHDNYhpUvxQSoZ1Xi/VfMUXZkk1QK2F
Yu173LugacxqnWDWpumCAu65drhhotCIxN5Qsnx3JDEQAqzHG1M0zp9dCHtt/ZJdVH2XGCUVl11A
bWLFoe/KsSGZQGDpnMIwFDQSdQQRZnPiKeZkgr05Fzn2Z2vfjmN+vIuWuBefYa7WmuFprZo/kmLc
h7Y5KYBdsjwAwdicixPwRwWrdEHc5qMD1ZEub8G23dC2fG/3mbBF2aDp9xdKkTjLwVi62VbnlJTc
Ipl0x6k/GXW0eQfzTXSPHjiJ/0psJE97piKqEtJsa38JpCAILdFg9E2KS4r/OG4lqHiQkHN/QJoF
GZZPL3vCZkJFl8DpOAaDdmoL4jjb0pYhFStEL/0c2DYeYk+nsnLQX/AQP6nMMheJDxAbSibH7BxK
MV4JDiEW9LHEihdgFuTyX34xVVryUM36RsJkZ0f2o1Jv6xN77f5suRQ/pC4OgUqqYIDtqzkKg0Zs
6xJOUc6QafHETOr09GlL1ugYrzZr7O+WRrTDz1az8gfXkNjOIgZREqzcT7Ittoy0KyLIbGEbiKkQ
kEQ4kvbFGKAkH6a/8CFTuoIZVeQBUWyMP5mODJ9cVQL1q4dPiR7Q7P2rgolz/2h9nEm9EEVOCqaL
kHKQ40KwKVubxSWH/614dTcC1kXOWTTK8cPyat5ejE5ONYKOUOYjOe1WQeDi5GxEEbBb6XbG1fz6
usg+yAzz3Ql7jshDLusgrisSGdSmit/MYSKgzCrUb3H0Yc/jweULqxxfSiJcFckbTzHy1faODunl
HV+Z/bTdur2XpAUmKJa0timf2a5kjZTaxdusXUOgYKCBqE+jjg8PWUNH58/BwZDGuYt12iHlQ5nf
jxpHM1HCC2ikhplS7SMq0IPYuftc9DKgLq6xT5xU1oNMmM+Gw0U7X8OLf2UvN1INL19iyZnoJrVR
OYwQzcKBGJsDfRCg1CjnJmPdNaQsDeZ5IASYmS0ZxFnj8AqE9dL/szhv65DOb7jQaLRoEL/JqMW+
jKMZddqC6myb2t5bOf839x/UeoGtv504jia2jP7FFHeZC1pi498JFfaas7kzwIaHbEeQyMCcNve9
ch3l1dynmESg6DysvQfxfNvTYAoRWpAaKghdy9kbMn09BGGqqUFas/88ComHy0C2JF9XPs/smKTX
KEmiJyr99g6PgIj6XEC3n79KLtDosCzcKwE/47DrUQyByoF8OdeejQgCaGEmDmJ/4H0uTvYL9U6F
SSDDe7fIKG0PnqS+uqVAVOwzn3bEJsfw/8qEaSHCcGG3MQ2I9oQZFSDOX3i5cTuPUR8q3fn8MwUm
mz4IdnjWnMcF6XZocSEsNPo5u/4z2AXHCJz4ram0/84OrNaKo/9+XynzPkLvyTSoO73vI+PkJNLZ
oy4hac1W/ZBXalwBwUqh4KFGYX3xbX3WALLkM6VDhK64kCuyFiWs+Sk27iJRZMDelSxURG2USsva
7JeBQbgyU+wKW3SqU0LOQ6hl6R2YIB+6DWEM9S3FJQ3LcHl/a0HVazegGFrt37yR1l0+5W41/6UA
2k1BsubcTCk7D86lH3VkXDZScolztuvvLJXqs/QOiqKdFaLUeJlBW27lh3VCT5a7Yu3ipdt8d+Be
UClcqqOyhw1PDCM4Z1hFSl0wvo8JlQwUC1kIjM4bTjfd44TqBfKO4nZFtHYBrzB5FXzn6U/ztwX1
BYkN/51o6rADlNANkD4GSAitEeNJmhph1IgRWxQK+F845xsIbrPE/JXiOUtbXH1MUatUIrDnYmak
yXaUOjcbmS03pLf7tw3ptOB1At+gd88DzjHRXf0YVVRwCWcNEzSuBqK2C593yzWZ+7HmkF49KE8v
9ixBAOIVyG8kr3VTfncVwBsjMnScAeA8iaxvxYFXRLULVEcKi2jtXC/Qtpa8ajiVkRntIiQk1Tbh
98Qd8JcibGZvGUYoFS8un7pp/JNw3N5HfF0djE8poaI8hh/Nm53ujZzw9UAapz+8yvUnGc81PN5S
lVg3dCRkrmmc+Q6cNt5i8eW8YddguZbO3hngUbjmbIZhDZtEISAPD7z0AoDMb4xzbUcEOjeozaM0
4LZcSNGdw/WH9pMv4DuMyn2wm64DiQuLjYP5oNrynTnmoRKReTUdi8fqIjkVn9Tx9DvBhfWHzkvv
rGQaSdQLo1vry92LA8CXkXiLz2wOgJxOnTi1nZwt9eV4i1WoqnVIdZxHRAcetFqOwGxlrk1NCqJF
NDwACXVzblh0hCefavVgPgu1tLPw8mvVY0DuHdAdjpLTriNh5BhAze6f7+j0r0qjQgKu1xdy0v8F
SuxUM6abAd/2K6b6M7T0gZsTUjYgZvhSUcBiOtEvgQVFHNXB3F7qLaTYv2ThBKwhLOfKxpqrPiPk
hF9bUQRQivGfRR65wTaSVo5DZfRZXdHhQoPzCpY0W8ly0UTebgmxWyY9Z/gOQsBKGa7poBFQ8GPS
QTyTR3JgHRTPsOa5sQ2oqEFOZYITJlGkvbSMSIC7Isq5ICf1zMRVw21KomyTl4v2h6SqGcZgUNY1
1z28R7MSLJ80qAd24Mrj7kUmzdXZm8WACL+wUhKW44EK+sYdC68do7peYvrDwAnKNBKIA86hVA9S
Bc/qobZzaD8yHzQmsm1GIpP6pdCv2aWzd4aETAIT6I8x0Gk1jgH+We8wc0q6YbUr9ckhn+pV3uiF
3RmNpSrg+0g78MNwlT2yzSVEPTH4jbwixnpHelbsp2XV+c++YFd4RGaB95gvoTwHux3ZLh1rUnwo
wzkVXfbe+9GS8UkScPyfxJ9ZLvBt/pAm5xO0F9Bg15DHq/SFew8CMauRKj5LPTM/2XWgXZURkIJJ
n+PKRkcIltpEDUUm0v1D7Zj9ssZ+5ZTdWhlJ2HpysVzgU1R6VNYD8K7GL3aXC0vuoxShgm5Ye0q+
gXqT28/d6Lt4b2rjxlGbYRxhH8t0m0lm60xy1YXadA24NIoZsXbUgJqH+1sEZoRMcL1qfIX+99wm
qcxplHH/ewKdzcGd/PMfQhzJYlpYnxs7gaiwLzjg+Tfs2f2nH9yTxs4CMdZrizeRLH5uDLskfgrr
lc48/YjBbeQatQGTXbsltHaPM4jsmyW9PGQt6SOmWvc2HIbrM+1sbyOj/2sY81K6R/LwvpI8fR3f
EKMC1GoZ1eVq93tckVnQ57vcZ54fjOt/m7DGmEQQkWAgP8cx6mnCI+zjKNWlxlwWgwPQ+fZynCkn
YNhLfbe2+LTi4rgxslNkTGQ7JSlkqXWfwECeAjiIrwNwVKGT/WqWnrf4F2P0OQsq4Qzwl8piep/3
Jx1ZtQ7K5y4j3181xxfuPVb3+hHgIzinq3zZOtQSRGhL7DKADtbmCmI9+fSXvwEzFpyN01qwdTbV
NaXbsihWUenoDBA4Dr+imWJhzrOkd0C/DiF7yYTn8UoqUtT4b+YKY4llNiGKfHWbVtMopVfW+Gf9
FtsJ7DEgNFKKn+KeVLeT/LiALbJCckbI1zH2mmBn3hYkRhbS+NaMRb+ANGEVgQ8tCgb6LKE/+AwH
ZBrjIDZ0/uWEqVSWn1sZnNiGDLpYjBRfdNwUCPUIml8zDxX1WYDBu2whgiRpNV3X+o4SWYsXJak3
V1suP03f2HxXJe5b2HoQVbVT036Iz0FFo1KYZ696NCBSENvoWvPPqigvFzmJHFKdPoJDb5Lk9EJr
JIHf/TFrf+EotCbRp0WYtpwEFgNjLYdagSUs28u/q92kd6Zdbnsg40A63ZjrZmZAa0Dueerg4M3t
Y/uLhaXkQ//Z4nCbFu0n424ipyrHIjQiElB65NqwFZtxXvIiewVa6ShAUlCqMvonhYIa1oi+ljwx
FCQaMziQHqmQJlHjbdvZkcPxni26DAIwph8awRsueY3DAjXmAPVNt86rJnmIUuReIwLvvlWxqmub
c7c5gRs53r3IEhvFKYyRTmYG1rrG1tMq7EYvM8LLq3btPKITVrg+MTQgAiZsHz51QmHRhDlgqo1f
lPcoX096uvczAu6B76bTCdNQQaFyAafN8qprzUoCWvxYfZfCoecDVWwZHRYDWmpQCtdWsCAF8/a0
WWJlnSm2hHdaB0Clh5VygW997Z0BLeC7jInsn91orMK9W+qaIXZ9BZvI9q224qZig+uFxIOSvDRX
8QZuZ5na53/bGgj0yU4UUEPbSeCkX/Xf6FUx4wOqWmHXi1HRlRy/3YnEfGFmzv07SfAm4tjUbJg8
fvMJPpuI2XRDMuOJc7I9519DeLSY4rwoYTbKSSwkyy8c7FqG/nWenDy+Ju2A7rjz3g5dRA9rG/97
vXKIquXoKONxQK8kbbXc+giqk3gbm9d56yivS8gLqus47Jz6Aj6Bj+RJbmNovkbIaQ17aZ9eJNE3
9+uJBKyOXAOTF5ARA1kbSKcH6G9a8vCpVCHPDmQ+E/TrJamqUKV+9Z0gblHq2V7LPYjOIcn13rmU
x5u+UbUiuHctQNgBe41surcfRQ9xM9/94sBrUixJQnDJTTBa1R2kQTOrwvN7ZWflj9PdB5NvdEGa
MpRXi5g/GpnpfgBdgnGANDOdQsCcdcgfmGM+Y8Ag8bIJYyNiRhjmMbYP0tg2Q9VFwGKsD9uSXAM6
47IPcEG+2F/LOhpsY0ns4rpXFe+tx+Ax/ybaqIdRxSxUVguHW2vS67GdQMUrgaCKFtGEoedyGaJI
mK1S3M3ZUJAGX0+R5Kkd62YnMemvDN1U08f/dPbxzvQrkHoJveQUp441KGVyvS8z/Mk8BfYGqMJe
NRxzLC/ROTG4rsBxz2x3sd9BeFVO8itTfCS46SilbMGRjfYdZH0+b4xH4r/x33S2zCy9NC60jpGo
2QfSK+HbSKqGz7x+XugdUs5/85L2WXOqf6dobApBfUJ7okNpn9GcSih0X/HAzMo9ICecQezXb3v0
U1/iHeJLJ/hxyVfhF2ZwJcMsnSzRbP7HvCmFTMGqioD867hkFbgsyMJQE8HnYF9o3GqXIxRirELI
/++Ciwqj1ZxDkiTxXO+1bEer98xKOFFPPFExe+/zAhFWZ+gXU8eCIWVOalolU0jETqPC9NZHTM7L
Exf2fWuQjCLYsakdV4EdrC/ZAHj0/5WTjs+T3bC3q7wE8E1dGSVdLWImS5h6qbj8m0hf2se1OFwr
QRQen0Fi6PFDWD7L00xslq0Ij3/criy66lQD6u3SHU+QHippJXB4W/qTGAwxE6d999H9yR0t6usm
cG1iNz/tmMoEWUztWfUiaazUK9bsy/KWWG8qXlF5S5yhWKiNdJfIh3mc2UxjFAUX+Kl8puzoLzV4
tKlC429XMEsiyb4LmEzZGHyEUQU2A+bMm2Hg78FoQRSKHz1M2BjSb/w06QPsxkpTAL6BUk6a6CJ8
jU0T7UmSWItVJwbMgIJ0gkgQh/iHS3yGJBD9+9pXf2mN/qnIHgdGFtvTEiOMzt57dleTiM/ILKWJ
zzLOyPP2WkSlgnxJ72wnol3kX1sjx/s+jP3UPQOp157j3/N3pGVIiPlI7uN7QYlw36l2Aap9vuvt
SPiRjC7U50V+R4MaNumlG7MHcKSNKww1xuvgOTWPURQeuZvg8d7uLVaChujBRrKCEUgGaZSZ53uk
cJYliIsd4bi52t0u7uXEYrSwy3pYXZPn/Z3h0/xBhdQiKvFiw+JdJzMNpIcVg8Gs3MM3yQrtB6eb
z2+7ierTE9A38TijCh4bXxi4drjcVF8ZYW/JmgN8IdkalGRLcVYauU3B9ttti82VN+dSZi/wSeBP
NgfNjSr3OVcAzJXmf37SWcnY8OZTFbPg4J/bOrGXoDvFpkoCHeekkxzi627pCwb218g9fewG2Fpq
EzVa0QZaSM5SsGGAEmoDwh/bbDeaKlR65hJw5fxjgWnSWEZp+D12+YzSPNcgls0GP9e8h+brt05u
o/chXEWXTrNOjLUzQu/6xTyuH3CMdRRujqIt1L/i5Wm1siu5qDxO87Zd+05BDaQhNMI1gR0M0+0X
sY4+DOPMsW/d6scAtoxQT/VvNPHyWV0BV8s2TdxNX39S0PKA3CdYXo1s3azY5yrbTf/XPszb1bqH
42HgDd9id8dv1LD7mF4RqPQcgqrSEADyG5jBQ0L/CoM30R9dXvIZ794HTSihTO27ICdTIycLiwRd
WEUfQDZiNuTYE4B5oZvGQ8Sk1hHIIQBz/hLI3TV9yENNesHN70eZu7cvRNow1OLbgX0XI6RhIQIv
i+er25iC90R4rWa40SGP0EwNvPLyLlYXkmToaRA+zAuGsZHWSesYL+QOnjUUOlbcHrKP0/8hU0Y3
uQZd1qw9BDZjHXAyzoMnOE6ITv5Gm7mGgVnkajwOB0IrcO/B0+ULLgx3NI+pM9PWGvevdC3CQXX9
t1luOC1ujjgahb1mP1QkOWQiyD5xs83FYZrg3KgTCrOyfX1/o7CcuhfmBnfLKPVo0SNJnHE5HeTs
XY0iNW2Q6WCpYgqVbHnWuLCBxWFo2fZveip/lv7EygJqiXXMmPAyvPwGbrFdwG1xyDQx2KgABG59
N71KuQu9rJwgZdjQSUQIvwvu4Q+t9Hwoi3GtMHCTNSrwF4WJQf7DWJalom2euTeGHEBZ+rxmM/MQ
GhRzUEiQegQNfmknrUB1FTS0IQIDMiNzfnwFt+sTrDGK+2BPiKyTIVxog86C+eKgMo+kA21B2kzJ
MQYWFtfZYsgr4OPK6HZne0LukKk6Sx6+Ko+bZ72pNroLnsUi9/8A7I1a1VamUYLl9V5pXYXF1IN7
UmUCgeP8T8R/XT/m/hDqxUbmdq0O3o76gdu1FhfUnvFdUqbEn+Jxk0hKuznOIzq5XYsgqn2tSPWO
P7Td5sL9vZ2Fm4ldm7CcMc3HKb2fnb2CCQF7/kcbY5J2D7zs2oYXJuqUcVU9kSOKMB2Zu+IdwN3J
mn2TbZnb9ne39aJ9kT+e7nuGml/qjHleH3uODdDI/q88KyRL0unNh8TMZI4SJOGC237fqi3mQZXv
jLx6MknIdUHs1eFM3vBE5Fn6VuXGMNY5mVEMsh4fr+o6h+/4zqdjAJYQ6YeUpKJZCgbPwN1GEYE5
bf7Hj9NrEy0aP87ydkUF0VgCE1W4UxGuR5vpn/nbHmzFAlCkJM69oRN1C+Cm18fY7Pig8YhYmgnM
PfNqEICQ329kXhXH8BobrIZkPcTJLdxEhjyZGohT0ukEe6k4A7Po4tUMUI9s1JnqXLT3fvvIlAZK
zS+YRLMK2ICeFUk94lu79QjS4s9HXRKpPrbh9eW38QNi+BRWT7Wuad+s+caFOXbwQwk/lYrjZtRK
rB0FNKJJofRzcyGMekaFb2PF9gBB4Gf5rbVea9kagF3RbuXg++HoucSbt1PVeZCio9p5Kel4yCx+
xZM3H3eyPowCLxGTrxnKF/9RbytPAwf6Br6tKNyS4UzciVY1ONqkefVmuXxrHsm+gBdNwGtCIiDe
K8E7YC+32RxD2qBwlxL0kYSJgi0hp6AQgwiSIC4L175XFkduLqnd6jxnoQuUNwpGg+G1ceN6E9dB
hy9DFc6C1O3tdax8+892K6KQnz58HUHDY0VXOq35AkCGEVnKfSPlo85PE0XWHb47T+fv3ateU3LA
260rW2gmeOjiFraHq981V39tQnGnI5PYir1E08+LjZ0WjJb5Kfrmv9vflbEluY4K9JshVnqtdsoJ
m/viKRDeicP1AQdzskVlyK9rx4fAC0mVgXdgIk3fWZI0EfN/oNToQp3CmomeuBAuuM9ExpvOgSle
c5/LIRVI9fJNt4aNcce/JAc+ubpeKb96HToxkaKk84ilF21AwbGeL3pkincYHdulG0X/ae0+A+lF
1qaF/XgkZjbjkZoGYRvTBuWnFKqFpvPKnu0DPfSsGzL3WpUz71PW35zRpRmPDgl0fO2ttS8EUv12
Iow48si/ykTd6EUYhhr13AxeflAcoWAhRyEeo1b/fD3RRtHR4TieTb3DsxBZSUNFyqE0byzBXfex
ufhVtE3xDh09wuldCJ6kWI3kvSjHCY2+9JCtcEC+UnUddeWmDN2cEACDByMLeoCRiwHcWJrlrLuv
1NPXNyISpjckrOko+kP9cdeOfdwE2h8+nFRO5G8zpOlpqDl2t/wUWPb+yokZUaC93bG7WzVLlNs1
WpbuMEcz4zTgrPwxlxt3KiaWI1P/TSAM+kFbNVAVsv6HO6K26FFZBcgu3gWlCTCyUkq6iiFfH1vN
RTA/0WVr8Kf+7ZCVAPyKKEJdmM6md3hbdMiO4ZNJHfp5gxKiYGFgpha+eE3FY0CSr63yuAcRmTO2
ARk2HCsf1txV5y/K1YuuRvNerSzDX4VVxlWJ3C56mV/Gbei45Ov5d8sYNL32EF9mnAesXn7NarPO
sc1HjT+jLjuesskoN+AvywMAdOOUY+k/eckjvvgQ+sCZVBISJkcYSPC093R1yfRw0xSG69a5j82T
1Be6A9w1cNC4qpePSo6j5+RKX3Oz91ahPSYWg/9Pmy8Z7gG104OHuraYsWVZ+Nhu74ttU3gmfI66
Boqrnb2N81d1uUhbq960qXb3/JFVY702GMZxfCkWhDZYMIkRnMc3f/2/lvhCv7FwBZ+3N0Hc0nNq
YUo2t7Lnfg07KbMHHCMXUc4/uk0WiXWwhfMWcAcWexzfe0yMlaak+j6prUZ5MaWkJAyVRRhsNGZ3
3nG0STEzVnzY1FAphoJeAtw3bQ3WLePUHD6g8DA7bf0Q4ktvUGLauBoZDeH/q7sofuRfc5OiEd2v
vCNG/UsZI7JOrA4TfzoN5SgCsLoqKpaSLc1yA5mzAW8Xao5VkMkz/rWE2yC4ltLw6Ha+/HlaGwto
vdlWeXXZ2myS2PeNJsjnraiTKNPPTb+9affbao6d4o18g4q1v6QsHRuAHbGH89/3a79wvNo05Bdp
OyTF7cu3661YJCK6R5Ln5+3puiCUWWV8+7EZpztRLSPlMpcrK9YGefVelF6imC73/5sYMku8oOMF
uyyE8c0MwjnXKfd/wRTbeUTLZhU7Pxgv7WTIYhu7n5H1ue5VG1kiVYJsgAKllEwkkatd0epEXCkl
h/N6LLweHVDTmnc6c8i19a6iM3UybEbnDDm/p1Pwq1Hu4+huyNGWDTD85ld4vwemqAlofHCnaQvF
ezR9p/aU2xqPAI50bblX4xJstzb1QVyRAIt4Hab5oy6JB3McX2obESD/QuWvU3qkNwD//7t2z0VA
BtYuc1qekWNX7/2taDVhdP8OEr/PG2Rg+ExTti2GetwXjhTsOadfNZiXL2I/m8PBu2/4DVjkqqTX
XZAT6fz5DvexjJtiLqc4ONqcxw72AAbuU1++OvGmRYQnQ3rn8H1QYZPsUPY/+1IjbxeoW4K+v+fg
Zvqz+++YVcgq//YnXg2NG71jIPzTmhq2naEcMs4osZDxO488ayZDll7cHyQ5LOLcVjTcaspO0Df9
z0ZdS4WXXwm/N6hMZIB0gmoCePyJKqsREPebKbTAw6bDj9ZpDIOl0MJJly4HTa9NrI9h0g5+JydD
UyfSvuquXGwiXGXvWqKYdhgSR+CY/AeoxwnfnS5QXRcov3VPa7lsvy7c6W1Zsvcm6U8WwzP6GUxC
e5/rvwnrEFZB6K8MpePA5WA79OjbgUCwteRaHIL1fQj7IRuLXwfp2JFyuYAQJzd1TOqBhoXHbVYB
0jfDlCxwW5JODLdEUaiKL4l79okONz7iIGml31lgWNV2avV+dHwxwLG3wbzQOyTDYfThIPFcOq9b
DFkSw9P0YjTHkKPLjYzzPjhTizRLzTSoIyORtwpt0UUVOPyfoZkKDZTe2kZk6r0CWMvVIsch9vOL
PZKTORHb/Tr9i2whKYn2dYTAw9xnLy7ZImH2JSNAtQDkzNuCNaq6oBnBGa7VWvXItrvuupJ1wiPM
H4+IWmUrAMG96Wfz1LZXGRdSxaibGeMtXW7dGKBUyaID5XvKq/50QjPzNdfuYvavw4caTk2QBDv6
Hkg81f6Hdb/TJWc0NZsnK5EDVKgEslCEKtdjnh+JzNFpj/elrL5TtS0xS16b8oNFM6pKAbwd6fu9
ORL8UqCUg6mCCotKmj2VrbI0BG9esBqQ5+oMuUQd8i/fcoAblkz9tptt3ZRvEiQZzcIfUOvcuN3m
T8/SzQ6Vb5lAhwX85I1PIA1aXCO5hRlDdsDL5moVusafIrSvRIc8IF1V4hioFYw4kXPYvqSc1a/d
I7r4+qkSxczn21YuxdUX776KR2bjVQ/C0EthfIIyBLQGBWLMcSrX1WL2iJSU9eN5N0p5C0ZedQmS
4PpIIootBThUPqXOqnIff602I52P/TI4dqgPRfgdbNbo30K4DTfXpSHDNVUpYrb5nPl6zND7y4Tg
Y35TBst+7+6OVwHa65b0zuPxr32rOCJmWg5RDT4Xj4fHeUg7pGb6mnV3Ny8Uym+g73IGhHMnqA0D
qihoQxa75sy5n/bcmJcYhTjucEn9RvLHR8yfqBuqZSpztfkGVmYwOE5+5Nyul3GgpuSxzic9/gww
DaEIz4G29fee2BHP0K0i4mlJ3EGmeVUSGPQWloZ4qWdITo5P9VQJQkMaPqCDX5hY4Dj+D+ugMgja
bG1lPUjrkRwfvYFMgdADiRg282y92e86g21XSLLS1RoDNpVKQq5M4bt9Ow8gYQ+VVW8WBd9HVlKP
FNgwdtpTKh10De+eixVhcfKo8jMrmABC9kTM3ajm7bi3ROOSCT+XUnGktTLBjvPPRY5MZuCyvD+p
F4lrYqN0Akf06IUU14ie6yuUta3t+c8vyep413a20cDzVPrQup6jziKDLOVzdrWsGcdrmK8CIMUB
gY19zfzS5jHYG6RePjRWhhQhDmAMKRNZ9T40ZvvIV0Vlcx01BOajEToOCdf0/kVRiBSJX89UWPPi
/zA59QLQW8WaN+MC7oPLtg/dFgtd8W8orj2zscX8Jt43m2Lgz/X7/ru7S7cVf0pu+Y5niaDglQeM
0riMLfSE3rWELqJeVBrTWkTZgw7lgTBSOTM9ClqBl2SNTfJ3uVYZsUmSU7Q3x7NeJvksJp31uwCV
t5HTFMQTEm3zVekmgrV/EDlVOIi8KRO5xeSBR4slbdcUmEvoZlvb2P0EH568BQFywZIs1hA2D+j3
yh2sSKKqnpep2tzAIbzMDOifRksxKzUhu4GFZQRXNYuq5qpulcrBSn/KQNL7cXDqatJtPb6JYd4T
t/skdAWchYHqIC3/bt3cYcU96VMlBcdqa9seiczpsW1WLhz+vu4o/QA6s8d+4rBHVNNNcBfhuRsv
QMka+OfLwR7mX3IY+rNsHNJB8Zh083n0HDb1YrOE1y32RKJTu/CjzqmqBHVW0T/fcHotsHlYfqf4
8nZeVCSJMCztC7g2kfTW8d1+hEi4ppt+culnIh+6pLpj8vozEa1PQZu0jWC4XdfZRuQrmHf9fmhN
HSQ93xwH9Uj8quLCbTcZ+u1h4ihxWFVjrbj1+gVHNn3ZQPXJw+L/hE7VpJdKhwtKa+9y5lI0UPOd
zVgPPQZhi3aXkVkKjzGbPdwzYCydRvR1yUbhSLQIYfYy6Sp6KeesZognaY3dngufvUStuBN5IY73
LSpuEqvmCqTCo5Mg94F2xL/UUpNFXC0EDduWUHXfqHHRkOvB6KVv3Ok88J143TE5QXRWjODG3azf
lM+Jr80V3gtgOmPLlJkGioQts6JTzwN4cx3VHpCdT8kWSrrg0IYuH0pgiX/3cPIZFgULasu0IS5u
kcL4Xi+ZatBw8hXCcaRpLSW4/WLZUJZHhPgOW8cRa2IblIkGuGxsmPX/wKdhFeM0vVmyX5z1Zcxc
gQTgRl55okGEYNVtgi+pCgt9a3sWY5lVgoqhYhw3ugAyma/Qdss2DG3bO92pLNVoIKXfmddDw9cq
Px8Yc3b9jR0XnFDStlxnjTKK8mue2kcE4/oRTPYRR7hchy4trcU+Ad4sU9NetuEI4cHLlKfBKlSY
fM/88FUKit8vR3a6X8CHBfkS/OP8szROVX/soWckZ01qx+uIvaiqdK8yHWSLxGsyIXnF84He38BN
N+AiTX5a6v+zDBUCuWiA35un9AgJRuKBqAX1lo7MI//8g7ec9FCeIwQSlkZ93u7E4t/CcxLpLiX1
K4ymLzAk7OUf33wz2Tw4fmQ/VkJ/wSulf2fWLz/fT2+OYVQmfeuNrkoh+5brA6TbFmg5IAML2W4Z
evMMtM3Loz3UawhwKhwhVwK5uMah1a2aVmZzRz97GtbVCd+q92ILAfUmo4Ba8lGSatiQlecEfQ7j
5cA0cHDftN0TPX7KmpIQLbcORRYkL4gHtIVUNNdV0k/0koQ6Amd2+Dt8fVE5bmPo7Qx+xqkbqU3/
1F10WOc9feT+Av2ptYI+gFobZTtYtjPpoqM9Gss1sWSAou4S5skKlN1lrlaSq/fNl5VMqOFTsvjy
4MG+KlpH7eszK9s3JSUlrvQMWKr1/bcwyYTvI0aOblMpkpArK4dzBgmRL/rNBZaTNwXn0b4nzebh
umhQZyRK4a9NJts5rdr6s/ya0A/soeqVoCxpPk387Px0s2YroN2A5HMZzm7mZdimkbVLm70nHVlv
y887OVKGs9okxkcYY/OE0+p/JsEkvBBu5B/QxCMR6IAhLwdWJkETYG0omMCSXOHzUpGJ2rad/5Ry
EWw7iaZ+pujMNW1AnrOdNurKmoq3cHoIDoWBEiQ1E3WG1FBlEbGhEreMUnnhwoIF6yWxkGCH7yIP
dh9W8u6L/rEYyXoF4Ls4RAhFX26AmkAxzrEpuhfsS4fFqxcst+ga6it8eGN8R/fvUkY5VzxuBFB0
+2M7JbX7E2RRptvi45wXZW1/+p7q3yxYG1cvcPUMFWShvuCgwbDIb3IqpQXleSA4MoZHLAG2kRQi
0GOahuteHaG2CRQ0GGFp8Kq3GqQhnD6HoOiJBMr/NWgF7k/vRFInm6steN4wisWfJuifOvhyktC6
sy7KqkvNTL8XzvtG7DLQdXRx9CZVouK4zms5HBqScYlrty1mMN/VrDCZTNmOnwNzUAxvWEbJZi6S
Aip29k2lyrPlP5tpdr8WudXtI5xZjMrns9jysRelsh/Gpzq9sAz1c1zJdogCV0Tuh/h1hTKpK0/N
6aP8twc+I4I5wl0bWMWkbYZEE1gy9JJ1A+t0Zb5fBILzFMEkW5cD7eqfD1El4nV7QNQW3WvRRWkl
tG7qDia/QmW40jan87FZKWQyesk0W7BmhPFz4HBeogsFANxhA5kg9mj3+yQ+52zb2Bh4sZSzTmsM
YQpH2ceJ85MBznVaGhD4fPBrwO3B76nhonXqsK0X2yIMOZGo9EFvGyuwSgZB/nL6F1Bx78qFBPm2
ZOOkFWNMuEG1Iedt6bcMV6QaQDYqLrN9hbF4zgF8vFiCuxj3frG+dOGOMQn6Q3qYgdSvDLojgFIt
UcMOWdFzmbT+b59dRBVKsTFhS70CAjgxK+V2mNol2uTtpo33ouZxmiiGeqGXfmV+S2C1u3+/m2Qx
m72avxJ3xqbPOyyi4O42AVvfHk8ph0CQtkct7xRVvqWrtoIK02RdSSe7xCbXgPYQlxq84MGu43qW
mtTAdStZB0aAOPBkRNAvOXE7xJ1YkNorQaoN6Sm9dxMa4afShaWorUp2cGhSkrj6spc0UeZ+Vidn
1rFnTXumgQh0bH67DSOGmkZQniDbJgeRtCl9DSr2M9Luuj97bkYwk5V+qlH3rYvSbm7uWO7XLwHi
hvg1zhmiCoS92JfmREAQutw/BdUo2BPK/uWKh83Nt+34TvbbWh8WWTqiPqVduucKF1UQHo6njKep
BTzTLDhSl3OA9FJksVKGneMMF0aiA4bIlouBSWQnhIgE+YONU/ljXbnk/zv1FS5d+tjunQXGrL2c
85MuKWPBF9zkOjF1HkWRZmfdz3N9UlbAEfq/ceisoX1SG8g92HFlmKbL3D7KK1EIqi3n55oDKJl6
kOdvyotUqTmEpqKe30KIca6GwGqDVTYGykGgtxgtSf/grZygIDHDinXh3v1VPa80Hsj63fb4GC1Y
hzN3DF4qZmkJudrxCgyHHuRGkhWR2NnaETnaRR3m98dhEsDYbFwfOYEYnHJ1fQREReTc1d9Lpq33
A9ECpW+/C8aIYcO6kaE4JNBX90vcl6wO5gzko7BsYgYRth6pPxBGMdaZzxpS7fjkNPhw+2jvQ+4N
788KD8lXZS5/ObnSrOXw7tBdfELup9OpxmKTdAwz4ePqfax5FWKy5Ew1bQAQ/aXgHaAqaH6GspEQ
6zVfWh7RRPD43Acjxkyh+GFGhHBR44wRL2XVjdidxjRHzT4vjjp963wWy3aPc5lK2043KQBOHq3z
dCbz8tvt9YQF33h58hRpL3ECJt99nlm5RXoGy5HKWtpHCI7HAbvi4Z2yQCZIfhAcB1s15oOGD/aF
g6FA5uqR+T9maLKE0Cm4EvuH7WUYHC5QCdTEMkQAW/YaBQ7PD72xS7uC9MKmcpTDivlq8VmhWH1y
q7nLNPPMVNYCINhmr6J8PCAdsaQkBJiuARcHavJlKPXQgV46BsG6I9cQQTFg/JUP/vtZgDPge0tr
4SNFPwmsYxBGLJuqsd35UMFrC+Z0N73zFIawTUJiLT69Fb39ezvS/u0yCZX1OOLQBt7VSFzsTxvS
zdeJLIdatHr8xxG4r4vJLPbukWTvz8E00CXzwe+nu1skNJr33yagu6ltHjDPDjEXB3MMXLf7LbNx
FJdsE2c/ilPtCcmGvyzj0FcW0yQcTij8z8UX7YtQdBl3OnCgSqWfUTnqhUKVlUNzE1KItZerlK18
nr/7kFd7uWJjO8YDhHU+ejQYSjytAqqMRLdTGC4XG/YunnDtKCJehB/s0SjBWMjNWKJMRjaNbCxz
NY9HDCp97Kc1pcWJQG2nALTALS5KgJ69DX9b29W3ahMClvZhT8iLPctLBQVp2TWxHGHMxyvg9Pjq
yTMJux5NPZEnY0Bq8GZ1F1PNrZ+lDjCvh0FOoPCIS6SzZd5699vnEUBNTmr/pvmYvZ9rEz7c5+LD
dpqLswiclkpTL3j79kS5moF+HuZvs7x6mxGN+igHJlFDcpf/Vn8xhR2bzwkuMkiqLmZdTE3/jbA6
b5f/kXXEqN6dpS6Q9flHE1JZiAZyv/nN2XZWybCnU3EHSaDuRNe/+s189lEEvMiD9/+EltTcRwPX
MHQ1x4fGCCGlUIYTseKwifJ0ztmj7EryyLjmdwM4Uj4jvy8GOhJ6okeDKz2L8LBEKSzojZMrr9Eu
m/TnJC5HbOXutXq7UfiwpCNeiKjbZYMpBoodPG23KAb25ezel0O058Qwe1aYvAElRo891rwcSKpc
XgvSD8QYWWuvepVrzz3d0JP733J1HTKUgWBrUpNjWa0wp6i2gZZdd5kVM51tFLC+CcJMfJ+SiYfD
RvZWO01tEGlakcLxVi1F9Xa5Lm3t8Ebo4qBGNPDZNcLFjNxpLfzHtdDTNgXHwqcO+vXKTYrB1WXe
SKaGbSh8c6ZjiopbbCnnFbbdsg59jBWc7Mn/4K6URaooVuyBMw5rxfFLlWspTOwtyqiH0LmT+sDY
DnUJ8oBD4UaGbJa00SkR6QPAQAmtdVQx/6Bxk25TpCCEZUYA4kFaHXqhZDxRGACH8WZgh9vq4CRx
b9v2GTFJXG9y5zJtkDNpgRHgAg3KgGociw6ffuMt1NuSK/7TzlN6Q+j3ydd12D7DSWOFt9FlsLIN
54This3Xz5LYhtAcX24hekM2vfi5QrPo6sNuspaPcpe6asiH8Arp5PjX3q9BcxkDpvjBMGHoI9Mc
r9HTyVvcQxLGyScH8mJuADN6ikWmBgFAuGoWR7F3CZHE3CLLLlKQ7h02mXFHckAFRS7i1fHEhhQD
6AZNeYgYRZk7jVu3A9B75CwxoXAOQ/e6AcPTBajcaa+FhdbZ0+siHA+eMcui8+grYqJ/aB7nZ2yd
+Nb9dSSdwn4Oqjm/3LQwVQ9YvjxqT8dc/NFw5ktaoYAJQ17yleIKJXoMYNVraPUwPb8biMAqDKnp
3mtFYPH5l9AZpzATX9fVbUxOVxP7bw34W+S32T4cUyLpvs5tb51tAVlwGi5ulWfgoN3tOCtwIsFi
D0Vu6gnWYVucC09Bpv9ccbWADdo5QD5BkevOZ03taKjtbDY/uEZclRxx/oF8P/bXOYZYRxc/onMP
wNVXw3TBL78y1z4IhVRKQPgfkElTrn+xcX4XmxEdp99WJT8PBIQbqJEXxu56dRY8AFWjS0kDdcFW
bzMlVfWiV1M1M5geiriyFpy2+stG7ssV4tc+GqW+62U5MbEj8uBnJ8Hm8ZakFuQv0duz73uQRT44
4nZJPqkbCF1sbX4ZmCSZ8Y7aWxJoBXR6/xWHjxvsyvuAZ3JH08J/lOSZZwmc8iBtkwh+IqtlAuS/
0x4tmubs0d/HMBUNavIr1KcnI3PZh5Eu932BH2X2JYDV7fby58r6SYvb4CY3Yaf212JHDD29GJAg
hwmqCmpoAj9j7mm12rICZRcBpGAGD/n6BTY/ElKQlYJHOasdZCls3mKK6fj6H6LljfoUAq7FjLZW
U/FJLLHUJDZC9hBiVCBScB7OSorQTwzYXDo6Aj9mQKIStf1IwVs71Sc6e3NfvcwUdZZbspqtqHLV
onyohZz6Qbsn3FBicOjUdZbpS0+9d3Jcxjl8NqMC7nlPitLJbIBc+ODbEYwWUsorY0azU0mCshAw
iC7xtqZ0ErCvO7QwZgSaFDjkIWntLh8dlCIvbLQZfJE9DZjYbsfW18+sXVWYBreeirx7IARVH8EX
l1lYt88w1fgOUThak6M1tqUEiVK0WmHQPMabVHHWCqhTinSKdYzwkmJZWAYncPxTT4SWTUYnM4QZ
+iRWT7nsr6gy/KuzbUtB3yMA1Px+j1f2JvQKWlPjhkJXupZysxDexn/P4Mb89Ksc3DkijiNHVvQf
cVjBAhDfju74ALHzMYHBCQIzLxKYGJLuuU1EGr0QLj66reW3N3ruwuUtvpo9yjx8fcS78DJarpc4
Busr/WjTL42MqxhfoFx8qYE3nT3c8HUq2IZ6WFBxG8XtD8/r1CXpAWor/VvuabaPGj1RQDTYwiZ+
qVONI2CxF1Ym1Yt4tOkf8ZJSUtsFTHT5plCrSxHMAvnTh/tDabouqrMNxa59IBV3ttOpZq03U4BU
HlUNJ8G7AEg0iG2SzauWkTuG6HG4qtyrvvVlBvkEXXm27tLu2AyacyoZFAeSofhtyIHAQA8Smd8F
eKp/SwhYbqy7GZ/bIDh4GNMptxAII/7+ixrMJ9oJFi9n0zHBZjSJdxZpQRruFogPJY6RCw81vttN
khJEGFAFYdGAjUrp9NiMgka6PwPJJ2JlbH59xe+ghufGtbTAj52Zzq5cgEUaesmJFrBDbhBygydv
HKWs1mNvD6yzHloYYtHgH2Nmty0OaLe96S8YAg2flxZCbZUTcsQvy+Xx2FSCyqFlylWmZT9nLGIB
QP3PIm3o6PvLbOwQ6sTaNvjOrlLEk3+4S1wd9+yNG8xxet/7zG7bAolY0hhoGCx3HdqSB3Ni5Nr9
92aXlMTQKaC0NNqWgrmCyVBU2ueeDmEQwenyaeUb4tYus2TGBr2CHpmSRyrOd7TvTJzmvbeZ3Wa/
ICwy3VV/ePyikWWq+NNLYOKHYL39gW0epWXRaY0xYByg/anMP8OFIsVjpxTMI8hXm3G94k0hq8+5
Gm4QD8B5b0iN1J2e6t8tLZKTnfraTAKgPrqJJUjvgZ4ZHEJWrpN0qZTiJvw88OGxrVo7Mcg8jz8Y
p3v4HYICbO8FmbEdQUEiBRewnoqd2LHz9mPOZlBKPxD7lFqfszBxGbyMWTwIoWhSnXfStklyKlcR
w8E7ZPFVLslBLWYjGKCdrvYtRE20TBsX7ImPwtcQbi77LgrouaSzILtGHz6pjQrbGW0M0Ls2ICzK
Dm9GuZPT/RopMkVegRop7q+6xc2F6/f1EA1TtnKBZuPvqnwtQfNhx4jfKFaf1Pepw2Nac9fROiuN
oIKoQpnfiWylcmIfIURXLOJ6jB1rBUlGlJvhU7hVEb/+a7r+39B+4wl9GdDHQWsMhVUpF1L9MYk8
CRnNAPNQjakJPntUJAbJpRil0Z4miScpm43Yv7RNPw+Um8zhu1rkoMgXaqSaxJBi4w6Z0S9ejts7
NQgF5tcGKdJpuvu6rdYv04wy+QndrHhRiKL7GPGrRyDZ2ns3qWLRsvmkQC8wZOGZzBHQKhut+VwH
E4ezDj5Pl64EZz3WUtdafEt7OW4iemMEFUrb875mIlP/tBjH8rEp4uXnKQVdqtUgkeS8bGh89V9u
Pc45uHiOZta+vGXTRunQ4NFtVG87H8huZqpdq+enzzaPEZR2jClnuP0CIDvMlS4ehYOGvBA79VlA
XKxF5N23McRGzyCd7mhnBqxCUi6O7faILNFTqgMkvFh6vKQivNOxXeYcOEd56iLorerdQ0nXbNwg
DAbMWyfFw2pHO3sakTHAkiHlox2R+V3Dego/UPd8riDLJXj15V1QiKGD9s8j/elfJXAGuOJ8NqI8
p64HHkwjMJ0ySo6oSi/aX0REsBcQAF05MnDFRJp07SLh48MjYIXqJ/HhEKX3yZJYp9RF/2yFplpe
mvOKbn6S223oW5CqpoZmPUO5contC7FE3QwbJXq5TX9mWsbYQvYNFdMr02tiu4/HrIi8BbWWRtkk
AgoWgNJ/euw/TxUGx1VJlAXPdEI99id2qXONkutHY053FvClKuRPDQ3sC+7XjK0miUzx56TskOg5
Nn8gt/vj6MeC67AfWGnXTynqHvsHtMqqPbJuq59FPy0lS9l37c3SZCr+OH59FtNLNhKOebrLI20s
F1lyO1CYa5mj4lutv3/6sYkT4teZKKvpdFixhglKBGgg/GjXkpeem65wPQ6xYC9xTfCr4SqfodB7
2D1iZnlfmO+Ecuhi6pOYy8MOkwRUqVW9aDFczusKZPAw2TwEsR+WkzEcx39kM2/OP3IN1zFTnFRl
rCUq/3d4VxzpX0eFmFMleHEbA3j74HucI2bYbVCBI4kIACMZtWvsaW9J3nbxw0iQQBgHfVkux7HR
JgBrF6VxSD+7tBHCiAnNGtpO0bnvVnLWuP4wW5oHihHlZL/Go1KZEwWI2OcgVxhnP7GqGhpfAAlW
npx2lde3T1ua1IeyA+An3ShlDAQ8o0UGC5wIVYAsxBQOOsdYI+WOt7g0UoOIGCoK5Z+3XR2mLrN3
iwlJ7QcVm4ElM9Gdh0suIaWHKxmSV4FNH0PsVn4q0qZVWRy3xYylmrPH2txYFMReOJ/ZNzTxpc6r
HXQ/0V0b2WWv5Oj/FL1QJ3cTA7vtWXil2LtVJRzljR5b8dv0Qyl8HFkeqYS6c+uR+533UJiiZyuL
lGXLi/Bp6a6WGJEujgiov/+9962TKuknViaNy7/RwJj6T4xqtOjGJD3L5i6iKR5KPQpF6b2SGalb
fuBUgkCjB+DR42A/PQWToyodUPDFab0Nk5MTyaQy397b6Xv8Eo5Q+b0IhCWQaEzC2/zwy7x8UsQ6
AqnwXCOYUyoF2T4AIkupVnnGoz4rF+i7Ma/6XB5XWmVDBIRPGas1/L+kKmN46cRr408pMGNntqMs
GObLYzWA5siuWPnr+4XYE5EO6l4AYA6rNTHAoASGiFN2KE7ZkFcfREKsYBMF5mpmVlruKt45VOUS
F5SenjDk1DM68rmPqkAS6ubuq5pOfMall7CUovPyuklmoAgzcBxlqjkHNyJsutA5S3V8ucagsDM9
iY2TW2/eQAlxxeumj1hfnE+Vp7u9XitxByhikIVfgJy3KE7W2GXoKXSIty2uuKSAmSGQtcLbGroy
3o3OEUu6anHkiTQsV5EsvyohyQFY9bw4lQiL4YnH+AV76cZYM4QYmoxyhhlz/XF75QPndgJzAZ2+
6UgqBByiLeNHLOpUM2QlRVtPY4UeGL1V5qgvEgts5RysaOOIcp1PWIMk8cwB1TW2gzsurTRVcU1C
5TuoOJMqnra/Nwv3qOyNb3xVR8T1TKm/g80Smxyw7YC8+GT35TyV3jD2u23G3xt7iMJnjwVVVOZC
eKqy/5hfqejtBT40zCBgqtjMfhiHfGK8uuNcypToMRZYU0j1LcM/E2YVQoOjlcfrg0yAGmfAzlmN
DLLfKsQHzx4mczJvCRw0BiEze7AJVZLDUo5hMJcgsA4garqhrtHC6CuNjSG5YSeLDbgUVO8Yum//
06vJRFtb/kGFllwE+nU9+QPrDn2QFIl05EHf+BxqNIl1cgNx+nEn8BQTmEk0T0MC8b3j0tdS0GuZ
1Piop/NZAZfmy+5VzmHjWjoPfaWR8HW7RSSS7NwMiGlaruG1kvtDnOlPdOhX6h6wZ33aZKqq0mcm
vjO+xmXj9ekT/HUzXWjJ9H9D9uO8zqU5iRXJLWJWNHFTBWm2+EfKDHMt/wMhnZghgZKjQnSOU+Bs
olymApHxk6dZuEIyeD9MCX5oaPvIA+7GiC4m38HmiDZRokDy9Z+t4XZql5TU0jxVHR3VqsrOjdsc
xPYDMyN7I8YgHYw1bF6pp7knF1LR4e6koUy9yeK9AWm9NqNui0LauHxx0/wVh+x+px/Vz4OXWQs+
0dW+HyWsndQ8zNudOLIHq1u593NCO41BhPVm4jWI36feyUqqj5626E74NHcMYmctN/cC2yq3hcRS
02yt0Rq1ik4lUgYDK+JvM0LdWmZgeI+azhTcUO7ginB/Ogy7Cls3LJ3CHZgD06EqjJoZjMJMhWW4
o0t0zjc4pW5aXJm+/4YPCIIQgqezEqjDmByLBzRJoMktTTlPlexBPfDGW3wL8Sdj5hDHtSvLnl2n
rfZOx3R2eiTqiitHlROgqNy5MJcsw4/v+EONld0D8pjLXvrpuwyszEfMpWBQCtPaH5ipAVQGAdML
rehsqv1IhQB3dtyqXo9U6ro75I4z/0SCX3Zy/nywCFWRrD7mKypYrI55OV5rywsI93/YXVm0U47h
GQpVxocRLRtor25nacaIY9xZEdHn1m23UVDlIJlQvzKL1J0gVhusfcSBTCM4NrJtqjonbs61GTov
9nEWc+lD074lNTXzq5d/u0lUq5GzhaMWcn12OlIQbTE6agEqhrVR7IurbazcWskW3dwSoPjqC72q
qVQW8Tp+pcNyohQGQMv9a7Iex8kN/piNumAVUp9OWev4zPXtPDez26yCTpGXXSS01rnSI3aSqIVT
xVm/g6Lsk2rA7DQNWphMNBOAWFIlwPb4mBtCzUPytCMtXT2/0r01Uu8IKmaMpgcuD4zMjw5liDaj
lCdJJEmdqI0+x9/IwTgxoy1Zp4YgEYFIKd807pf7fQo6atUHdeGra5q4rCDPIA7wEcM+xG0qLKsZ
f4BXxIX1G4jvxGChkblTDmdsGysE3EGXDemkG4XdOnEEqxv6y2v9w9IFAdk3Peydfva1aR0AMD7v
MEXW1TXjz1CWl6dgCtd1C37iv9lQy4u7T9UHSkmKXq26xx1b6Pz46yJXstkWqFmLM+IvMzCsKSeO
sO+JlCwk26vxI3FR8Kpl2ffJmL80tF2fDao4SqDYpSUhdtK2jt0HbiKZlX8aBOgBTzU/uJJtUO04
rQrrChzBbmoYkINPOqs6VcE281z0Ui6fgMnIdkI37crlTKltR6UuEkBxYVLoNGVDf0EX3kBpstUC
GdcAGN5uWyUfO/vyyQobGKYCuZ2BoFoS72juCXMZHyRaV7Ke9GTJqTa7R1JGjKQpkzql44lIdng3
rCzMB4dPOCo+lVjkLhez0xvahCAQIi6mIbFtSbTXPz5W+X0HqTldI+V/U1tLao1mWMtFqgoAdE0b
6eMUP4gMM+BX78q2RdXvH6k4W+cu89TZ3i++bcvOqKAcC5ueR17fokPCBdtlMiWZVORIyjc81UBl
ECNJ2O17MsZ6ENAc0mM3I9FKKbfj2qPhU9GsBgpDxP2dYZfRaaPlUnRlkSZEfCEDIJIcsmabq78k
oU7ho4v1NkAMdekiMhIFaOPpbWRh+GT42lUeS6dXg3Vy7pMXCEkU1fYdwicv+BHrZtWuN4X8ITFT
FA1pT1j9pgYKHfKeBeDeqdco+iU6eB4YlWrrNBRpERqcuk3531xmcRz2MXrR60Aj8QY87zX5KQX/
xwM7Dio1x6x1st7cOnyYRYtVoh0UFgvw1D1Js96KwIC1uJ6uRPMRiZhg0i5bl4TG/9J1EwZ7cT2Z
TT85Ea0mZRlSt+iCF1ernDOnb0b5//U+mIpTcuOqNoPveyqwJL9Q6CLuMa0Bab0Vq8FkDRq1N1wc
2JPxWSf+KK/ZjNB8X2M4tD9FgE4Yffv5DEJQ26xwi35v+t/uCbrtCqAcmA83uYVHEdbN0qy0VSiw
aN9bwDVKPwkxH5xWDBjpXq0RaR6iyIvMurvKBcB2RPRLLgJoGHQSmd90mmeosupPMtXT0L6Dnob8
QHhsISkmBlnA9e3Tiokoxwxbx4hx11RBAIFj0O1lcJrSa8WTV2QqduGx/zSqqmIKzYxeT4CsZvS+
7VizJVgtYaiSGgAEgvRoy9umVtzzCc8JCILVdLArcU5gJtxtJPIXRHS1r4W0HUbPoWc3IU/8aEpJ
/hEIzZsW5DnxPDuwVm/kXqvR/UdqRDZNIZ9PCXzbLzhn4/dg8oJl6kSKshau304Hz1717c7+oK8R
c2XOBXiwYfm6HvEApCmsekhY24B3HQZj1E3voiBtpYuqZKAicX/n8DDONQNQhyaJk8lHEzpqMk7l
GGf5GU//uTT+nju7w9rfdljNqY0AJCeYzMkHtQw9jf/DcRNvUbY4A0X2K24JLGieFw9wRXYWnHJ0
Su72KtZBjHsb5qMYjvXmO+Vi8pG/8861OisoKmUtgbZli1ofQ1BytE9qJnxBdXKgoLysnHKVtXRE
G5k2ZpKWcxZrIapRLVv/g1lUTKCH/TOv6ABXb6su0B+eT8udi47KcAwp3lYsDS5JgSJeiCispz6N
rMHx1jVuqV4femPDRG7WR7fUz3odbmae6uAtDfV07GpHQAQX2AB0nRjQmW+hAp9R/99E0dOGrHDO
Rj884YERZ/bX8W7C2jCQq3u//xv2B1cy2lrAMpfh54sWrt1ucbsNL1VqCTjyV0Uw4+r+yapEac3j
27T9pnFBeZkwijuCg4YygckRtfDWZY0fyOEFaXRHOFgX9C7u+BJg+KT3e0ZWt/oB4mmej19M92LY
h8jVvT+rIEKo/JDEug6xfaDQa2TTs0DTiQj/3fjrzxL33ePLauztYDVBKuUpueWgWjdpqHp824yK
h530eHI4f67dwpQQM+p0ldBRQcZb3Dhjx48LkDcCs9BemR37tOoZHrQFO3qxwlwWQNcBwXrE+KBD
l+/YBJMWwQ8PPhocCtwnZ8d6+21cXOsygJGtOu1Z8RSmrIQLQlF1S32JNAbh9vv2yufMcIaQFRV3
lXWCr2jFoFw3rvPdAJxD98dr++rGaadHZsmbEgkMHCKQYPFG28VzaWz8Jky1jMk1Z5EcYV/lMCds
MlZ5nZfw03Z8uTl3Ow8HDAuFhsLHLeAq3/9vLO8oK6hZpvvcvl2343LUJMHGZSeddvze/xyNpjJs
Ex0m/PZu5HpeTjhggIFINR/7pW7DxCr7fyn6tQauYwjfDFdfjKiV4ysbkDnShz/8PJzsMHUM8jvg
Q/wL7vAZNVSSBo+vJ7ZuYg7c72dcOwaUpAknPdpCsFihpav2+uVLOYgR84775HwROpBvW0ZxaNb8
s1q0k/S2FcoKPzuHSUd45UglnCHh6hclGSJchBM5XzDdUNIrd0qkFnINxgXlIVGrQ+/q+aFWMO5A
DqubjJaUX0zlr6KHeozgCPjonWOzE0bN23BNEW/dxICncxIzZBzLpe4mUims9vJTJZzwI1xDii6X
XWyJIcalmQ/B6UQoYscrHG2xDkr89GUZoo2KAbeVt5b+9yypKqTPXdHPISaQbVdB2YfetKmEehxP
HDXMwkbdHJWRdJy6j0eO7rEeM3m2if4UQLhGXJN49prIBzDLIADk6nIhYTo5TMz42s9YJR6HiRs7
sq0p/FLigLOTOC1C4rBbBlk9KMqvXTa4+Eucg203UsYl+inl5qah5WSCyRzf1Gihgdh64PMl+B3Q
TGAc8hWRHzZB+mfmzG/7Ic1vOVAd6yssiqxQvd2sBXS9ZMO5JqCW5YEbffRkv31pu4/bZ14fG4eS
VU0E9zSBsZAjO9BDHf1Q9/t9ARbfPa5E0ycTaAPps7eH4M6f4p8HoNQKBNl616l9cVk4U7O8eFpG
DA9pHjfBoKsUZfcZEBF9sTi+iyux1UKqoZzXagl8NlGEh79dgQelPWIhxXZvpCsovrTQ8iRrv1fg
tPVogxEfHtVrgj24KcO4+Ha0PqBZeBP1BxaDfAIW0CSosJO7bdD386zbCuQF013QNu69SRbfe25N
FAkVhUG/2x+rPSz0grQgV1jYQwwaB1JFRXxLAShBpts+g+xU+J7VCzAvSh2YUKbH4ssQjA/oduWs
Otq7Z1fHr0+7ngBIbiet3dMda5W9X2wEtK3UvG32Kjj8F0+OQWiQI0DP13TGzVVEj4jFUOZUn9Zq
C0FB1m5kwVFqLddEeQULEBz66k0T6+gfItz8ESvdZsSBkXq9koeJKBixNZeDLl9VPLXVBq7mPQSo
UZznXzDGxc0NxrOQ/W7cvkSbjhbAMBmOIOq+0RpZHgpttyK5hYebv6oVFiTQ6RsLmGla2+9IDHnM
zyFJBl8ZgHjQ+QopGytoK8vXyK8qncr3hgZ3yaYUxsRAymoequAP0WsW1QZCKuEpBpqjE2d93XK6
L77KSGLeOiH1QyIC/VdAYU21yj4M5tEQPVDLLUVytoWshbiIrs/5CQo+IAJcNFNDsKtU/DsrK6ae
agsV9z5jXKgmLGiIUdJ45vpCYwvdVWa5VnFjJRFzicvG0Ucd44prRw7mx8iL1UuulbayM074ndXE
2ptiyKlcKXp7OiN9630W7uVV1SwF3NkhR6mDAsQfiH88c+F+/09dp/qDF7YXsNPg2BqUS+x+jxCP
DK4CFqEHUkLHT58enWKC17GGqkdGTFD59Va1PLtUX8DbQT+a5RQcLy7d67BkW5Ve4kXHDw3s71cB
gnkb41jxcHQhhLAyq8UrNBFamp+jQsI654JJCU/sWTxu7BhLnz1Dxi+7OMQGhz6HhKW0CUFVS1+z
tN83yWwXfXPB+pPboskscjaOz0Gp5xigwUL0WjcfPH7PwuFqKM99MDUH8gsODcr4syd/Rosf1DLm
ZIqdqz1QEbUGLW3ma/ThGPY+PVu6i7XGbNroB9jSEGbEsLbO44OIindgGSdJqp+iYOrjuGHpyPsd
i0H+OKeQuGw91gCt7/jIbQI4R0pnkoJLnZjejgReNH6vVFXVELAy+bcZQM+FszSR6CkMxsYiEsuK
kDOIN5dyUOvHnwdBV0aRKBsrht5rJc2wJSFVQ+bAOYjXsQCOUdqUcq2u5Zn3d4iwolYoxo1rG0+w
zvqYKWXhz1255KIfUhJzEhwWmjbCD/iO0/QKQxJDXCAanIyE5wRDDx3tSfV1N9OaHQLemk5Y5igJ
nDw/8KQu83vQrAokZbqCIKuHgjAlp3GGd2op6qoPaPO5HhQjeZsjBK3IEZgQW4+RinHPYI0gQ7NT
y9XzFS3lEsAIqRK+C4wY/xjc0hj6Kkq666C4aqhqFL5QJFbFAYppAv8AZVYC90sH8fnd2TWZIodQ
EL+3qUZzCqu24D/eN2muCo9jDswZrVw3726p+PUz7GUrMnILuqyQ2xN36hfdluzMi7IZhZhel/kd
1PmDu/EmLjIWul/ZNqll0gytmBt1T9uucwGjtr4tPCpJbw5+TfA4/BIrfvqmF2hy4r2ryAoxHdn0
xTqOjZwAsCMG/EsolAndzZ3ThJYAULesvY2L9WYgrW3eNj5k1X0Fo/5wF+jIOgoHh9p6N/9b3Mu6
+A0ijn9JlaVIfRQeyHB1PJD4BhGj60bpXOAmJfHv20SRf4ff828C2i4EBWs+2JFY/uSjOL4Hm2SU
NJegBTtgJKAH1RClIIsjOKTkrxWEdxNFw/O7mJI5VpxMfv3qFBzgN0K3c90qfJbnfz5TRsBoc4MG
y71UB+i/y8u9NTRRVOcVRY3acImdsd5FW10WYmM+QR2yFQ/GvXbAYHfYKrA6zGSb6So2Rsl5YxAm
9zl9IG3R/nThg9+QZw96CWQISFyukx1BL52TdYoyIQtFhQcYpxoUAwcmGsiU0XG9K63dfbIX2ZKl
LUbriO9mSWjoiqWvIn4Z9yjeNP2A8EwLnlYDEKXna6mp+Zr9Vkmn2P9Yk0Hgg/HblQnADfTx9nxe
AYWymFZoUw1qW0u0hFYZiRIZxqFcFlqClTo+IJT0O1lyuWqQGM2z3LRvanadFPu/QK/3ZsSwSmK2
6fvQnDLwfnBRTXvDjIfOLsWIkNTwdnv6AxdSGWI3S1dRpR/TT6iKivPHR0jSNFfTLcXDbbZKDRjB
Bp0fW7PuLDqr9gYRElNFOH6SKkCMhSDT9+DQ8sSfho7KTDN/WY5aJuiH/28PYbx5cOQyf7Oyfc4G
YdwvLrrKtlFygFvco3ZG08nlrcb2Vk3elUK2lZiFOA/uJlk0CbaMjeqAv28BOppdwt0M14oPZEuI
0qlvdrWwjEaOScBG7IRFFhe8k+vjjRSsIrpmGcbUoq1RTvXcZqcsJSSauP908kd+PwTsbE3Y02h3
MIRPmT80T/LrBpGO5JvMXBkSIThic1QaUt7123z8V84NelEwpieSkTgxY7uujtCZngwouiIq6fLI
yGqaEvR7+zrWOkUpbnaGWm5b4rymUkUprv+8HDyU3J7IaSu3fPmtj8eFPMc6D5me1jSrImqPF1sD
rLVv47bbgXQKdkeu+DRN7zeRpMWwCGdNuwXROV220GVs1getbIAMKWrJmOKjBQBgX66oqbm3LJDH
Kn7U6KKM8+Vs6LzX0Nayb+Gg//ZjGrDnkdQooISAcWcECZO081wD/FkRIljQe8801pBVzQ3Efwi5
typ9JTZ6EP6M3QwsJSkhNg7FPEgQXpZJQaMVuIqIPXEQ1BBbz2Gz6QcMmM/btSP7i7pHyZGk/JR8
UXNP82uQO9LeNcJPrRifC3KELid36nlPEPuWy1ePU5f1960xh4zlGgFy/4An07Etlh2uPlKTSXwg
OeKtPUIIOjMGjley+NaDCyO0PQxoXLKUes/eN4P51mw/cfXXUeQJjLJrMWV56WUQQr14Ro5WfAv0
InXbw7+FciGIpXBh6swisuTSkXBbCnUAFIZrgGgOtYdhneoDnrSV8yH9rBgEbyudwJb1memdVc7B
A6GlrJy237UPvPO1muKO3y9vfKRPJyxCEA2rrgjDke0bllANilGK5rJWaNvhb58OjAnEMo/IEZwE
1ZdNPzSGCBrQ9iwo5QrzYWaH6Cp2tocPRTchuUzS2lW4qITD6tznXZqy7oLFq6cdpbtwwTK39dLX
Zo1KvwhI6SWms0uNf9uL25oK613Tii2pZcgAvZnxEotoT8p0Cw6I5vesQ0vAl5T9NFB5eog6D4gM
3iDrFUhMvhEp32vTeuOo+1Jp/cI5kZzUSMKGMESlMz9KDKnBOca8uX+LJ5ELiTA//SF4hG/uFb/b
xGOc5QwPssRqMLCq0BdEdgm3Fk3WWGrL0yJ5e9iLb+BBZul+I58RXi2U9JTvoctVUeoGBnOOBVTZ
31Y4QtUAPlql2gZQS7LS0ElqmPs3wTVePF5eVL8Cpz0Cg4U66k3soySDsV0d3yorFecH7nz5wQwu
hXNEeNwdJuePqKqAiANbbgwxvc1S9snfBxNjqARKYSNwiEWcBJGpU3u/U6xd06yur1uLJZTprphN
4U/IQe2iODuC/w3bwvoSpNIW2lUN79kFWhTiFp+SXzbRq0u1V6eHzQViJwa73b2TqKM9Gqo00krq
XwMv2K1nFJqBI8EcvtjKBgbufw10k32dI9axOHbwvaM/9TqJcANo1Xe24nKO6Ka2xdnuG7YkOCD2
bfzaPCD7ZIqoGn7agjxe9CAF1cCmjCfvex9LywHzsDMm792+hfZucm2VgMf8sdOj4BlbVjGAgJCf
GLlI3Mgvw2uUnWyN0z3XjjpeWJAeldMujBmLP64DlGGeAzOoRQdDC6mLWWZDfvgIOG3sr/bCi8Tr
DSrOYSwGEL8T3CrPwUW3+P2XAdFr9XJWBMjyUfeWAA1Dtc8xoZZgHgnZL6yWt03WmNja6lcXjI4J
qcXSWsNbH+sj4dXft/QfWJ2GultHodfxniNiDUVUooAZ0vhxVBkUBkLU1/mIf794XCyIGjSwkRt5
EP5kisxbiCGQAmXxS523Wtk9LC72F7Pm/ncTi/h5UDAQmpTbzbpbdCBELFsSPFwRfc/5bXMsPXvf
m0zMJfcbVAwIh2OTK3MHNGhk6/8j4cqmO+UKAEHq0FcvpeA9C9VJMdDKjGwynS1UFy1Adsf34fyF
+AdUI//nOeVsH5mhccwFgGFl0XUN+tVMjdd1x2F2aQAo6cXv63qGd7VzCAzsI1z6UznVLBxEWVgo
zEnfZTX2T5HbT+9gFtC+lz7Ud4vQQcnSXP052TVOU7PQTIW9nQ1kyTvrkZzAIDD6vAj8DElwnAkv
3QbGbPm311Zjx4CkRlgPJdEVr7kaI0t19kRen+zKAoIlc6RtQM5KhtrtIEfGumsSS2NRfQt5ytAD
0FNeZ6R5BAMBMnmtJIKea1fZ2Z/cKjFed8wXfj8FLUE4zIKJaWftuulni0bbkqfr9ysfMm1bek75
FG7kKNHwx5dH2dVMRQUSEGSPZCUampBJaD3SmYQjcP3lPXJjbweT/znFcqjITaGu+VUVUwTBmxzo
VJ/g+e8fgIYBlCLEBTHbAG9JgnvUFqIoosZf1VAm4/vzp7BzAiSpyCdDUTH9WDh9uA3s5uJKAIU6
d1Aa8FxghhpqKumKVBKnSFKg7Qf2+h/EICR5dWQCdujyQlLnm7CoMJqbE3XeUFgPsYJ4x5tCtQhp
Eify3DeTnKknuwa5YafDN1ZGhVOxmU+eou5K/gsb7DY2vcM5GrLE8JchrFgQ+e6/oLPP5uRhaziq
Jy17fZTTmer3u05gBXfwjfJVlgfj0h/RRcf1gp3RKo/MTYAO/zDdqFQuzrOUX/HTkNDPicCBzTlG
fzy4axVSpw5JSAIo4HVgN4aCtsCh8/hpHHFKqU3gTxYsm40NYXD6PuqUXlSd20VY6cMdtWL6e3Dz
ooeXHHMi+qpi9UhzajMXajBp1T20yyIxujIdqwke8tsK7j4X+N+uEFXa+W7bf8VMLjrcFiiujxKq
53pDpSXjsXYIouypBnXari+xNntlLGYih5dvLoxnQ/88ENWhiMMaqfmE0EaodPkl/vIsm2JdlZOw
43P75TgkXhU90tp1F0oVsQ60FyZlRNwCsqjslY2UpLDqjtuUirCFDYHeH9EhAP5oxGcd5V6RmYdp
2v8eJsXN4lmUxYm+zAiuUPuG1gncSqmCtGl28SxoLTxcInKFE3SJT091qz55VHrIHdbYqYRSy+X7
EfJ5OiKw1GeD15OzmhsnY3Wuk/fCuNw1fkRLg1gGcyw22koX7TkeuDWM2CuxdrE8chvZbG9bNh0q
75MbWVhT4DjiPKpzlNxkwR+1j7OU5FlH5WikHMa5PlbxSo5d3kxwW7d+Fagzkk2ZF04ZBh/UXbi3
L2bkoTB27ogLsl7rvX74U7uYg0YOcod9RTvfRJSQZiUu67D9EFdaGH6Ftk/8DGD+2P4+PHGaH6OL
MHsJvvLbGSIrqgTX+egkITOe/RPrsmJXDCbKq8S8hq64a74P+CjeXnQW43mYhwEfm53xqQuXsyuF
yCRtdIRefq35s6AQSFH8gElDPuxLFb/6FPCEnnWdArWBx/jjqb/oGuvhJUJnsYAkcg+f3blyX55m
6N3VCr2L4adIGV312I1rK861/NT3xsQuppSf3xg1bbBHbkC0hvYk2Szl/WLEwajqDnwID4aErbY+
J2yY27uNPFMOUHL2uyPUxsLPwQTAmoNJfBrSXkUYhWnRMkJpMv8z6QWKSXEatSDPbXHDk/CQLFf7
bbdv6E3CkhpFdnLb290NTLveiwzaEE94vurFsFpOoqIjswZHIG9QJs6arqRpzs1Zuh2hm21Bw7Le
lyTTr0ejfg/z2SmEXG/uzzG2Fti/YRgGjJPe57iEUaTZi5q64xPjDc6UdCfFILNnfcmbql8OrlTo
p6pBBfg89Igf81EPSdLs0VP3Q3/6UpRicKq+wCGhXRGvOuPqXmJq4yExSEcKedgMdFJbpBE4dNzY
KzmLoC5eVSIPshKBLPLqQbR6S+GpGHO3hpd6Z6MJDO7q/5iw28MdG2IKTTsJGBeNmG/mBC952Pxd
GqKd7KyHJtrwtJ5wXfiFzG1qN/lZ8mZGN3EnC5p0EcVLepYVXsY3kvVgRxLNdaNdt+B4txEyREFK
T5Ev7DEkIoRI7ZL9F1o6GfBg5q6rlSpNk4nVNDMeI1bPsO0XTsAfRlzqoWTmow8Or0mgryt8lEQW
SuJXioA6ol/ouLAlRzKVmTweV+v1ZGYuJMx/c/42Bnk3LkMsp+2opMHuUkLTqSPVkZGF1fiYUPWc
pkk/BizR4czU6zNPkQzpClnv90TWC1phnAD08lOxccqCYzCO461r/XmBqYmOXQY4gqj7/ZU6VkGM
gFqBk3WBWZJxrBVo5sNCwl3Ow6SQDYFsfPgZnq+KxQRFa9v/BP4m7uYX8htGYKBB+61woWHP/Oos
EmvIq9k418RjA8CR/GfEJUNsbIxBDKRfygN1eIeQw1ICWpTH9SgT4vot8h4hQjsJ1WIk50byN9Sm
+Xe+nq923HDvYdzX0I+EuIbRobmfwJv5gBf79AFYm3YbgH++vzG4kpT8HwDNW0cb2Pchg2RMp1Db
i1mz/lD/x9kvlWo6Y7ad5oxS5m2o4RJ9/F7FiSzT3HHnUALjIdtSAOGHKUvE3dEz8CO1sZAFh906
kb794RGzqj/ajMkYbiuJFYaGeDxrO2+f7AJBH5aSumVPdAevZaM2yfjl+c/xLoid5Te34aOyqF6i
wT8oJeTeKw2iEHqsss2GXmGNOJV55Uow1ZdIWl94eCeNe6YUc0Q2WR77nBZnBnqmS9zvI7Vg5IEE
LtGpmm34Sm4VUMJvpL4t9u5SWsqfMJGYF0/i4bGFCBeczlDtyWk6ErkqvPsVDTmWljjkIPWtM7o8
P8JfWtzpjX4JAl/SlNqZ9/nvszFNpTBkOtcoahzEZ/1u4hASr6Gsl/SrTcyoqlOKwz7sHi0FIPvG
TL/uT7mWyjIRwmPdxZR7hUsh5lXd9LjI364pzebD6sPF3jMUmjf4snN6kyoW8LpCiRUB7vWRL5tx
7sPkIy6+oClQD8StFOtZrg7kDpwq4ZFiv62YkF1AupG6JmhkMjzmBdqPmYnShhHZk8CbtO/N/XXf
72G9qu7UeUredT1BT1sX1d0ceoZpJiSO7nYCmDSqATImJbgU24tgNqg+kTT8sO3Iw5yOQjCiYGhu
73nW3UiJOz0DSajvj9uqKwAT0BHqufbQeypx8Bkknkc17EoXkKr7KB0U/Zy7dVWNlXPQ6LdQeF6O
VCk6vOXZUlX8NMtRXO1iVbB1SpALODsoEvmq6dZ2qkdiXBm8JJ4pKdHTcZuOwXp+uG5sae4nPLQm
kDhcgFgJpO7fQ3ayAqAQKaGu+A8XX+9CziT4bwhFKPSvM1Bmgv3dLrtkDckC1GBr3oK5SdPbxoFD
gRJHDZXgLdbY4iy5Hjh46vqwMHxZ0ZkrNSAD+NF3VXjxe3NrCQ9CEbSl7Zr5tuZmAIH4ZU7+BlxX
qNR582Zcl3A5H5YP2QmA3EUY8dGC26QMrmQwy4X7v9DP/owU5eL9toJCNWYc/PbqJuQt6cit/Wkj
zW1PcCQpn5sNr4MyoSS7RkJcyg2mraJKQJO6ptPnC9rlYlJAb6e9/xGOdUAW0z8AdRwF+RAmxOe9
Sv5II0A5b+mnF06SAj42rPn0VHAqvRCkgAjIF8suHuZALyini8iZ1XIiDfkeb/WSpJpNUGj50izK
ovVF1PhGyYK3rfCrbIIeo1RlVEU7DCqP1eJBptBFnfUwJMJw94Q1EhToL5Cyh30F1kvN1MyTaRaY
fxE/d87XQRxTW1373rhIp0qcY+n11+WWQoDIUvvQfhab628xPmU9DC9aeAmyNcts1JOIMYq/NF9+
XAWqpkVOS/O2JIw82dNCLkkQ+ukZ50C7BweY2REdShfxYcw+RD/UxBlIkhDPoZyG28qcbwA2ZgFt
qZGxWzBIG7xiFJcSiMwWEjkoHGwvaD6fHkPlTMue3bDzvgTG4zzOoUfEKSofhQA7/gtKb0+582cp
sFTr36gGge8NDZbUOmVAV9oDrqrQRLrMYU75fxIIfrGazsKo3+KFcKwYtuwNU0Z54vGLShHjJcqq
YFDj1ujGMXlzlzV3O068jTzEU7ZO9E6NUE55KmAfDla9/d0LDkA5S7XdgsIAz4CKzYrEKyQSXStK
3MX2aDC4Px7JIM+z9TfxTC940KROfX1me2R5HcqfdahRm8NI35P1cYAzJ1OnnlNdgDRQuxIcOqpZ
gjVXcyr3j84fEyDxyb1jKAApOisxQ3vgZ3tzaD4Qx8r3FeeKiW6ie9l6FlJ36nV7cKApNuterLYu
Pdi6EYBmnFe51J5zIgU7XA24N4Y9Guwos99qe9EnctHCgvSt4EA+ryJUkW3+wFl5BHASYAdEx+Sg
vxMZcqtWixkhNukM0ashjFyxz6x8o55eKmo9nlQATRMzG/TYkq9S7XTjzrFXPKSIvw3IyC2eRUCt
StoAZfqFIjYcIJuxkWi95h57rWl4Pc/77lr/o+lvoBt1sxwOm7HAbmdpmTFE1Od3nTgkaG6jCKFm
uRuJasrSqFUSJ3P6/UDiwNH/JozoPinHJ7ZkZ6o4+ioqrqY2eSvvewaT42+usfPtRB9f9TxJD8fz
8S3GUU3ygNSR8CFOevFV9FfkdAvo+/aDNG2KILPQD/+BfY8Q+/dNA6Xdn2gYV5LLwoDHeHAA6tTn
VVKJbDAz4wUAekjkahHKIR7m8VtsEmuuijMkqlAWXg2qV7lOXSZMvUBr1D7ZL9thaBdBij4NNnDw
XlKghGj2mcrrl0qxI8X4KRoH1pCGJJj+5TFafYHeKZhcXuVge9loOj1WaR95cXdMKEmV1yfq1a8C
HumB+A5+VrGOHL62xKT+kEVo7JTT9CQUh7NbxiUXya5OBfE4vgObvg0Z+x1ea4F0KYa6XnxReD6i
Shx6NupBNQdtx5+merDF6AdIGB/tk/C2LoGVvegCFoQUdKGZQpay7d0hXp6GI7Oc5hrJr9K/cZzW
HqF2J6EOhNpfYkZH/Bp6C/wUX5yaoVJfBsRVTb3zvOFJRtAZJJXRZOOmzdENgBPXmf6B2Sm2+3Iu
uhVgF3uR6iQOkWh/UWQKp2Pgqg7QHECEeihPt/82Z5DJQwJdV2e6PpAi3flWNlk4OIz3G1YUfU8B
pQ6huCVjquXKt8387fhbKxTy+sNfcLAF3ZemGWjVOpyz20H6ZPAm5yHjQ3mMXJXXwCQ0kqwDANra
BTAgdQbKiGYYuy6lwbxPZZIHnfHaQ+oxTMiMIPX6c0ci1ylMPQ0B3VoOULQkoPRUmGGzLPlPypNN
+BD9BX8hRd8Duuy8VgH6Q+JqhJF5Y+xl/6vFhXeRT4/k397uaXhYkI/g9BqfDbxlEHJtLmrTf4EJ
8j28niLkD1NHD2If/9paTSCSNrh+H0qB6/1YJSIfiu/DAZmIFGT3eLK5RuFJNHwUCAXrBfZBrx8L
bW0u+umboVqxHXJjhgVC+qM44FShgSyc4zo4icmL1pgIsLQlqVC3fNTjX50pwwmtxA/0moSNbQQj
MZMFCksk3GmV7FFzegSo8rGfeXaQg3/ydLf+O6hVthUvvhavB+CxPLTkN5otfWygYaXA5xHhKEAK
xlmnikA2VgagmzAlEx/MsXh/1vmhkvY93y1pCKj/GuNbRtqUpQIH1HtLmuJdpHfqWCzktnW5otuF
Lmkk6t+VDE6KKr6lxfTWgmyRYL0rHtTDWJe3WmkSlOfZXn+8KhvzMO1YBH+pHDjCdwKzrZU9nH1v
+EEuXnT2muGujMpW33ziuyfJtnPAYVakAnc4izLgFo6u+EWmjzJr6XSC43fyTP88oJ1Uv9XX5o/+
p3Q3YHAfxqgDMU2Z4tcPAb3nc93CPYzWBOAyo4y86Cbhufmd7ifGIQOM3CLTrBqqksRyXrF6LQKP
VjqIoWCYzw7fexH9v+hu+PxngK9Pk/AqNkAqKuTKlF8WhsgXJgRAycf+8MIwdI24O8kkwXID2gc2
wlMbcct2Ah55QbkPCh6zMbxpncncBA9aMrqVF3Ls6Q1ydc5tsvJ2DdXJLcCM3TDKSuLLSZhDkGsD
cK6pAhBoVmD6+tzPZMHcN7r64JqhqrKrve6xNtsVwy/LpNFtmP6FxD9mAv7YurFEf6mvaMbDsvke
vm7fYPfjyjkso6iL5TbyDsMdM/NcHGEOikjeY1pZBt91cfmy4VAlGc92yecttvxsmZFsYX/933Sp
nyrO9wYcGj5bXrIzZOZ9PCzD31mOzOITGbbC6TC8yDAVL7fofmmvZdE7ycQgb85XjFSk81gaRVYa
ukeAfOdhJEXOssMYpSWf4WFxkbdfXu67B4O7lgATdjJpXPUoD7saSgpD59750qUbNBV7upZcZFR5
n3TdUx5v10ZEmYvghQ8K+ugT9+34qOR10J0x1NltMagIIohNSOUh8mjMUSZ8P7fMR5psqOHSut2k
CeOwd9NXgix43b+EyJi48bYPXiWVtfvzpR2MtC3YsP/ane/we4/ks1HnHmWR/kWdKIPCVSLpTXMl
b2UxNiHrLY5Y3AaWV/rsnrMRcnqfMrdxNa6RpsrnZibNHp9tZX6UzUeKfRIK3OqIZDd2C4lCFg4T
oDfVKzfEnYzwwG0/hYSfvs4pA8mtCMCA6ygtRTllt3SQ65RT+hWoflLkF+KZEcXBx09pUHHBOiIG
RDXh9W9abThXt4ed5Bv/o/5Zys4xb3g72nVb9vHc6IorCyZVli2eG0b/rdOUTB08zj/LpRPhsHVF
f6Vp2R0p38WGV/0+wJa54DnSZJBXKebjoBUbLnbVoDWuHgfRtcsVyUzNG35UM/FuypC1Fe0LR3SK
r5IuJbXqWwiaPR8xKDtBTpH5OPnB2+LmBlN3C4R4wkLrWPjlaMA1KVg2BO2g1AfO8tcximbgAlAv
K7fk4Xq+AS40TJG6RKNUaOItxa0ZAqbySYIJOLfIieyHWzBMke+qnjiXiGEG2e6p2wb2FDVFQDyT
oiIew63YbRCx2oOC2tTkp/NV43KOnIEJUlaBZDD51nQbWJmSUes9Pfh2CpYj3X1EHzamjfYLASds
82DSXaTCxhhgxSs592wXY+H03BogEfFc6YZVCfwBkfsxdjWfUl2ZtXO2XUDJNusz26DPGwClrvPc
46CYZz/CFHXHDQXugD3DpRAJPy6YKgAdPoLx09VecyW4yC2g5NOkfTfmHlQr7sq/baVTNiSApsJF
CXgHXWQ6k3KKfKL2S1RHFB8lR1jE1Fykdfc/R8Ia0FneyPovWaPEf0/FW8QpEIuzJyUixUZwv/Go
gwIcfTbdvRfhGax75kyod4D4hXcD5/mDChHDYmaEgwOgKdt7F8bLU9W1/XtyRYUzLPWt2Qg82KJG
U86MaXm6EYBj7Yb6lXcoTDGZfcUcViBx0euAOuEyDr9sFhnXxB4+Nk+seCuTNm+YDcvKKWwND8kL
kEz0akK//bTJ+NToOB2JgOSbtB6VMTDzUXPxo8FM8NonzhZ+E94YMU9zfjPz20he2J0gcdwT8HC1
nv3kBS8mXZlKwdnNqa8ZM1tsCIzzKH2WZGT9z6qkjEyRWF996/cw5eoqvnBuXJmNKUY5GjInd5yh
gi+CVggSgiRKZGdrDaBK/iUMd5s0/w9D29Z2yimDAn+vmhwmT4DZIeYIhVFXsV1lFdhkrmfrJSww
aLSfw+2oW9hnSQzsGAD3mFeLx1N1kodTR+rEElTUpf6tk2PVeOwk7Xj2ygTGaedtW3crfDtk7ov8
T/VozTcUWs9TG+UOrWWvOKyJAog1ZVHkVfG3d69viDmfDuv1zKCYg9GRvxodDUEFY05MjFL/Vcaa
Zsk7xkKDvAqi0nOZS/JVcQ3rGjlp8E4jpTJDRaZfeLY4cFCljCTG55qvs4PIBV+cCetqXswaqBT4
088BQyAcg2RLvo2kxYYw2sQzFdwnYkBUA8zYX1QCeefGuTywSOrLmZk8BdpQMY9s83C+M+YqxwuL
V6l4H5Kh6Ri9q1C5fYYUG4RI2O5xIBSFp0Su2mY+vPsuNVi9Ul1+vs75H0B/TlIR9HqMZFBbiABy
O+y9bwHpYAcw2UGfnAokliVvqysNjLi4ucp3ElAjfYBLwB9n464KiIffxqW0RAOyOIUVswCrqMm8
3qCVl0FJsUmZJ1qX87gL9dS9gEHQBXZVcTrLhAvKyOPsT4SQTgJoAASlXbAj7EphfVVHHQFCck8I
EtofwAfR1LmEVj8sbgIdQ4Ax2r7977qnBXq+9VmvAHvR9gpmZ89sKtsyYy3sAgB8gadRRjEXT7zp
yoQ9ZcyECmzEk3SLSaP6xRTRjHMdLRZBhpP9v8fIfx5QGItGAlz8MY8hbPFWHXkSFkUtugQR3lBE
TFPwIZ6XodYkvtbkJy658xI2LtYur4o7IAhNkaEtnUt58ECGz/6SWa2JUc3N8e9OG6UdmmK6CYUa
FNBxGXfL883xWmxYk2yKzIuOdLatYpE/lCEZ2UpeQSih5RuTQqnhU9RBTyW/1OXC1XMBqXWksaOM
rKfdH+Mu6XlJFf6wEMkSaiiPIitdHyXjH04lM8SVk5ZLYmfbRe0MqmhnZAl7cg9jYjaRPIBNESuA
aVzIPJN2OEsNX4NXSNJMb2pR8qrf8SsLL1611yuIv7rxqHKqChNzHB5zF3WWLpYDUX+DE73eXwcu
YZe+9Gm0KsPjMWtN9N7ivebk8rc2vGSBNgJfp9XAn165uDQRxAkM/IndTKll+HPlS2rNXn4VlknS
CQLh85u/oDDBeyTbrz56bHc9WDQHnTkJnq1u8S3/4FBOgh5VDO065f5t+/zZ6eeRJN44oRnKQ3qb
alkxAMsJmvc1JoaTDkLlRE65+XRUEDk/dyfa803WdLuv5hoZ9M40WCg2A2bHAnNf7Ha1g/e9wz8y
S/opLYq+k8Yw38mlH2th4ufHAfIU57oqkPDStNQfLRzPvBk7Z0O0KagMvOB+glKfrF3Ks0U//YGj
kEe9FNB0Exo4Ovv/Hvdw/EC1pflNor409VsmG6R2oQut1dF6AYq8KXnrjbHqTTB/SKKN0+7seyYe
tjZ6RQxKht/sUe5g+DjO9zHmNHGpuojO4l6cWgj5SGDaxl2w9c+skl1EP3Ya7JlMRCrIWXsQYjQW
h4efe5+Pdioyx0lUCS47uerUOLL25wTpWBH4akJwVR8pO+nfG+FkSaBJgL3QmXMB4zP5zyDQcyM9
uSXDGhZVfGmi3JZDwlmbHcOazOyfQBqoHiAgZCbegV/GMwGo3yRp1CkYpA5w3Au16PHhTbaIsrko
3L68SbSRTN21W9boo0Tn25+jEzNInHPZRHr/X3rg0S22jdtaRr6Crail1i4ueRE/5t3QeGGigasP
VRkIyocR9u8PtAyyR7DSFcRXNCmAb3iow5qqpffxPfO9gwB0uxde8Qv9L7iIdkb/Q4supZM6TeWv
ZzCSRO2+Hi5UGN4NEm3WWiBfUSjuQks6AtIxeCty/G8nkiaYNRiAKw/QPBTYjCbIXn3Oac4rvIF9
nD1QgYDjoSJNhuf+DC1Irblxjzwbc7FhKIDh1YXaQ1inlvC7kOoyyFI1xAvLgy5+M/45BC4JzzBJ
5gYwse0uD9OCXjDgU439GY9l+eQY7WvRKFDVs5WsGXI5sWLJGI29zW4qbQ4PUCPZCiEeFR7vFgqG
pyjjShEHmd5z+rFjGImSQB0PNa9h8jD6t4sdeYeXxMVUuugbenC6fABLCJcGjW0MoNzePXgX8IYQ
8xT5SLi5hQ2nzfv5JKsYzZxzDMAGIxQBzXyzVGuAYl4kgUGkRh3+6xZJYo1qTyzJYNlLLfZHk8QX
OvJ/+a2zRpDPLSjECwakP6sePQhtlawxtdtLj0xJbbahk12TqPC93nn/MD98z/SUOnU5GXHmlTXx
PyVZ0hy7/ER/+dnw/2ubhAq+/DS7wRL69sfDdGSIg5aF42Ju2jKzUgRMI6WfPf3xU7db5FaaTTjh
wbpLYX5GmNv/P5ZMvZ0Q6aNKf8dS6t/pHC+kIcCP0QNeDtwnAc8lacuBmdHU2Er6VsOYSiEtozVK
th2s7o8XrBHNIqhxS4qkCjLBnqhdQbI0VB6mWocMXFyAb6QJ5/2bMPSL/s3Rsl/VW4vwMbje8AEk
uDkrUcXzBc9XoeTAld9p83sxnucEnSCa1F9W2vq63d+KE5iu437wVH/hyDcxr0oMlJmnvjPselHE
3u2KuEVtEi2w2xHju1+RqI7O4Cpf6ju1mFyfYi0iMTARnSWeVgGkkyeg4ZKC+DrlvTbKuCmhdXOp
HlafWtzxGB3kPnoXVOLFgrkeLvGXIJORi04K9XLfLjoYoxNogU88iLg6R/nQM4TBJamI5X2W1pCK
C5GUQUFf7yDVVN1+gKN0Z/tNpVNaBSbnqRLigcQAhMNekzd574m0CIixIzCcZcHcMS4EbmPj5Xob
S12n6WNQW8PUOZIoSOunRMinpZr+lFZY34ztdY+BJ2lN17AhVlRYHjBFHxfuaMGGC67XVT38P6Fy
gbGfcDPNU7r7G1LraMCwzWzYwQrb2aWGHMw99CoposYeYd/0PVtXEewMp804sQc2H2q+EhQyIKPP
CZHbJLOA2KvBhZb7e45FJIc+t8SZfCiF+2xW6vpKH7rxcoW3r3+Q5iABJBHTZPN7g3aPMsHu+ILH
/fh+xFSKdIK48UnRKA2DHoF1w4jXNPAXH3Nf8SUWfzCgNad77pezlAU+6lDDQYubOo3c5VcjKxvC
C542kvKm0+/GUmEfolVSzlUXQAWkdfuT0JH19ISOB1AEQ7A9DRuN7bBRVf2b+rRe4rhhL35rp27v
yh3nDmx9sKcfD7NTqmURW4yZ01yTCkqdilguYmH3koDxw2XYF5c4jJaUq79BLdN3pTQYovCiNDFg
kJfg0Kg7NpKgaDNgPF8EJEm5Sf5kRPP/4qtm/pY7kFnwFFSPwpU71g9h6Tht+7Ap6OXbRuoYiLw2
i+RY9e3WshkUNPLYwAMTzdZPU9P+Q1x2Eofa+0Uv4q1gAQ3Cm5DfYvcOZt+EFJG47UV8Tn+Bh721
SfqJdgZ26XiTEZ/Nr7kW+JOo88EwyCBN8v2m++SYndPtz6T32pPk/a46lYZ/Y7SmgnuMZj1PYmm3
+ECYdPeZPdh4ogVfEMNoCZNZOH/kyCTQlJFNZPpDxRxTSqhqZFAUiEtGim7X3/6c6F38zsUGs0Gd
3/DQulhTqCDhGPvetV3iLOwAFErMQI62UEgYv/ZdJrRpwdLbEp3q5SDIrikfhNpXC2FOTXxO3NQx
B/RrzZPoLgCgiNc+iLMCkvekP1kf/wK6bcJ2dQNMM3HU+Qnh2t2dgQyKRlbJY8uHYlTDxR9MSyDN
7/z5gjXYeHvZTjHFYo93BDFzGxSRnGEoiASRx+pFznanVylwiYysH9WBes8SfeTFmFPoo7I4j3lW
gAc7eV/gChwM2K7l5zaOgNp348kRC47rRw8p0lw5U8fVqfgC8d21+mUQNEkDFyuuO2UfQnvuyQe7
BGW24oX5iEU1kBH/htJuSaIqWHooTpTyEQW7nakX2idf83VmU0EhsLSC3pJArosYjlZmQS1aL9wU
FOCmuudGWx/ezjuov5lLEgy6CD0Z837YGMCXwA2HIhA9c+JYrJzHxCdNXiN36e5ZNtifzTYS4jPp
TOI6LPytyVuJIgaGYCvXU7+49Fcr5B4+uxpYcbqsi3/TAZQRBQeyQCyE/HS9duOoWTqHVOPpxncM
OG0sW/OQlDjuHAy5xIe5mtlahR1eG7XCQPa+V927KEpUcojDEZYAGrECwqLHxrPDm86lHCAjtziJ
m+2US3pXH9C7ZKgzetW9GxPrkHU7wiLAAGrkt4kHl9K5wU9NQRxuvkULsXxucqRXBi8nmGAaeXA5
/YjoapsMSgkvlRvDKISnUzW0pOjcInIb4A1/OXmjLxEu8dvZTyvk6AikzsV6nQMJvqXlrnWxnyQz
Vt5rN3Lc8owgojGd2tMBFAKN//GEkbZXkHMSUvPvpSuOD2YbHWLOwfCFL4QvI1fNFAuLWbp+Oe6Y
ovXSRr69qB9QB6rKKmEGUuQtcmmRLxR6EepE/PdlcTc1cVjQzVHG9ymwBaV7kmryVG0+yRXNsWyu
ndpaej/7MmGmFXtygCKBw2DOb2iWSMaT5PCm3OkRcf78rGtzGVxVP/5juzh320tIp5BTW2g3xcYo
A45NNxUTqFbVXxKVkU+MZ2fsT+/HoqjrKIIkC4tMwyhM9OBB5hRNQlDYWGKHlYl1hl/sDgrvpV0P
Atj4tVhky/8ElUh7LPDiQR8pexqdcSi2JreVak1vaCIyMJ7lBF8OMW3DeuRxEZKjeLkzQljbpB6P
MJBHQ3GzqKWMhM5KdYpPhvqMDp1fgBugvFZ5yTEyKIuRc6LSfFkWqo3UI4DVpQU6PjYSlsUgv5rO
BwtC+GwCTbR1bUClvdLeEX6rBIZ3pEbR0EgVjkGpS3BX/PYbkIDEbwfYSnONZR75kq10cK6d4Dtb
ttJ3Cy4sEB3ZIEWETxs5B4aHXJBXqn+BQvsEQ/H9QuVX+Wr/CWrB8F7FkNdOFASoQbqYq3zBb5vt
kduE91s8Y7xjK2czbwlMUC8CVss1Xqdue132QkWevZ8dJDvJkQ2L3xCPvGw0hIRbM5xqUNf4sXIR
B/3Y4Dv6xVUHUNWXV360qM5iBkCqLMQc1z+Pl0z6eov9IM7ghz5xIAyvvRP1BFpCr5ofmVLPweSe
wsSI0z38PZadkiMRt82eTSg4RV8W5eN2nV6GGzMONo7z3cK6JMAhO3JYhKYz+DKmIfAqhtBQKAGv
fIKoXTwzEtV6cv3fUAcAlsuLJYwfeFrlufwW84YhgG3wpOzXEk+Mjz/VjVZ33CCDuTd5jji2Sev7
d2OM4nKbfmMxr+9sOGssjSQqE1+Tt6n7zhOSM3LpnBiX0dFgr5bBM2hNgxARt545ZNv2agkDgsJI
qN2sY/HZ5s2HwAkkY2d5XV6kPWTi8IBZQXqh1xV/NlT2/1Tu+AsdO31vVxyNe9eK4/XGMjVnqxVi
72GNQPi3/Fkxy18iorSTGiRqJJLEbWAHlvetI39ddT9SX17n+cwLsbd6N4SfZGZilcq+H1+FjnNV
R5ZTrnJPXsgvuYWcxu8H34fElNLNuZ51AQ0QYpTEpcszSdz+j8sEIECQAjTeXZL4m7yGqMBQuIj3
vWBrtygN77H6qUxnWvnUdOQxEc03CTNX9ynJ2ySXnjhzQlLdiRuhjxpRdSzhM/eLglA037oMKcPl
BoRhf/WZfaly/6tduR4SEPdwOuI083cNVn4Vk3/7ZZkpmYui7bDHquxS/T8XyCF6M8KaGaYlwa6A
fGYVTaw2qZGzVkZ4FAJrzEvSRnx/rbPUHfPGWhgKtkAOQYO9QGeXqB85bo4ZeYIsr/Xf1NmQeBDp
J+7lIqjXRrzZk9fK2vSls7WL2nigm/3p+WhGzy0iDnTgGBBlJcU2WA1Ra8PjbgTFsavBOEhCLwBe
JYhJ4yY9zQymnlvkepkkirB0UZG/HcxFbKSQ3+DP57T45IMcG7MJr2+lmphIGp7VRcfz4ZlMw4Il
RelJ2T64rdNNR6qcbHag0h9Ec7cXgwrof0hArEkNFqIbWmwi+GPhY+GaY01lEMyDxCt/jmq73ovA
/sGt8N4KhUmxzktC5h/0LyOXg+QOyiE6nlaIfQWXKCOBw9XH8DCPzRwpRdGFYSKukwHU5SbZFCH4
mFydYMmwDRxDJvkcTauA6X+zoiRHtnyU+kxk9rJrVA98U0yM6iMe6lBfTSS9iL+Utm/Fv+29S4EK
SxaeamgmlFkBsddHgmh/B8MgBrgMirJ2qddls0xtAxzYeSzsIDu8ECmJ+cCjzxnubk7joAW8AJmp
IVrf4O8NCzM6bTRHBTp+mrqra+e0zHy4rGHlCuAB5lhWe3DFdGOzTY5XXmD1hhLWZkuiKRyWSzEr
tb9blM9hcDT82GcLviALYn4VR7Fwqc4SC2rUiM4FdGCJ3fmGmj5Hq+Uo5+4yFuXx1Q4+UGd7kVpc
fbrTnWaUim5ZV4gXNPDdEo+d4zPXoZiLsQIjVspcXq8D7HXWS5EGHALDzZnfcQi2PQFbyD/d4UyE
hptW/QBybQ8FghqaiPJpmLLTohkkF/1LFjWEP8apNAqWTo9sqoYpNxEv5p7u8lJsi9tRFE5DWlkc
+VTNEeC3lWIKvKn9xWgnVa4f2fpxRNXPLEYoHwinQ41Vtwqc8P/RIHmbIpREyiJgx5jjzTSZNifa
ICP0g7tzxA8CK44OL5xtPI921zrv+EclKJeffDvMlkSUuYnC7ceU/xV9+S/U5tWsSb0lGMWuPwhy
C7xLnAGguybyMM1Bpsa30z2F1j2en6ECIzUq6TB6GgfBAbCYE0n+6/FvFnC8byyO6H2iGgNQPQqD
KbsXmGoZQBoG6Zc8g+WVN1eaDRLOQXnDAR4V3pHw7+vP1ePJngb2tf9pNjCF4TfWrx4wLmsrj4TK
7iNU6cb5qtb1GFrOISyYWVIn3rzVlH7Czbeizve+xm5LW3KToAOiv8MQK8vH0NrgXXa438btWJb3
k4CxQnKro9F8mH7dDI3pI+IoOh2xrSkG/B1PnJnSqWe68JGzaOLQkqyMdBpwyRqKlx3rF1Q5tDug
kDrbx9CuWgSgYqXUmmOTC2pLSwyKoXme+1gh+PZgtbiueXXTI/pvL300KTeJy9r6JULJJc0orxBe
jhRxYGGHReEssGowDOSkHfooHFOsCYCVLby5M/5TWi1PH/ksKd6+hPr9gEsbXC1ruriHrDL2pyoq
+4G0SXiu5qSLM3Ly/eO9FAZfpL6r9A34oVZwzJpno7Zvzmgwbl0CIsMtyo9E3NErUosxn9F2G2VV
ZlfBT3NCvJsPl7Hz/N4p+R/byqVIBjExkYwbDaqkFWpM4zRXFIX5yKozEcZZlVv0WmiYZZsw1Bcp
YJirXfLeT/2uXn1By6iFMmhJydmO0+91/xlu4LgTEquCstMYO2EQXXNnhRGdx/JZ9c2WSsP8tzId
Tj1v4QM5z/l9hOBP8IXNNE2lvYBotmGIl8mDn0jLssV7aO72f73I79Dey6ewWpGgnlNUvCuGmPHq
nuuBd/N8DqesKcWSS1JSqwfyqupg+zoXRdeMAi4X4pRYj3L13zZBuuER9VRmT6YdYZ8bpi8QCSiX
M1Yz3zUaTeicjnRepzdT7LfXJQYqM2tSKmUkh0ACgn52qNeETelEPU/H6prWzfK8pUp4ufpScYpR
tXDc8Oaxzt3qK2Lc/RDg50s4e7ruF5K73Q+pNJWY0nNVfGIjyEUXKMNffdKtUkFEAfzJbpWsP7fW
zDCTOTVNc/309SCL8+EFlctkbXKikp//B5yyy9691dHdSKg4VM7CXCTacl9DbcpKkdpe9Sd90nm+
m0DSkx6DR8/eVFZ+UH2uNEWyO81dNPOqMkl60BZqDcVOSio4q96XAn8CaNlGV3aBIBH23mqKPANT
VZ/cEv2+7gsyAiRNAv4zxmiNZUzHr1O/pDbm727EFaGptuP6aUmF/MoSPJhlJfFfRYjYN0cwHfuT
E0B5MBD0/2ll+yllIk064SY0Udok7Jh6IaTxUheES9Tb88KxsOvswDlpRZHQZzlxAO1GQa2rpOR9
FIDPe9Tn9wy+5EpoSKtKl3nXwJVB6ziBgg5qQcfiGfqMzyuVKOLY1WeBsSmhiXm0zpFNfy6fknKH
97hW4sP5Py/N8gM3dRI7rRXSUlAYEY3TCYTTnJYzAhRjmpnq8BJWVztSirmM9Tb5h+2kmdvtM6MY
zNTxK3btL0xKhNnlICilraz0v3Nxm6LCMXH32sP8Y2OheNlfvVdRbzyaNlJyQxqzdZMYnUXoFF5C
831vFGn4BTufbQP8QTLgeuMx6C+WZAbzL90cFalYSy2zE1AOTWS3RBPkwULBRdD0wGLgRepak0Ur
9+Z3qp0LCq4w0dIcL3kU3h/50nXVrjgzZTPWx/j5+E30i0fx+2lcqY+9DSV80+jeAIuY5/D0fRxZ
yDT0IttNkqYV5L6oBc222PH4UTlRa5xuUguSf3eW+DUuSWmDhYta5GeXsvjvDxphQynndBeLFjvN
08RcfM/fRzorSlzaaw+b+qRcF3zpZ/w4QLOcNxQgM9SBPFFheQRXur9JutflJ6Wlya/3/XvBin+e
8lhvnfMa4ENCojPAZVqA+x797qvtsBnQW3UK5n8GufbwWweiFlkDANQSMb9991kCaHaSfb/zYysa
UoLzwEXJ/Z0o2gHghEMyOSjAJQsdAVV6MZZ/sX03rG6JXr62HLwDydaxgKbb1nK1ICTYaitkLPTI
ydJr7BRZExH21MuMYKcbypZxHXCo9OtewUZM0bKdsmZCepNacJEPpHVzThqSggZgdiGVqhWKySFR
PpL6orDP7jna2VhUniWHOuXfMJR8wtjGWaNgeCjuEvqDaaogdqSCQvxaZUolbgH2fMOCMJ2SeAn3
/mIaLlD8b0SJRb9vdQKOm0iNhNPnPQ36JzkP2H/7+NGpgpDCEUpAwOr8AkkoGJuLBSK4WV9T7Uwp
1BxhDaMyM13KtEq3Nv1JltVyNqSsID873+WYxWeB89RllsoYseL+pBGKxOlRkHnhgnMlYDR4YNDZ
sG29SevOcmsH09tNswe3D08klNlhme2wuPaPj1M7yI7i0TWfoO6Zdx67HapNkVIKivQazueuh27B
TIYDfcATF7G26w5GCZ0kBFbOZ/QjrdtbFU58nU7+yIIJzLI8bi3G28oyze5VUIOSjPdqLhcjg/te
Jr2BjgdFY9r0JK/1rd+fa0/GFKC30SrsiPRH00kkoN1R96WycafbnEfINMEBVy3/Hts4boWumHtM
/QwBmyQaLoqvwYhRW5MYP1kf8M2+6mbDUIimpOJzbG2JYz6usX+DwpEsZ8AG498Z0vBYZYl8ndi+
H0u6CwuCXe4gDKEQJt6JDHFL1kJih/Za5F1W4Gzqtk8FT19lvI76g9Ty7qqOj0yVRGIbYRvZDDaD
dQl0klEnR4JmfUtTYeG19Tu4pEaBAM7Ubm9JmgBj7ssGcUHo5UUeqjZmd0Yi7M/3j6zCRqFJJkX3
laGfmtJwKhZ4X2lP1BfF6cr6A13C/lExMhVh/xUVXYmwIAPSbDTe4J3e2U2jLxlQFB0z0ogU/eAw
Mz/lOKXMpgDJnuQTDPJX5V6KU3d5BFhnNgdKV//hwTmEk41kfJErQnUZ4UriSnNDCfUArHtKf5rQ
yKzV2mwG+MutUOs7txChUsg6tFXvDa+bFC5IlTLw1SdBheSsJiDRWV4X1EGEzh4MNsNk4UVB2fO8
244Xz8S9aKvM9lQhFEgTUdykADMXez0JZlSqW+jD8WjU60ARQMhUMy9JqrkZrX+TmbedrannpONo
oA8Pu8vls3iZGANFdNM4rep8zSv7O/fWV4WXLg4AaeVJPEroMCFvUGhDqRgJ1TuiJCCOq++e4mZp
RFTvoRLAuwxLWcDNjPeNcYtHOs9L2PCTLjBl5Tulvjz76T0tSb0abL7WsGdGwDH9M7DDwzqPE31R
IuICVgusvkKjzNY4nI0ahmKCB8m90LJZbFQSl5nw4i+0EE7XFQ9fAWbY1Z0zO/HzywkrJe2oq0KC
896RkXNYKwKgF4V7kHrehlIrFwaB8r3pyOoVRzORRzY8ns0Y55oKM+hgk7ZFUnJe8p7pZNqqUZMd
9MmHmXlEllteydqdp/5usppErKevZN6EMsTyaIgrzwutDkd4QuVzwGFUtI3E5Ci0O67oWwBPAd05
YjQugNmqgrSZuInINou3Eh0fLvi0WRcVh7HXgSyNL/CIxCHvqS5/grnVwtKrooZpb/dYA8wgIEqd
jjji1QBIQ+KA3+Cvchna2lGuyFsxu7Ye47NJt/2PNqa+tVSHqQiDzdm4zajRgUkqQLKC/M1Qr3VV
O93X2YYKJpeuy16MMsbZG0Ui/JnIdLoS/UMNkrMQI56v0BeOm84Ry8ZFNhp0Kd+3h3fSVSdz0qj/
m7aRwjBmsmZlWXRn2woZ9QMin7cXxiPMnss6tdlgFMKtThvgZPODcwu54otj76VA1+Qf1WAKZYG3
Frt+l32qciC+S6Qjhs4W+3UKjnl0LoR6lrQuMp8PH6z5aBmoIf2vh4m4B8BGhU3Ok0tk2Dl3bZRr
3QPPBVTkaDtmWePYZH90ePd+yz4uZWeawC8jjFhnmHg3KGtilNf5pk1M33dDfo0fdQZ4Xw9ztDF7
1LhLOaPTx8dpEqhJROvLi0Nb5w0zdAnz9y93MuiUHoEb+ywc2KjMULGhEm5+n1nWSVpDOyfukVbB
Pi4q7jkwztDrGNTN5Jtr0BQ+SodamSyMzr2dyBQKsbdM0jAX0nASGYs+ijOQUG/e9gL51f97UYXv
GygTmikiOKhGxhv5vRnEDVaIn5ZyRAdbhJbPe6Osku4jBkA5E62fYbxnx1syoPINGJzGEpJbCoFA
CbOAdhXqTtTWp+r1lFUYqjpiAKouI7B8r/KhJ5z/kYH+bMGf2XIanujVb4F68BzyOYRpK+Y9scaJ
kX2cG/zLwQ+mvQkuapGN9AgYgkwXUxG2UlRa75J5LDgCbiL0bsHXD7A0yQ1lZa8kn9sgCew9Iu8I
edZVNhbKAlbunag2SbI/i2BlMeYMe4meVYRg7CkS5kT9RradY6XgsFmcZMwtXUqQPgQH+5efkg9G
MzA+rMLnn7gu46Ry/YSrKdnqIAjm4dK/Zo3AUcD8E8nOWSU16K7B63nxIFaaaYwJawmWo4ytex+g
N6jtsfRpWU52IL8d0VgU+CxMqDwBLzZzsq77gsTpg1NhQ509eWvx7OTB5udgnFnK3gc1tg0eRgVS
NnbTkBaq/moZwJFwHoNWjMFUZuwEzXDp2fY9u5omxAIMCc5SV+g9nCTCB8ZwArXyr8A1tcg3qqwg
BOYINAIwyOIxQ0eTuwCRQRktvmFMvJHKh1qRKVtqlGEK/jrU7QJSW0oJr+9jle2YqL162gj0fvPG
nSkIZfZcbWPvT0FcLb3LXKajBUSGslni4x2+k0S2EIcyb34Jub/nv415fQpccHNLOE8pr1BZHyHH
oTh6SEdy0j55gkDvy1wdJZj+bVznCvGF0yYtuG4jFlleT6hxVrtWkvwTEmuSzMUI7h/LHG+luu18
aRT3XCxjDqej0eTCYMYym39ZB46BZbJNam6Xyr3mLk/xMiBT+t/Vus4jXjuT8Q05i3i0N+AbdwzD
LwcrVBdttg7HeAYf366OPHpJJjwTnCE42H/TfPP85sXkDZSK1iQ9pkUU7ShfUiupHfxb4Mxa/0+W
mg5v0oIjbSog2XNRijV3ZS+fJ4th6SAiPn6lZnYSCNJ+QX0KIeKeLS/Dfsp/nGoqRkZw6kUkyqYJ
kyPpi6hZ0dj/AIABDUXGJKgow7Y9AiPN5t+V4xJ6rh2FcAJOzkKcJEPSxyUz2IrVM+C1n0sFOjZa
4N2avHxTbhuwbmFaqavoF0IJXEMdiq2rdWnt3RKyec799SpcFuzLfa5AZJsztyVfTIQHM60Estxl
hEoWFfh8ahzWy3E3OwURGXtT0+//oiRVSeggqbrEfZeg3J0v3OpwotF/Pb8NliI6/3LrjOvf9xON
FKrjIGvg6xWqZoxMIq5jbbh19Jh2Nb+UcnrfZAYcMIrrk+l2BA0OjwOSPZEnpp3CWerA78SDa3dv
G7sai3zsAhhlp8su9xycL/jB6VBSKgJo+IxVnYsSdUzxVUwZGwbooqflth2ypJA5YPEwV1aXwcqp
3iDiduzp1kTJWtir+2EzR7pqiwuClxXy/q1Wa/uSOXUGlusoc+eEOucvI6EMEYM5mgaDqF9nodmc
+g23UVyoNOPs1kIC8yykaEfIUVqxa1ysK1fk6i8akp3mX1QiMPEMzeEOhaU9f3hKOqgQHASOIrXe
Awz+lP9egXrh0O9MeHWUAMXmcl9iqkL04oJjutOYsr4ALglb3Xj+Nb/ZXxW5hUxG5fJmBA67uWGG
Ec6Ey1JiaQahzi+yyOIr5i3ICIN+hFzQ6ToUvqujc0hdnBug44l0XJMn+n+TrtoyqWTYbqDFgTDT
WZgNlA+3J7o20giIQX/85Ro2xysCg4GhZK4WugSYjdxDSbg+yjmDakWvwsrraudlRFJdd+Wtkv5E
GtIgFYd6ZEj4ssIU0Mh1t5wQa2Tdot7XXxzQ0sPyng+v03l0dA+2IX4IiVBcvSsRrMWOI6Au4NhK
6EgjGogwmK0zLYLwyp5uUxaDg2O5laMwK+DR3asXY2sZdw7STK/tLFpKoGU1WzmBnMDGkaaNv/A1
348NSbYT/r01R3K84qeIZCkj4gUo1mHjP+nnaVMKNC3XjIlb0ZndGTBedsMEnyhs/OmC5+J28TH4
miPdnMfHV2xcTuM9A6ed78NSJnZLjPBNXLmkI9Pn0bmJkaloSwW2ogNqlwFRZGbIH2NHrWjPm+El
ySps5eyaF2r6P48RPfgIcyEiPjQgjBD2mfc3bnfyd4dkvDRFhF3sUQhMHa80PL4FFAkJZoj2T/yO
Ctij9imgqzA2fZVgsjr8rUzZoX73sr6rxGJ1+3Yt3lN+OVuNBHuTKJx+tCtviShi5PiTlhfzniYQ
6IcAcHgSBBLinWjCCt1RER8SUhHpLr6dV46Fx0BxqLwBzpwm6nLW4+i/PkD9kiKBetvoXU2DTIgI
pfnspObmFxRxV1Sc0hg9aVUWZ7X+1405MXJodmomqCvi8cycKMudcfcPkSsKjR574binaCqJ+8Ss
Uo5t+cDxnlefBcmlQem3OEO2DPiHGw0nhw4fStODzJ1uvzqICmGwc06Zxi+48or75ll4crsavhXk
u9sW4dIeu4WgPwVK4jfRpCsf0bYMtnjpI9Z/vrL+Ifv4GvfCJNiZb0i24luZ+SWJtrkvFEWutFbC
90HdoCgA75pIjyPySnanuBhV3lTf9xm7tAqZcBgYGipw6DWb8kOrvIM/hoc86fp935Zdun2/gVlj
c0OnpaT99mt2MNms5Tj6VyifYjQ8Kq9nzw8PWSrgeUrxiFHMaLz7VpAmjenwF17vMAuHUT3/wzxb
VfxvCXtimdiQpRM5o9dQOrnc1qNh9/WUhMiWhd1lkZenRRbSFuYG3KAcVzIu4jTpt5DLYOsAQWlA
inGu9vVeRYyR0KPC9MBPpgxrbGZmvmLtPRPrPM5l4e6DAZJV8+suD9zMEbOuwPL7/I7a+b2+Vj+U
liZaWVMtq8VFWRTrMb1YrfvVfCfwPDv5M5sBaqFL0Tzu6W1PgepQb6SPvyrR7AAqgtwV7r2pNh/6
Kn8FbCu+P5RrMYk4I+oRpkoRboNIg1+HmlqfdS1s02W6Po6cJVxvH7TsvRXWwkPqdRFDGV5K3Xsu
c6aeLOtO4KIYZGQiBBcM8W/cqjJFi4p44dggkLUyWPOH5MTqJqP8mPmsgWevoiYfO9Sdtzpo5gvq
Zcy0xFc377dKxgNOVEh1WVfUtzmrfbxxAcgVOsQ6yYPMAAixBRdIAsskhGDMQ5AJoGVlGy7pI/Yz
Ch37rEsHoguqa7E/Imf6Wq48EPYpSgkLWZSKucseWXhI1bn3YsCdlRvWHy5Yu0x+sso+TL4FURH8
9I7RoEQnst5CVxvhiHSuXyBMnvgT1MTqSv5iyB+G21mgF0vmLGiUPcBLfPj88UulelkfIJGfVzyP
hH09JkXfMI1O8xOUabSDkyvERPr7SjDAc+/JKbyR1T9E2W/OTHANBNFZU4vEf5RYqZj8fLJZn9jr
IKV++/P3WGVd78FPTjxB2XklMBVnFR1zCtsjF3AGk1WAN4InsqpsiZm07YjswseUoCS6d2O5Z/AN
Ms+89fAYxtkoMDp0qPQJLncxhg6SQwtfoV0D3UhDQJmmqwiyWKFBVkfm2tdKuzKNMcvBRRqaavKh
Ju3Z2UF/PN/45yygH8NaQVJjvHWF+7QiSILkZHi4ECJDkPq1GHL1WNZ4C+oh/sl8Oc9Y4SIyNfIa
nmu+GpY0qeuHL5PeHWNXLSkg8tCmCGnhj261yv1DKwOUJA+uOMr2uEk/ZFLAR75+iMnTMfOD11OW
pZdf1POVUzHq0B2/uImFdu/kn19HCl/n/JfJU0vfZh7zk1X6e6bZobAOVvDupAsQurLi9+kZWCzV
5hUMv3GBsVjA/+/Jy5+Vhtp6GaylsvR6TCqMBTrEqBIiy70S1JYArZzIFB/2b4OqrKWfU6LMAyNb
jTaQrmn0jHPPmFtTYXDS+G0ajmUEV4KDCiMaImfp9bdSFjLozktgY78Y/IL75RXXOcT8iEgTj3jJ
COwLSPACndBxlt6yYtpJeMPd1/xJUoJii/RiUtyKjES8vVDCz3vTe3r2e78OXipIvIma7w5cOaOy
x6ntdF//KXFLZRt3rmSVvFu5DuCDpPFnrsk1gZ3ruF1rnrgZNKX7ChJfPj6N9gcozxGTgk5/rUS4
JRXcX+Kgn/5ONb+cRtpkOugjV1SjPVhGtmGDL9ndgM+i3s5oXiM59U5oa8CgBrgOe/cOBmkaTLXh
bzOL9y6hAS/9/zD1Ps+2hI+lV7mJa/eDsTSF50X3cZsPjTDQhnwoh+Htm0bRjh0jaA2h4cJBqLy5
EQ44VZcAp1SUYF3EnH3ATX/6NHJU2uUN7U3YoxB9fnL+CKCo9I9l5kkHpMfteVeGH+DrKw1SRnYX
qLeYFHCEGLzJTmuNW6UVTeE+lF3tvNdbxvtY19LoNIpslmHZju5WXityIaQGriX/VtIrNhwFuDpW
c/UKagZa95MoxO+Tm5sX8mKE/adZWUp7esfR9c7jawxDcsX6D1Q+fKG3izvSxCG2EIRj6KNuFddz
WXo8FnMmHMJdi0h8nRn1fwBNQf0HVgSMBm/8wsOPF88ZsqMVMOlvlku+BMcEiRIvotvf7t5c2H3A
mvVkvdwWDn8w83HDBy2hfmg3drdlikyIJnEYmgAGGpVQ9wIbmX2iQCIVAbtqo/km8s+1+2i2QBVK
o5DYPcL8XO/E6V4F59clW1Pg8ZMt7zevgqb4T8B1lm75Cz8yL4d8dxF2ZG88gFwKe0EUpqaIc+uO
J9itKvK2m3FSIIeOc2eqtPHc1EVq8klWUn21oYxE3Io8XbLihNhie51fSf9c40+RP/bkCgrECVR/
t/nSvb906hP4RHEL8wDfLwG1qm1JzTxeDasHcMz3MRI595+t+B2Ua2I+MCKdrs6CyMzJ+eLt0gYW
4WFdNqEbCc4BDcpgpDi71HmZtAhzSNKa8ZkH6IS/APPQ/L4y4yjejFARLnjg8pZzLjbsqop+wgwe
IgrYA+jtjuEgTEZPRIbVvJXHO/ap+bF7UMXzQ1zX1VOykpQiAhedwZTn1ZGI0pgr5mJrOvYtvejh
oQpR6m8Y9KGlazSaFeH/ZHRSTYYtOVtX2SUsAjvBgVfbL+qvEYXbuBNsbdstStZjp7gukZPCDEVF
tBpFhub9f5Yfii1JbTHFAFTXOeHswV+0GR0fP2YFemdx0ZsKIrefw/YIfl8R8V5evGdwH+aYbFI2
i+lKPGc3zkgSM5oAGRrT4jmxh2M9+WlYFLnfy6rhSTPCxwcK33i9n/cBjRKIJFThNME1ZKoZO/yB
T/tHd8/E6/DC5JJNE/Qgp0NEQayAdl6KpdIrKFz3n85liTwfyRSTEiG4ZtRbtvtIPdhL1KUC9Xak
DKzR65+dsBdbEkWrcXF0hgolzfbnfWCVA9QuDRdfCmqDDOU45EA1Lf2Smlbq1tLRQAhuNUW7Yg0p
9OVAqGqm+n0Iv6UWu/sc3FFs3i0afH36/R74NRA9nI53piYymUlGY2NXKeqeOC+d7B/ja7SOEPOU
ERCWEtEOa6vCXYYQ5/8qb1DDAbzI4lLl8tFPmr8X4O5i0Xp7Byi2EiB2zF3sIl23I1e4N4/rk/GD
bdZs9bztlY552Vq76YIq/NWpsNLR6eMh7MjBLfhf2SEPtgkSEkCQvG5Ls9Mi9UcjClB/vvnOlcXB
r3bt9iU36bECyDu1iT9QC0FaeFya3cgv4MQw3NWpEbWxdOhartRKqi5+Pqcv0Dr7D42ipprbIQlZ
yumolrACyzbaC/LpKmqwXpw3W+wa8yjcCtj1j4zJKpMUSObxZARW3KeDJOxHzjTWqLSHV2mfMK12
UBlkOL5Koe2IGdKAvWR4WubU09aWoD/3+q3XwAA5TH7KEtibVIONb6mYR/62IlMLT80e766piIG+
m6RdYTCqsLDZFog56+F1oI7Dx7ldZDeFSVDymeSphUwMzAn3rsG7eLLKhlAr5gNUuyXPHaa7rYAA
ijx34DN9n5INEP8KHbewqGm23xIAz1I7Ul6+ucLhLzNec450nk8GlkQGPcDLeaH1fCjGvbxLu/vN
3+KgUvm9dBdxKeu1peAxsSAMOnBZuJo7hb85D4QfmP+leWDkljL4/9ZhqeEUy9QP2vSYKBZ4reNA
4Ex7x0bjIBRPUYkuZcpW8FVorT1XrO/R3f8WThdFgEINFhDn5S86ju85fkO/w0eXGy1lyCSTDMkN
K//y+YwiOzSvvmicFHvf7ntZwVc5U8kH5U/gSHixUDSE5c3OiC+Iq18ZCxg3ZTBRCAnU7Ie7DeQw
IN3zQJq1joknLbOeZLENFLYuVVVwcZ6Dm0qmiFWYbUPxZYmYFy9lLo9716gYgT9NZ0ZYtaMeCtFl
gCJPthiAx4pruyGiL2ZyExhiZNsszpDGT8OzdXE8Mf1+fgbon6iCBayICFWFEXk6mY6zIqZ9Ep+G
NnTOOVLQSXSLiV8OCYF1r3qsa4FwaJCvqtdSY2MVlHT7GM4zncgd5HSxTS+SyS9ryKOWEaSG02Fz
J6fYFkeey13dko7J6NGv02AeCRGrDV1REvWv0LVYpjeNld2+ZCX6r0hAiqntBSWs4qndckkK++QB
9rBA6e+DCMYzJ+9suKT+CrluMEZjdBl0MefPVp0fcm9L9otc+32k6FxrFWMiuyx/OagrO9xBeVW1
x9lC4hS/EMhreWh5ihJVl7oE6jhwsfmoz/Ne4Z0yCnjh3VsNAgU657MhVX4WHNJ5zYcSeXF0cydF
CXCzX4orjp0kbrs05JrZb9ggx8DeY6i3AVyTUBpQwr8KdsuYdjXC+2cn/j6lWK3AjUhAAj8zEudV
CHf+DXacYBqReh5W4L11j9yutWtcCUxvDvBmpP3H77XmM8W2ggNEllsnOesktceZcM8k6L3U91Jy
h0FqG1OGA5ZvmNnCyC79HHnZ2RilYF2+C4k9damFtdvShwAccqQISzwetTRBu88A7KhFQ+YHOkxj
Os48uXgt/G7YFUkCpqQWjmRmo1SgvxBAD4eZhqSfHEpFoljz6Z0dLG4OBqRsH6V6a6reOsOHLfgv
aRk3h6qRAdd8eZhUoxXRxMZw8kLEOJppb2eLzv+nT1/8WVX8ipE1QEnDdeHVBsFTLtcGSxEygbKa
fYI70TmeuBfNluTB2GSArlVuZnBIKkane5UfK5Ii+FRzkkYs/fDwbkpsKBoo/hcbrjG3DY+zNfwt
g/neVozTdCcMqzAN0IC3Yu7XrmyLhn6+pFJ7Frf3Nhjypg8P9nL9MmLcT4fPLR7SwbOWz7XpwTrm
F32HtiEZNv1BulOTCHFmKHsjzIoIKA8tfukQQUjZEa8+9wo5q6XNqqJlZP6XRnd5BOZWvIByAyUj
07QmJEKUmBHmjW2kgIwzRZl4g6raZdP114gOO+0WM2L0rNE8ixNHhfiqiPVU5C9Ft5axX11yi2Tg
lIPOA9k6I/3QiV/cjHAHSTsO++VYWWpY+9n35m5mIV1DCTq9gDPIfDHjfxnIJkIBnjZj29M/k5A+
b+JaSXfz2Y6ts5iz733Ks+M97WWiu6x/XArMBuI221EvHvcg0Sh7ONSVcipE2cNa80ZIjllD7Hk2
KwtU1DmmEYOPavnwdmXvp2EHIo7G1i4ijguAZ8k4FLqW3pmVa+Wpue/cdk2EUvvvv/dmnRwQIlgM
ijhJP5X1J+0vze0dyCkx2OGRKrTQR0j5rrRUpg25pfnLbhCs7JA6Xob8cSDBlJY8/QA6cxKnFUPK
RqR/4B5GiqFbkpPb+aMWf19VNFDsTmTfH0G4dfTT+j5Sj0k4Y0e9l90ouH1fgI4WL9CpL8vtlX9Z
KBGGVC70gxVA8lw9qHr49ao7WWY1O5HF6Ykdx1gzS5kHxMI703M95NxPsGs3lbMI82Ln3hRXrEea
BSQzswGHCi3nmr4dIjanmmOYBpJ+fJsg4E8fkUUdW2taS28C/K1VHUjNGRReoO/6WEfQtsB22h/i
1/1HnjUyNfHs+++Owm1gFfxcmoXxJF2deEgSZpE9Hm6nBJ0g4exZSsS/ANbN6N+/CkWyH71CFJDl
xsU/HKBEPRPJXu4WjxdbZkyMEQtbWPyK65ZLb3u8aZsxqU9cNscwcWkZBJGQOjQf4l9uywb/4eKK
EgN4Y1QPaYefVzoModcEG2kH36+cxVncRpTEANE85f7miZHUDdRacTDWP+//p3EVqIejx4oE2xsk
v8495dtkVlJM7JV8as73bxK+L/QEQUksJxq2qu9aKU4lsWtvNNV2GWoOg6/ynH9WDdkxNFe2eqIc
s4gClJ1Du3HSWH23XyjcYPgMCTWT1Xc2qlY06Vb0aQKATg1sw349l/ZtqDhLwsixIStRMqTYLAjV
FHoxXzZGYBECsZuyGE0cDJptW37v4mcEqoSIljrIdNoCqqqvkQkjmYYlkLfCvdByMJ86kOeu0pem
fcbpl9Lulz09wgNtTtG2rveJLCUDJx1d53TIfODgGJWcvi0VGybTjfO7UuKyICsAyZq+kR6b9tDs
ntua8vqZPLtHTwEA+9SDCrKaude1AVUIPKdXcviA1p8uFzGMiL6h+aEdnkL/VrATBbMPn11vuSHA
6u5IuYqUO1iBOqQQbejkbdjvC7xPrCLrYRMGIGnBvsLVrV5YRGwf53elm2Il680bL3uKy1ITDP8I
97YDcRPJY65K8DcQNzlhN3nz7rZ2A5YTaY4XlGcd/s8MtulwIfgIyL4prf9sDSuo4JNGlvmHHtDp
PqQ1pdii0e89S5k5hfsu5QgYBMpgKUWTJJBEqJ7jsmMrLuqqljAfUGW+/RGhUXSmHVBw0w21I+fj
EfaYk5wqe1oR/K4WYjlVv3m8Ozpkk6OGNCgaBIzcOHSfZtca2BhL1NrJU29/VL7VggCAUYjJ4pF3
iGp5BhWSBt39OQRhVzwxtD9ZWleDA8intNpM72I/zfFJ9pei7n+yhl7IJ3v92m/c8O3HcYzOoGnj
0ofVsqeXnpoH5fgCuvnDLSHDaaCV+Ctv9Goh28lLqYv+sjOBWzaeitqspvuPeYZd2QYlkHXRHfPo
0DKV8a2DfYcdiz1LfMmumnqkjpCjcet81ZOzM30K4lPOJA+LhoDd/Kz7WxLimwbYntgPdlQEPgdM
GiOiz6OvTGx03TOmelfe+JYOSu6/NmDSqFkebONc3aTXGMmsvEHJTL6E3pwkaQqj5e6lh1XKVyNa
TlM4Ry9vT38wEQj+/VSOnnlc7hO+i4cd++tkB3seX6UjPLbN0m2GSAKABEaDMH0BIUwMNDEI3iVs
iPeEXWkbW3s1yNpRCEqT/zQ/xOvh6aOFij4a6RBKalEt6W8/tXbOt33ERE9SwtgTDYAC8m7IL4fj
DUGEnS1/lC6hFUDL98ZM3Od6Cm6YF0PEhZTvYJ/l/XN9jG2Cu2nEWO5nUFJ8Bsa61Z7FJUfYDj66
2lX6CPSBCAQGkPtiYv2PhUFBEfRIItPK1VpfB2bHg825SdTvqd8Eg6Ir0UkmyRHtSJhFf5YQujak
40ULWenBDs+wjnmzozeSBn35ioUzDfdjWWqu7jbcDQ2R35C6LqvPjEH11yKMh+Rtv6E4/kWnyrz6
S4U7ApStP/K0QzCij7qXaAYviQqDZRt9M75a1nT1/316A/yK0oiBs7bDngNlfpPvU8/jbh23KMCm
v+83cLgIYjnjoA6bJGfuLWyuUSMp+tO94dopTGrT2aT4kGVwiFA3BNt+XHVJmXQ/Of9ciMZTqV2G
5RuZqB6krf1dUKJNUONChn/pUmGzbrZ0Z/gjIOvVXo0vkfwslZ2v/XhjVPNJppUAXaHsaIN0djhf
5rMFDemDXNYLucbjE7Gt803baXKyP8bg57xitl2TWYkTQ91VIrdfE1MZPEL5UnzO7fq8wHHWlFQ2
ucMAdZ+H6Ti92xL8x6mu35VTy8zNNBuD2/tdfCkTWnaIHEt19knOgKZJkcx31r1wDRciNppTdRwc
NJf+TaZgllP8y/ZhvNUaPNWhmB8GhKNzvw3px94PyvNBQP9QMg3cO2jjRtNqPkLgpMeJzyPQowUO
a2jwz1oZ63t0YrCuN1qol/H9qtNfRwvWJZcRYRRkD8oNeXLLjhexewMrVP1FUyYIzQ5Lhkoai1Ls
KTkG/wxMQy3k7A9Msil4KGsGT36ZvTy3WTfElHobZHbHfwVCylWBndTiwioeHaQovFPIx+2pKG2y
hub6XWxi5vThfT5iBFpR+t8UPkdWPIAk0nC3rB3rLg+GN2SKPDWV6U6d8YIz26/hlZMkw5WIkHin
GpqsFi+q/bWKKRO31VyvuPgi15hlkitge2mkE5GLoZb0fA+2irHqdoNGI8OdSPxDvCmgp0hT8slM
T0do9lx9fJR5Vkl25vFIJGyBTtnI/ByR6EmorlD2qQeiO1iYrBWL2UW89az/sRtjM5mJ0bzCKT4x
DS3VC7PiMheGxn87kEOYy3dNepZEcjzxRJ34c5W283ilw9yevPq8AW6tGQTklrVCEX2ozo3WEoN6
ARXTStJ6v0t9EghSnZQoc7gIMclf9phVM6E3/b91z5JiFss1qQxtd/ZZSWCsXIpp0IpcabUQslRS
T0lmZR/Zk7iBjjPCLWHGT1s7xupkOQUVLCGnrGLoN3vdXAKTZ2xn1cJFcABrRvh3/6PVI7Ex5nKR
PjQ1Axo/Bw4uWl5qsRVLyk9ZbD5bbnsfo6AZzFZdmnsXUlrfnGmOadWb1EF+TlWmLRKf/anPiB8X
1LF8t3u4wmOstIeSS2n+2cuFPmyGbfBVZi2u9ZATerARWoB3U9M79YxKB3rT0O3y0l9CtBfrGMmD
9RzMdlmMIiT1T04K61OFMZFGXnlhPtpWfh/+dIeOGQojN7zhpuBOboDuDRKfnUrdCjffSx7vrvrP
xI8PO1lRvUAKlSOPl/6sKkp9541ZGGCVKJN8GEEo6Fb6wqpLTXHfjMMeDokepm5MEd8SghLFWRQS
WkHVAzXeMbpChETO+Zz8PM1n6d7xYeINRQl6mnUs0DjKyvdBRSwxU0i/QlNhyGRgLbhtnGUp4+HH
6ygYS8eBGeZ5WVJNBRVAE7TqdugWAP1WuLrvmtt4Lnms1RGu4TNSRIdv7cnH3zLB+KN7He9KbEiu
y4ftxnVRCnSvzwXdffCSW7K6BB6gKJDopFYQle3ZcN/8SW9nQHY4c9NGgf2tBOu98ap/tCdXZYIz
0hswuKuHn8i7kjhrWx4oqeoGk4VbONAQocI/i/MpRiOpSMiYRiHd9XZ+K17xJS2aG/W/UVFCySGA
Sb2sQb77cyMQbBsDr4WEpszp4ucTMUrbzNS6lZkZUArL+aRlVV6cIMgrYo6R/6Syc01C1LOhY2+X
XWixL/N40YEFbIrdzpzKDTLJzknGbNqGmllxBmPqAwpdNE/6XNXqr1pGFfeFN8uXR9wyhUSTlNjR
TDFLnZ/PZ8dKlBbUn/Omkme4X4eeTyyS1SJ+zCBJCW7+HwvMeyFn2E8J70D2W4f67QmOQEJH3RM0
Nm1Lv8WQ+NaKKKaTYns0+YJvwcCG2DUBmFdZcu+Oh9oPvDW14H0m8vjW82J1/WUDvIX8pF8r9wRA
zQhHLkiFlUzJuQYD/FphVkj1bifheV84qbm9xpqg/VXHE/s0V1eyEXm5i+S1R+uJ0OmeYV0QDgS4
BJ+5/2JPV7NxYo4ey5FYi72KF4qTR2McLSUcmXwlWVkTYGEweDTtlKYsbYOW+04r3RS/80zkc4oT
KDhGyHq1OfbSw+gd/YTK7A2izb2vDHNhhRLQNWZAVqpoLHYT1xkRkuk0rrCUNB4Be483qVV/9YMG
cy7Ew2/e3oX5/NLCHVUBWuKN/ZM5rDylZT1BwUvEbaY0Qf+luP2mxhMcBuQ29NOCeifMr26Riabu
GZJPXOiDbbysSI06+Sovh9aSsRiK2QS4ZpVQCNeT70eCxR27eBZg8bfU9i6kvIP42iGnB6o7Op8K
ICBzNAyuOSLX8qmwupkLas8nMN7F8Dn6v/s+5VVBxuMps04mn2LOcf+APMZn+vtxFPCommW+2Fbn
08JGgKkjYcc2CWYNys1uFRCMk9x1u7yyHY5PrWDrmTijnkdtYjznuN9IojSnXAYfGI/Fv1hIuyZ3
MRw6ZNS95IN5eCd559ssocSG5bS1m0SHuHXgpZLw7R5FxBjHvGqbXEb/Yo038TPvK7plvtf/q6GN
iyzSEFXcLjD5PgLkvVikgfBUksF3yn30qgd+bFVLNfF49wcG0LzYoiRvAUFPaLdYpOq1COnm1VnE
5Je5ZRg2hXYlNIaTMq1o9cv9jB2mKXaT+8sShwA+FYKPYX0AKa1PJPjCKnQNs7VAE/b/WvB/6N4q
JEmSIvajdNn9XBW+Lnt33s5/jFzcMGXJMw4yqGzp7rUTqBHRql/DCyNnTTl1K1Hbv9hPgCddYydO
R0z3FlBcDWZmM1aF7fsuEQt8kWDqodGqQysvfJ/TexrWoXlXkCNWmHD8cwm3go9RqK7NAupr0n5F
S3YhE0yn1exkupKXBK+H8hDqeqmP/W4snRbd4yeufzT/J+csEw4gbpJ3905cW9QnU3O1KsNHmQB9
bXr7F3ypPmv7Grp/n87fBs8WFQPfT4lHVN5u/yP/h2nyJiBrPtfffJCFhnu5E3bXHORlnR2Rsaug
ADFQkO+VLddKlWphGumTQDkZYplI8FsygTpTvGFQ33gdbpqbYZg3MuoWmERQyjAs3aiBm5dhLMgN
UBLsfS9m4GTSkkGSAVhxjGkpkiC0E68TUTf0Q3gned+91yn48VykQvin0o1ST7VHOL1XjzQ0dnH8
bqroT7zxOAGiiCNePtoHEurKGQzmS8efQqEtvamMd1Th6EiXYe1BaCCzIsD6xdTX8XogOjlzVb+S
cWY+ijJ3BrUrT2zZc8Coqej8y7eHfQNgfuEU0+bpYt0QNc2lmFfAikMwwIJtbCc4A5XvICletuK+
tBMzeh7qmprGdRipthF9qoliqun1MevrzBxCYgYotoQd8Fwv87TSxjQ/sREnFJ2aYJ0AxBfAi7Wh
c7Q26WjfKBGNRaWFAyD4R9XiFyZjvOlvgkUqJoxbk9VXlPWd8iwtp2daB2r05Trd2ZxIiAoMYdMI
aJOVJY8hd62h0do2AaPMz0MeEoaOY1gh/QgFcHXdVGUbdKthu86EMK58Qvezfk/DTlucB48Hbp/M
AkVL//1Bi6Q3XxRnuiBuKlqHXeASObO9psLV2065ufcr0cflKU/NeUirWTxJyGn9r/4/WnEXRvf7
Yuuct34N4GxctAOsN+91Y4mEFFstFXPapeO48oDxm0/JNjamBi3bly8hSmo8+RvTLRTv9sTTEqgd
0xkOjKtYj6Cq2CftBSf+r+eBNZCfRh+GBPJL2NX5M//jA9iq9BNB+ZKcqbbvOQT4aHyU4SNIfRHY
D48JtB/WKVirBa0PeDN+exi51WnPRQVMlNyr2ywSUljp/LZO8OLrmDxIT+rMHuZMGEc6RrHsNoCv
/a+DVxt1AdKpFisIFQUmalzWcP5BZhVXyKrt/WHbjsdzW7TQAJP+68BL+5gvXgBbprUG5+/mpRKT
6keprM/DqB8OAZ4f4OuPU8LlExweX5tTLlbs7FYSZp0hcFhWHQ5epOxFtwER6hEAfCxByjraXui6
nhx1ZMI26qGnLFhhns111UOqV8xlzoYa5/hf3c0GEUG6I+9PV8T7xKfKUZKy8Fq+lYF52XJ7yTck
Hh5ZWbu+nt1qBsvVL/KsrsISTsX+jhjR6RRBel4W0H/NYk06s9J3bDa0FNj2Ieu4sC134AbET0El
RoJ6Jvo+SH2KIQihQxwnTikvsKBZEi90pcN78UP1lwonxUIcPwPOcb6oIGDlSOslgqIh+Q0a6hBP
bgUwYsBOsGUsA0LQusjMvpcjwLPEmpVCtUEmjzNHZxEOQp6oGEcrL/BNhe9Yxa4TlcTQsLBh0RLH
2oahX/A8+WuxV6sIuTaamqTrHL1mCue/3707fb/B8VLJ6Ejru3yW7RVN/5aqRlQqUjDtMobcWLok
5HeiINC9srMpXYKQf6cmMxOHvWxcLhZWG99BYx00BGxSnE+Jud0KPVeBP4FjTcXhw12FjjYvRuvv
k4R/earnTI2uNiG6hHCAualtKZjmMWd+C+HV6eoJkRjuFtOF9ncf1UyOeZPMx+lx13Z5k4I/drvX
o761pFwAe4rVIdCdi4G5SvrnIH8ZhdtjMLHS/shg1u+OB+9Xg8pPc3xewnNYQaKHQkqXwAUqxzhZ
VXBU8lHeYdsFf/4zlZLl2ino6721e7QSKXVQxTqSQI5QjDVonUE43mujKJk16kNVMfjg6MRs79kU
Aadk7tQ63/NpeFBW1vy/BwYnx8BAEN1I0WzDDEpy7yekoYRW320vBpU2LcLTejjT93RoZocQZkVE
8NyCS4jG+vQzQANKg4GfmCfukBmWjEcbcPoVY/NcFff5eW4xPyTP08k5AvCeNjS0qaODB4Bn3RsL
tMGXwjp1wUNRCaq9C0SFPfzY9c7neG/xUpqW4anHvdotAhmFIWtDiiYlCrzDgRmQvN7CtnAaSQQ4
5FQJM1KKCTtAyKXm0RYECJtH7VlgB8zE4lTPqLipjQtRuS9nEELSCRzFDgr/0lqM7QWuMayhtNex
pTVYY/0VwjXfMvDfs6CFi5/uUqhcxI0lcxu3R/6/Ml6D+h+3XVaZE8B9sW7vqXqLAwFpNDif2xhy
5WOWaz/QmveOZJa6El2nwEX8oF2ibp1yHOToTAj5Fms4YdHKSVP1GAf3gQEceZyRaUR5J7rCyKWG
KTb+565Z5V7D1lF7ZJrsETA7M2smvhgM1Y5f2Id7R4Sr49pKh3hm4eq6G6p+RrV6tJw3jKjhmaLO
R9DR99g5WXLRO5baa8zt2sVxg3dVlPf/xJfk4spPSTVoYkzArPD7OTGb9D7KOuGykySJWoxqSOY8
d8d56PElz179tbMoTPlxzID4iiZcP9zzSgaWGM9u3iofdYVIfw5T116A9LZ5AbbmUhCufO3gNadm
JAjI5QOFOFfNhzoIX/Q9U37o3RgtjRIOFG4EN4B+sRcn8l5UNLrn8jANQjz8kYAqRpqXD5h5j2kC
xXpbWCPw7vnPD6VrZheC0GgDQITpz0zIXZBGwI72YC8NL8Oy18QzF7Q9Sk1qlh+9Owsa6WBSsVDQ
TNAPojwwB4meH5Y36dTb/eLY0Kw30N945rCdhx17G4p0DuW+p3AWabyTQgKcZkKmWYi35s+6cxgC
dvApCr8NbMH8xomsweWPjg5hRocwR06gwVv5peGCQ/mwsOTlGNxx7N8zEDEi+nCnkUfltgG0KplP
BZrrYXfz40BBH6dsRqqh4915t13s8wm8Bq8W8BYV/0z69QPywdYUiR9/AlceKDTp6+tm9qWzSODg
fXejBigVFswADr9YAU1V2qKwY2Lsfz6pAWmBpQGvd4B+J5yHKyK4XwNQBHzKFT74h2FtCDc2XOX8
UmvLdCrY8MnaHMn+2SkWuQ8OWOkNTaPkK1gZ/pVfylpy/XUJZcv+l8AAm9Vnk3vbm/G/imUI2XMg
OLsdcJUWbBTVCvFM1jCoclknoN3ptJgmJTDvA5BmBl6YQmkL78KRCeLksx/0A9VabLquisvZop1h
Cw6a4KB0GUwAFX7S8qv4nfDJIAgSvFfD7vL5FhsOQq/1rmp/HCPdT3BgmmnVyKRBUvMmB/3Hb+5x
b8UwUY2gmNvki9btTP3jPLBKabzp5QawNi5S+b7HT+t70n03ButZ59cFpWGhY0pgRqxT5wLUI2ZM
gDZ6L1QitvepNn+hUswBUw36UuBShX8NUZ5jbpw/JaxUrB1GyvYYzPUfathsapyJdE8wb1Nazx8k
nuPycWWy/OZAiWmBGCPbT42RCFLkCVtmCTibeEpRhuX/IL3+m/YCD1/zlt88+cXZDhCM1FhQDmmB
1YwLTNtxXNo0eInXYDOt3mTcg6RqT3hfYuPjRzSDcJ4QXZ22XKD5hvlCnlQSSK6nBLQfx7t50vJo
ya2nZVWd0On/p+MtnNu5OOSfOhBmu0q+NI7iyGSokf+kTSxmaHLfhf5BZWYdIhYCHsq1jWhpqdru
IsPX2X/fvbj1C2WHChCF/93jRCTRaZEOIsmYJGefA/FKYLDJuzNQT2GpzUj+4k808Tfe6zI5ctUE
xOAhoAU1bJDtobFRqEJ1UEj1CkSzjGR9Eya1lNhhKzgXGmPniiBzo4lejMlULHH6joquQxrhp19s
lCSuk+IogB0vXXoeGDCnXzO8Xzk6LatlphgDtl0eai595BmNU82wAf/HfNN6/5aXqJS0IG/z/ja8
ct0XJE65lC4sh34ydBOtdUbJXGmg3QgUhGAnixb0EgDP1adSvS9hFaSulFNZ55go5gy+K95wcK1a
R/X4M6UL6PO/9tPgeXujJknPPZf+v7+rc/fnYndXcIsstR+ak9YTqrskiLN7FmRx/8VkQGuXgZ4/
9ttgAFtROB7SVCoSZkRIrd831xSKcqiDtkNjB+GoRfq+lu3pR8bja3/E/oUO2K+Wem8iIJ2loMAi
4HKWLjeVxh/DKKEbptJnBj7UZguVwH5zZr3CcAIADFhWO8XcNk8adgpClnfzqhN6XP2fhrwMOJqs
0Z7/G+hBB9esAJqAzMTxKamVNzAGp5xz320mnt+U0qXsbSL2NDckIXENuK8mn27VSTvtRBN1uRKF
ZossEz9n/WlwTlvYzhv4Rw3GAdaEv1dO1JOY/FGQ2pyXlgKEJcLpz/5v30QupYUSNhRfBHOfXEev
ALD1kejW5SSeO+BaQ8wz04HR7cw+UizAwWhsaGxWxteL9SnSYhmR3nCnDGBcVlA7cNnqbME0luk/
OuUYBVgiC3ncrbYanyn+rWmO4ZTInJlRb4gdjUn5WZxEs6McXOZMzawzzyjEOviQHzKg1a1QmEfu
Rw+oauoBHyrP4JXd7JMWfY64/pT1/l9EPi1tHHfCQ7Gp6Wz5MaTHqAJWB8MXl24I+LS/yJbU0s7f
7EwNy/uTWHYhGZK6Xy8qc8YMbiWRxBkIMBelBwC6PI67OFlhsRdBoMLYTCOtaM0AkRSschOSdN+q
C/0khh4xq6tlbKiQtJRPWJodh2pKkmIzEBATyVYhYLcX+I9OndgFEgGfuPUgVGY1KDgQocozHbjZ
U2Al0G6zVcJYBDCLFlIHj5IxZyY0KWLAtc2dN61+x4RnAevNw4sQ+MyLlDAzfCHdGNL4tJip8ire
vz0FflxwX/X1ekpnjjDToTMHa++to0SR6WyufTj9+is7KqdQn9vA900ultCsjujVweSJSuicouAt
e9LIXj2lEM2E1gCKYV0SecWD0KRVkzOiC0bmANRipLs37NEPieKjUk5uYRctNUrAg3y28MpWx1JI
zvIjTsKgfLGEibNm+9v4dSVaMiv+lccP3KesUZkwqoKmL3Zw1NK5PLZ+57DxYvJTms3JluCtm7vG
CVKkGgv8ILxUSI/TM96KnxFR3OSZE8U08aMbuZHUmgIAxB7H0FLnAED7sx7w2ROWR9u1hsqW/CKQ
smYueenSDq31BVK6nnNR85EsB3ffwLF+Lxo61ZH2+VqYAHz7vs9yIuzEhD1/w+C6vThCoHWFVayZ
WdSkHKhXPAz4gw5hFAGxKIeD515UjrisECnT9uNhHR9yg4CxUVGHJplWnGRRdWbWhhadPyBgyfOE
uYEDc3w/TS6MDUhj+r6ZKp//uu9W/x49ZXhZ1UNjYy+aer0K9Pgl5AifKotvscL/E69cURuGkcUK
QNjICba/BUQciADQegXpuiJS3gF3vqlJxpmsiPWj+I7io46UyFROovalW+s4sAuNHrIFtJPV0soc
qt0oGAZ+6SiM5Ai1evH+L+cFrx5K4zG3hZquzsJZgNII4VwX6H3Ta4WeXpjSocVDeAwsqko4BW31
Uamo6AoQhXNWgMvKVtXPB7wPGRCwctHBuNSRkNEcjLVFcIcn2VsjnSDiPaQXLXeoMpBp5ZgN22XA
caZiPSyxLZuT2/L8Bf1aEwwx6AofMxfs8xoOZgfMa3nybgtkJ7MSV3MEpW69Jpt/25ZKrTi4XCBv
9nN4BX2M0l5vGwXiv/KL9SC+SJ7y3q0tPXCCcjI1WRGQiqzqaMGO1KCudAKqWvhdAwOFm+jmB3Iv
znk6GCz4KUCx9qbrfkwd/tGEZuhL3qw0nang+xK6qk/uxk/MwjXn4uNl47ZBmtzGd15EOpJtM/a4
tQ1SY3OaiG4OjwzhaT9RRueGD4kq/JueEDV/6FfO1BEBG842SEmWGRk8OAA1V+1pSNY/D6u8GT5V
p+ogtP36VIGRpFuhOKEfyOvHjPeTMlozmE1/WBnykjy9FZ6XuH/YwVq/vSdGE7WJ9ZG1Eqdq9rQt
OGov8FnDEcBjSdWs1CxATfc9xyCZYCX1lY8OpYFpJQIBmLDq+ufVXAYOIT+PawNa1/z9+hQNqD5G
RYkvJPfeA9NkBPjHrxk7j0pf2mCz6WujDPWdCKgVZydoKxdfDSEscHxC4qoR2b2lS3fin0AqLKpO
nK/fJLBmv/x9bHA1uXWc8DP/AdIqtX7+tcSn2MzvxwGSgRVVe/GKqjkuSWWAed1C7aGy//dX4esv
/8cJcmfd3qqACKw4adbY9rfBpRWHTqnylx/1OZX/xW/J9Zb73k1jqy3LrzjL703NFpPhpWduGtWl
DWX0Ct4owsbk60DlWpxf7XJLalJJDd9SvG4iEvRTGODkPbEoGBK8WYauUvmh//LYPYaAWMvzl/gL
/DaT00yWM2VJw9rfbA6j7fv2pvX25mt0XBe3bcXwLHhUBEAKRZFgjw0SMYhmBIqwdmVtuCVIBhx1
iEvZA39fMhKTW6ixwLIwcSI+GhJp5DykLO6YimKmcLne+pfssqUIg0bZDCgUxOZ9KkqBm0E4xZpA
xUDqyIG+iTl/Ozdx4CIGNfOaH6DjbwbtbWpXElwg7pruJE6cKJDV1BagHunImDNyylsvDna22rGB
ai+kvOOQwlosRMQPjl8i4+jwt+HQfGQKFAJvnqjk4w0wocddwsKUhrvt0ImdwwmAd6fTxiq6/lWF
b0yD1Kq11OqZrbizNzo37sX1IH558983ISDuXSI9kb7v1GK/kemqlH6TWrmf5JhS5OAkHk1nl89q
djy020j+oKzqHyaa3NsCcgiOlrsRzqcJdYEXZrPmszav50CuYouLdnZjXiP4PDBQ/a+mAeTL+O89
SR2ZQfp5Vr/3LeZgMkZ6ZV6CuyBTuVpqvRAlZWEi8xKxrFsQJ16eFQWXgvnX8NdzvWC1Inz9jA8f
kM9tzTW+htPqxthEiChZbcWLAG/mRfm/f3cJX/ehynQVsej1cvr3cqyD2WkFKLwxqZ4jfupPikmv
6A6FpT6fXs+FrrbXu/lZH1nMMBD8qpJ35c14kT5ve2XBHwiMCp8LSprpibWovAB8eMEmxPSbEWEC
7IQl3ODAkdg8gDvdN6a+BmaJ9DcrqQ5qAWNEtNS+0YQU3mQ8ugfv8hAciBdAKrjzF9A4WlRGWi4v
hE1mV8jAjH2Nr3zlnFpk51cKv8TAvKqEAqWo+fJiCc2ZZR/rTJcKxNhk6QYDFSq+ZSvBhYEJru9s
5GNwswuyyNiheDjWoFNa4wCpDTHTorvko82YTCo5hcSP/wUZ7Q4j5xJVRizg7AcZe/26kTXftwtn
StCON/Wo+LLxytT32nsUneMha9wMYZ65i7A5/l3nb5tU7IuLBuzvhlU2vKCDP6KEWtmzzazSZ1NR
54dKa22334Dry+vIdgThgNWt/7AU2yR7x7xzewwP/gxKC674OYbFWOJRltgf6C9/GuK1ImKptbEm
uwI7GdCw5KtuiAvEC19T2266Np2oDE3sMp+zukzjSvwxuU5il3bM9GpYwAXq02HQb6ESrp2P1mEP
19tQYZjqH0eXd6wt3FU+kZ08b8SbHZCdlJDaKo62pCGaPfDMX3euKjrRiXekmqBRFJwtaqYDBiIe
dnxDv6knDFd9Cs7hGr9YipqVSSt7XNjrvxQp5zSpjcZKxPBU4YCN2V5QgF6GXhRS5bQugtlCJMyc
dS0YOfqhMixuWGlj4sjLFPOtWrWxY91pyzI+I7srssASElXn3yPuLRNt7wURtNjO3MwuFZbxEbR+
WaT0Uqe8yxc7b2Qz2+7xjbI2E9mwRyUHEO8xjAcJ5a6g3M6rtqfX34jHureX5wLlTEnRPFOXz6zY
ysTzf56M9WQ+oisY+CyO2L6dzWZD6J/7Lfh4mbYNFVpSbVYxGWvqU5/eyvwfZp6cZNaOxtm2EvsD
QH9KUo5KSfZJWowRHjfizOVJMTpCOT1LNd2eLZOsVL3UHb1pHAw26RgBH6Ib9PdQ56+RcpPn1mdn
RcBGudZlvHYcEGqtodEvvcOQYeokZ4W4tf5YhBB0VXv6v0uMlWGrgGsfWQN6hHTYfzr3gvjSMLvT
0KQfsstse1YIZRhFvenLXiLPhyroycctYJUpeH/BrdI8Cpl1PHGmJoIFJ0SuFTo5GGnzchccuN9R
kSz1KXTD6+7WHJOKxp97BMBvBfaotDGX1LgRCdjP8W5gbIaHqvrUEt4CzVbsZ9h2flPxxqxrqAy2
AI9Q6FTXawAd6aqUrBwO6ddM/BnzXqz5+iudFfma6j2f1av+Y57B3It6NxuARyweOmL+efUlzja9
lM4mdEJY9mXz0bn/Fvu5Z1qMcUsdscw8Q8j5bixCQisrlWWhSMBVwA5MgxKZ+DvSN65d2as6xMxR
EXeW0T3ZrkyGlDr7l9ffPCxBAZoBL6cnq5gvdapJuekRglZp6Qigd5+L8qAxhvmDT/51rI+AnplX
ISk6anQTgS2PmXsFN3Qi/ju5xCwR100QTzHHBY8cNkhrAoo3Xl1Z92C0zbwTqDTdJ+WrIxSzcrge
ZKEawxZt14rLJk2MaoKDJ71P5H4K97mT4lGxbWQlz/kCAOtISh4vdPbPJrsHzAQjGQfMZ1r0m+ho
JDGuzpyeYiEiHmh0k9UlOCVKktvGg1GiMghSFECDQkkFvqTa/2admCqjl9GLEkNhrvfUBm3tNmQn
7FMAQslK8WQh5oLLvDgsCmHKK411S1HKYynQztEKp+IjeTDgMw3bA+veFskqewFZRmdFvqsWkkMu
8LmPBpITBzFhGLitgVjQPoWJdkhFpx7WxGUgQDUGfIteYf3ZTvUqjIFxhbmpgJKawX4OPLSuYETG
7Vt9xatVU45JPL0RF+aeVt52Ht0Ajr23q77XiMfbqyr3aGdepL8Qf56PQ3zVBS+UZCrHWZaqpJxz
crCfsiZzAVmnUVOYl4uhi+YI57UrLx0wb+/lzy65F4w18iCQAD4sXnNRzjxREd9NdIFrdgvslVX2
Zt3Y+R20PGkO/uoBzpo1TZUdKr9AirVe1JPsFxaGAkjGYTNcWkkzAjMkfQVSLIiZ2QPbPCGR/pJa
OyiTzfDQD2ZmCvFMDp4n8AHiU2J24F37J7jfDbcKZc3dp5T8hWX+oF9y0rPB8K46nnLOQgs9GvfX
BkThdXTG+Vy85rO1W+7Bb31TFdjNg6YQGwhqLOxSbpPSTNJFMB96n11nLpDwyEBdw58OoHpXZ8sJ
HtAALSzTajZnKtEyCnRlIFTTkABlI46d6md5zE1vjxijC99pXzCUUc3eAkUVH6RVUIeJlmdX4plZ
sA76H7aYIG7T2jDn6TKJc3llb1V2qnmQ+rtcAsOpxFbF44IH2wIomzPJJL5EICZkFqP42XP7LFUR
Fya6auEJNdIwdFe8KasMnJfHwMUVA6DhK+iRCXYq2lZo7yOGK6Qvp7xTr5kbCwGQX3t3lT7chjNr
5Oo+cYSH0RMi5BROdCeNuV8XGI6GUoLW5dQY+QVxkB/wuTXggtldy23CjJIm24Nie1B9fxZc4RpZ
FfXGVe2dVOqE2G2gcEfm04r04hgDzt6njyLSqTcMo3bU0zSgLBIMLzxs8c+FRucKyFsS3SvV2gXU
Pjmg+zMB1gIMLLBV7rvhls9fV8Btc3o70GY73T7qPbwtu3KBiNbFM8/xfihp08p1PQqMJDZm7Urq
nIdaD8wh+yuOo3GbdhBlCf/qTLlT7Q05iZsxlv8R+f/ytNKIa9DHn7wIyLdgzRtR+1qpK8J4yMef
3/geyyD8i/HKbXJVH0p4GZwzFMR1R0ARNqz2WOGzrrqAi9JrJhlIH2Q6tKSQY1Y2Hke3k14IKb2l
kQmR2oF/Wm5wNW/WJgqlwEdmozz6qS0O08VWHBGzCm5ja37pm4XIjBCwti6txT0ol2v4p22J1k7z
4m5bVRENMPx8DkvfSiXj2yd0vhU8YM+khNYnoEnoi+PjzI/uUMamu0MaaCJXQoFN7ns3ZVYMiuMG
tjEfdxxXLm3jCs7GFAO3Txzi9vhOp4tEf6sHi9Guq/zah190UCNHJcYkP8Y9C39eQRwJEZPO5xz7
mtTNxd6ANqlMKK7QaFZ998Ys+fIUyYq3WaSatKLOTOBwW8bFpRyy6XLMsIsakrxaKRZ2C4tDKecl
tUgiQwoFdcXEX1qglpzhtZzC5e6K2Z6gyBWG5bwxJGTcl7BF54zx7gDEg6+YJS8ElbhcNzpApkAF
ivkB1R8wSX0dCImeN2Fj+hSGKFxIMuhpZudaO8oLBlCSmkAr7d7QL2u6wymlRIyAsYX7LGm7YioF
VXIOUpS0LHlCuk+kFCaRASYJYD8aY0ONMZuHniHqS31wxgf3d3GRiwh1o4VSRKX8epMqbZ2QUetD
+jKcLAoXiEebpbHd1tJN4biuwfP5Zy9IeVyltpQtxWbSMNVTfZ2bwt8zyZziTpL/Iy/r00rW5fAl
790j8Qh2IGRE1E8eek/pNwZK/xLZcSQHTC5PqS3G/0ed+FgiXbRz0FSQ6eUjGugtWXtOaqv0dY0g
iz5R0mjHsf9HOc3GzIB2KydCq2IO+4vi5F7ZbRVz5Lt4tcH8hF0TAOyhRxV6Z994l0vW6GFAstQx
G/S+0x9X6/Fm8DF0Vr7C3oElXdfOtAbwN2V0tLjyzOTfhUnJAy7Xj8ihLSjqMGfqroqokdbLBBns
e4edZIush1mAhA3tjEd4XCV7qf12U8Cik+gdjOuSgZD21lt7bYerNOdraScvwZeXPWQg43xXqOis
nTGHiYt2rEUNrinAGJvMo+lEmD+zfOsuFrGZnugs09PlqVCQzh1oX3MlrZSErmXJ1icxgGYDgxsC
cjqwLCtNq7t+BeXMso8PtJ9QQOehEdOM5bSdAl2wlELC5RQ2a+XSrbYvDR1tKAaKj9b/OcXtIFM1
X3Dhr/66rJ3H3KEfXX4yUoqBMm+AYXqV3WLzrTe5g/suHKILz0ErfU0dOYcjDZclf/3wOgUjqQxe
hl9gpV1vzQX7ln3/fZfFUxtYJX1vIRUIoijNYg3/xc515QKUShM2ISyiwDnLBMG2ajUiWJkjf5S7
Tx2moMdjM0xSRgLHGOWkcF9U47mUfFBh1HyzBAbDmtUznNIMUyLirhNsWSZOtWwDoWm5fEYE4VzZ
ZVFerEmRdhhBkE4yBX8U5JN0lFSUOsX3GNGQI2qoUkLSlXX6euTIu1cdzWobfmsSGj96KVxA1FnV
P1P97VqNTUnnmj99pSwoHqdkg+KEchXsV0k8dh4yaR7pVY/830it8mDxiiAWTiKokbwsBB1BCTco
M0D79GLity5DbnlcrIs9y3qXsbtw4H1FY46co/prxMnm7j226eBkZs/wAKz7bgVXvA8f3cKuSB/H
uhHdbEcUnL6qnzfa14xQPmKk7u5Ti27+Bb1ouLo7rQy7VVK57fxfNYlqlMj4uLps6C0+RXWq13kq
ONVueN2YnxcdfeBUgpPLxTFURI1+mE1FinUdOB6+6PryztmZbTF1S1HYKvcwS3PL8ibqKyAuWeVM
hXIjrqT7KGeG1R9/hIvb2fe1I2ND4EqockNxiwhZluj8eETkPvN9j9Mp352oEPrWLJtwoJlMDhGr
ZAw3TSR4f7Mrj5WBJqmIi3glY1kGs4yQ+EIkTaDpKFel9gp1Jsgr5XoFPi3pm8fG+eOGmb9Xkrwk
9QjXGZ/SJyysBRLFSSwxMYOmRBZB1g1ZKgnvKtBoz8iiSJOjqt1WN8jmbDy6NUoT53HHdsrHxqcL
u9843s76l43fo/shqcnYspUyqKhu+IS87dmU3eyLxkJmqWU3qA6gOd4nIXo4Sm1dIFJzqlSFuk0q
Vx083C61b73KvGIoGwEveSycBDC/50eHN+3e1vLquUUxuLb3/K+6Shf1VhUdSG3ZcJNtYkLURQaE
6HNyYfQz0SI/48FtPhv8TsdBq1NzmmksF6szteFQV+yf6cqiGm4yUaeHYQRRXtIFQz6xgukrVg4K
H9DUBMFau24/YNSt6ON8hrNyH/74gF/h+YnMal3N7OzUO1rPq5ew6FZWDzjYvljMsRYn1F/oEv4C
99SsrWNvnofWt3z1QKW5M5AJPyfXPwlnj72/oVMX/rK45nO6RbnICdsZaatd1Dkz5Ha9Ez0Bbbve
SQsYs/haA3oYXRQN1uIfoKuFf/0KZSuqiKYRJxDgIyg0xhMUgbBA9wrBdbXznGhGLoIZkExRVRok
NvJSs9o92+q0Yyh16ukmGtDpBQIt6EWGzyZJpvBmlGTVyl/JbryLv40VzDYVAyVQGVFQyrxJZNXM
WLx6NsRfTjYZTGqj6z/rp5s0lVyPWHqTEUxjeh+iPhaBOmSdqp5c//cKJ4+AhxXys4sPKthMfPTt
aXFefdSKHttHADXE+SBCSOTvP04VSMrNuCq3mXgQ6ZlfXv494Hg9Kyd4a+nD2b6uR6WIR4SUp/T/
+s2C2F67ECrJ3oiqO2G+dWDNU2rW+g1XSoUCWdue+kBkR3fad+oyAZAmZ2ui6DFIgzId7/zsFiHe
Q8zFfM9Vk5osc3AC/5cvqQ7r8bj1V35B6ah6cxsB90tHZfbo3a+AHzAF5Xkc0aBIqkOR/nD7goCg
u0v7yFmijLjeav6Esu8HIgb8lys+Yur98+ynpcbrGpzxgONW2jxmDjV64xiYBlzfrZA46x+5egkt
QG9/GF32jT+tzmGsq5PtYxG1R0niqUQYsV2tWKrZOT5wK+YcYgenkuqP9k1rhCjq+v5qfXtJqaog
78n6SL+t25nAow/J/P68ubgtsk282tG7i3sQVp6OGU376vqZt/KODDNN/MpXgFfKIsJSFeJ9EZiP
27yZClv6JgEXPBi+FpDw82a/kgcEYQaZyh5PzSdHXhv954tO6uyegJa8vnFn0ts0oyqPykq/GGFk
VhHppKmoGUHKn5a8ZTOkLylkTqqkiDqqbzOiXR6Uv66YiwP+7VdALeZnc2Whh2AC8ssSV8WJfge9
JbA8q0/DwFOKJxOnwfN6p81/lJHPNt9vtrV6lL3Nc6djD7KCi9gw4r8kEXdthxUUElgg5RrHDB93
lsVp998MsOLJ03oy5lwWjkBWg7YTKxoz5jRuzZRL6+Dq7fTdr9M1yQDhS2h4Vyq2nrfj8OAL0Cm4
Cr1YXQInR5bHKkIyPiH4FhEviRyFpEOK8uVECXyQ5ifpN615WcMtXOHOqL1NTfA8fBLJOXgD1S5Q
uEwKP9tC1kc7dBISfhhC9pWnRC/AktjlxkwFXDeJWKgOWCf2WzX8Le0+urpme/QZGhKw8RTf83qi
+45SGVH9K67cJGgv4UnsG1ApFA5C0bNGUNX8z5vNxMFZ61OLNLAgcSvs0O09UZbjS4x/uZQA/Sl4
pRIrQ834IhWxT3pMtwmfIJR8UBLeYqAZGvHg5utG6Ri8ui5PvecRa/VqKtke+fzKFyECtYeHzt4/
VEtXXIDgMDQnn6HLds925l6fcUykoXJrUSzK17qHry5eCjnEVascu4DTGHWnOdT4HeVy2WO9wRpa
VblJ3b+TO7ZxX4qL5GVcFL+GLkpMhKy0p1FkXfmj0Qo88zLGXuRT5mc+/xEn9FSPUzfMHveiK+LB
Bh8rp9f7R6lJgYLfNI8s1TW2uoLDXph/FVVUZiJ60RtvSqtHFNnB1noFpjRVJpJw7K6QvVx8zvmc
6cC1C50+jhNFpgWLYqYkUQbhKMwBLKNU90Q7AHGHO1B6S8nQ2dY/H868wFswC4RcF284p1Rf9PkG
JcgZVdTnDbE/FVuZQ7FpzHikg27nz93MQhN0GDuaQ+Jy9LSTkUNvVmV6qFI2m+ui5RF+A1znEk2O
lelSgkEu+a6CA6nZ1nmJO0XWrVlUR/dCvkWhDxkRr5SyXuRZ2GrrHEj+MEcbHOzppFmeOVWeISac
flQoliVK+gySjjrlLT1vHEsK3wtjbhxLvkn3YChkEYE1Un+YwoqIlNJBPC9w83DYfyq3elyc4m4X
vZIMLkun0SrVHz3m8C8gOEEGMSVJDrReXpnhKxSplY/mYhsGT2ltDjV8Y77gflrOstBbBti/9n/N
0qMNP2JnLkRMvuJmgmbDy/u7bQ8d8jIV7Iwe/klfESHtPlTBjE8zAlOtXspwYuK0g/ssPsEEvQ7Q
7wC5y2VQ8+GUjgMQ9+XuEeeUQq0JNhN5DGaZ+CuE7X/cRY9Us2Wp9yK654sqIiaaxK37df8TZSRd
glmTK3x5c9aQIB/C468Islb7DFaP/BB96x2GcjV9Kc97OPkiHgN8oQyrk8CJSZE4VXTxsX1MRNF6
HCnDRIL8p9B3PpPNQQOU5GKjogVVZ9ZCxZYQHLFCP80zE4QBRJjzwrQYS/2PfTVUsY3eA3AWsioa
gq5aSiqqD8/eISg2zc8eblWt9xToiPKj1Gaid7TBjxh+tbCzqs120jcNbXzx8f2LfZm4hIqibveV
qkT/fBeE86ZVwq3CIF06b8daVTld1zXiM6bwg+PxppNaWL5G6hFCqJSanHlR26svIZx9CWDCtyN3
uvRUm/AWNxs66M4xSI9dfq8LONXLlCWLGKBg8vr0Zrv3ukXEjxuR7RqMfT/5bq2y5da3PLA7JiDo
C7Mmk2EmRVaDoyyIliCmYZPg5dfpXEKL4wEP7MGyMgG8aMmCOPv4vExY6Y0QifH705wGdRTypEp6
1RUuDVNkk0+K0AwpXoZFm5qL2zHH5mosv/f/yOAIpMGP9rfD3wKcPsLvMMiWxFyfWFpeCKelc0Hc
lFlxyWymS4MIomKMPpYOxP807ybv40gEZkTMfB5G2Ui+ATts/Syow/CnIe0sZrCOVUNj0kgJeTJm
RYgn8Br/J7VF4dWOIJsgX0ns4FUCvfo53GoijuB0Xn1suraZwyh9tx/dthd4wIuZ+raR8w3wDxrU
7+bYN5F9ZJK40pyE21LpHoF+kiHlzCZ+XTO3eah8wX3HjxXTONCh8eeNMltLlkV04skVcWrHEsPo
RJTO64pgfqZaCkokqUQhAjGTahpGBEVLHHr7+DCncJQ0ZSZhIQ1YJ00DqZghFaFk4GC7sXuVNmxD
9NgrPC1WdbTSjFRHw+1BFlpbGOtfUpIMPeQJrwCZ/M4EOvS/1GgDyb0pYFfSOHXYM26PemvHBSyu
U6RIbJIf929psy1eedobncOw7cScHK1XCQQmUfPtX15gV6hRkmtIu35h9ld9/s3qsk8GdVc3ZG6f
6dcxnGDt+P1k0v2G03AODqS1Wy/T2Ji1fVSqJzNXdoCRID0WgCd9ksh4cmk1xYheIr/Pq1z6IeHZ
KGadk5DxqwUsarsvdP61zEM18yrmS0QS179dRZXxkAoLxMjbWb9NZdZM696REG69+SFLwHivR+o6
ATe0n//254MCI86kmH2d9641xHnfheioJXdt2mLKNGJKmi3Fluajzuu1HEhBzctk3VOilSIArqn9
1whzFXFE0FGZvFa76m/ua8Xlh8awsK1+WOExAycrcSlZhJXPZhdnS1HtdNkSy1PUiFQMFqDaEsOo
Gz+n0ofiWPG9yhWLjxxVh/PxHVH+bR2oHcyrY/H+a2i0o3K4Qk6Zb1zShnOA2LTEV6A7hVngfoET
/F96O+0OGf5nGXMWcK1m+ro2E1cICBTcaY8SXPMnbI9NVq61bW7//FcYEtCvvV+rIhnHdo38QSBo
9+fN43axu2gcKzParEFxOLc7L8kEbaCqP6jbHA6+nABjtMs25YlyfEr65ggCw4DRRz+BLdZC2K1o
Ad9+6R8RPo1U4GP8YSzPVMum/3jCQTmbV9MeeJ3WJRgiXmIEvB2Fn/veSkKL3TE/jwCqCbkDiWjR
KoI39TY4v1EcMf7T2ocxTDi15cUAsYD5ge/mvsmJCzTCoVLPrdP+X8f3hLfmdHmrOtwBshp2YfoN
esSFkg6VHyJ+c7Vm1t87zw74zLEMzTRgszEze2AekHYgxMuYBpNhS+hgHARYhs8LlVYHP+DT7TmI
6+fy736lPkLJDXhdP/2AxNKr0MI4RFZmqSh3maqQWhJZvxvXDfaRdBOcz8kABMniSKnPxZW7GgZw
UPK7zVSVhApN85sLVytxGGP+WDo+FEFcx5P6bHD7RP5Voje07E0IrtM02Zef94eSjLAaZ3bwTP2W
MxXCzHTVxwh3t/98pavT2L1iIxHjtLZ/Dik1I9O5oo7l4yhQ/2A0oq1QmdFgUEH4srBZkzhq98Ex
CVCDam9w2s364tL1hdpehvLfU1D6rDD0oxVPQMSlwZ+EOwmlviYA6kd3jW2nemJMR7XyOPV/cGG0
6mxVbfThQD0HV5Ne5XBBE5cXbLgvqpZMnClPgwX+Cj0F18ENNgz9ZesTKSMnIq9puqmTLKS8EVmU
Ikdk9ZAXYO0ZAIhJZdtluIIlx0N6YS9Z8KubHJ5lGetYK46+dZEpOqaqdtCSJ6GAZkpzCRoJGfLg
VEwEF4hwcYPEgL+PfK217Ia6SgmA9doCF9ONVlVZMOkRyf3bXXsadwny2WqG14lCRUnXURfeir67
humibWVqG0dKNoSJSexSmaaHm73reAnjjMD9EjIy4tSm3HUgq93BYfzDkaLEQnNI1NTw27/X4vQg
yNihQ7K30+8KTvct+Q9zxHEa/DoQl7Lr1FZsomxskcLhcV9AZ1HXyQNdCyS04P3m+1MTUg+DphGF
ic+mq4fFRJLPFq/jVZlKPS0eg1+E/fIPFQdazAf0SNksNAuOXupOSnNbZknBM7aweY1W3EJKZit2
cWWkGbgbJqMytCUcaS5NzuB31jY9pOfqd3P93nltAM70PhJrTqkx4se5tpTg1Gy/1xhHRgayERYV
6a8XGCVMaxz0buZAlgmG0skQtbJpOQNdEOxMjPs/jIONVJTdC9k0s2Cu0Tw52ItLfr5igU8/lfoP
TyWk4jdM/aZLvRc5R8v6xL2q/AsFiq2PPbCzeFLlVwGZbIycdWnQZcRRH1ByQaOV0e91wrI4B1d3
eYDIsC++sgNQ/9Qfw1ORoAyp0/Iu6PNfBUD9S0/j8yxXjjkCS4i/AgjBFwdPmctY+p82sQBa9OC4
lepDbB3UpIKz1AtwJUt6b06Dwrk5uptR1ySSwpdtl7odk+wTWo6IqslFxry9tGPNYNLcGhoM+yYN
N7SvO6J196Onqymo0GIXuzsThu/ZPh63mwz7wnrHHreuhxOWbz1vzyRnGETK1r5mVCKnmZRWhUbw
T6szwyfLgBWE3ekbDS6Jw8CH2Gj+vo1b2ZNh9xDcuDGKisWAWh6kmm5AZIvkK2mVbcc6u2Dr3He2
NNPS6rQU82oWX1FIOSJ/svSNycJfuk6He5j3f5teFYLB1q/pEMoeCpbdFFvMc1rdeUGRY422aXuy
F7y29VQCeFGmO3IzImNsRyIfb+4GC87UD71Rge+zP261E+8yj1esCrDmWvWFKqwAOxN4hDpfiscf
FmVfelhxyk7u4kdO18nur/GGO4eKXSyccV7NwpJFkcJPsvrVnwwyM8KKaEH5kBoSaEbr+lN6xlq6
PiwgxqYWOPpGIcIxDJ+EhJl2XWNxZnWWejmnutgmLutQs3zPJ2KyTi1SvVqEI3t16PWfKfRV5MbX
zoGmW2HGzKdYdNqhyWzZMrxTaaGVkvbLiSkjobOE/amvp5hj8gUYwm6rGZApvKM/Nm5/e1VKKWw1
DhTpdFz5QEyX3wyPBD988rBCWF6pPrUBfmu8Af3jzjb+lGERlUqgg13F/p6u6wQld5oFNsn2JyXc
abyy4cjK+1QUxoy+FYMFdF4A3makAROot5jXNH2cZ9is0JftVTTxuwiYHjXNHZVXPPAXFltr06yR
9+7aNjwpMfqUUm/qhM2RHozft7P3/QDzqFN5ynGsdK4bNSrezi5rL/YAshKaWgBLET+oy0zNb+qY
p3FjACUKgWlkKl6ypzu0vBWw0stPQnI+bDZvzhyJQz0i+akKaZ6TyCIHCwhwxWKxOcrUtdRs3KZE
lJWKv1+Zk7pIWjLHWrGXBnuWRTvRI9IKRNXJqgMWvayB2zFXXmnSL0IuKMbw3oRyplZUqaNn+5oe
cWsh8y3ZV0Fx48Jw3VODejOLkIohtGXINDaQZuyn5RSglOiPViWKcTw+2J0pSgGoljt4w5qs8lhf
gcc24maPDfbS65PA07IQHsvt+h6ZV2zuN/Sb0uMP75C2VPVgpo6LUZ+tEfqGgRDuNLHLMEPDfdVJ
oM+8UrVbYV/UJWJ9q+XKY0ceOo0EqJ3yWineD8ElL+TEhLHH2JHRe28+MaGxkfkV+hqAk/cy27xY
OduqWgKaFREwERYpyqmqGt12OHuJBAQbuOFV/YVJBSdq0O/vApyEHXnr0Zhh8uyH9Ho19Iu13ajJ
OH7V8Rd7DGlLGUqxHyWWCB1AyVLxRhajR9dCZ7Btl98pPirWrq5eGvu4FOr3aM9sMvBTrR/Lo5me
JX8BwfsUvdQvy2R6WU/HY5mmIhl4LxxmOhpIxGYGPH3bFTkKDyvUUlnqAHof7drrowUgBZWs8iM/
TJcaDLs1EYiib/42bhAZLVf6sTZ6b0r0nMpChPeiirvzeVngY16ZPyIs6dYQgl1ssuVDBkr7IgI4
lBZ/cb6dJkDUdnHBVvzxXKc+LMLtZ9IkYNa0I7sS1E7civcBF/HuUrJRGjlh4InXaA5oywkWC0qg
sqkgX29tLc89VMNBTI7W5oacYW55CWkpxJyHeDEy63dWNrJVkl6jLhj2+8es2Xar4Cv/jjkUvRz+
rYEVwBSDAQw+/9kXZW691mRmFMgWJIcYMhosGUm3ubekhGLkKrj69E0pdMdgBLh/pLQpSvGZDYOe
7rFN4nc1ayXHpXVdpEOm0bfYwVdKM0SArsKPtxwv8nqXohDJuKPZEYYAWJSY3CDxEiNs0We6fD7g
6AXxNHiPlMAH5Py2ujmkNz09GL7W8ICBMl64DVdkoqNARGp/+TS9i8sayqN7UFsbrgcWmWcO17i8
i41TUOjKW2xJ3aM+dPdSCtdYHfvR4mo2+vD7h49aQUy987Qcz18CKWeHEfhYafcJjlq830oa+SFU
B0X3zcZMicA4Ti8s6GD4QWMR9qjoI3rV3wwKN7Wix+OSzt2pFcj2hfQEcGYrQY7mybNt5/SUAD7P
IkqdZs4tsLii0ccm+QlGFIild0720g9KpJYZtVXdnnG9Oln21CGKZFWg7IN4hDbFkesXOHRIeNkd
KiKS6SH6s6C2JepUnydwPSiRKrvy9GW9Tx8YXCMjeNiZl2PbMTqNd25afy8LZD2YAb9nGIZed1k8
Sq7ZV1HNGIS98AgUfxP/gVHHdyLrwvzvU0+4bYVHKgGlbs+yeg2unyRMV7dL9Q73gK3hFg6XMvql
8lBx1L0n2g5K07mrpq2McdD7QOOkt7owaKa6aDowIEvuQ534rNyIn+42qkR3tZkbRPAu5+054E8h
Eok7iyKzpLoQkecwwwX0QJQl5tW89S+jQM4wMAuyXqOqyA9ykfDDe3FzrxZqvSDr0iKaFfL2hTox
ldVuX6Qdma5Gbf00eNzvKCWjUTulOl7vnjh/miRt/spfl1Rp6XLdicqSzHFBfDIM863oS+WGHucN
6Lax+9f8ONkIxUUmadWPwSDXH9UW+CIDGpzeO+z278lZxTirQBSDwbA9+uczo5qFTDdLl7H5fpbn
LtAOdw9560GHoidjSs6Vzh8864wxBQsGcojhWMbGhpe46XAtrk+dGI53KTUXSLUdseVse++1qVdZ
IqHemeWsj1bEvXWol/UI851NMpAkKBnU0i4tYv+31jQR/ZtvXphAzIukRolMGxCyhn0Qq/ZlN/Qr
D1d3Myb5mFtdhPHWxiUjwMYEhi1c7y1dYo4ibhKdjhTkhWTiSuOEmMyREFhVNH6jTtFksbAc9Qgs
DQv2pAFVI5wwojXyl3W6N+i9A/5KNQTYdL7Sr/W9yJQTDh1Ti4vEcsqQmJGjtFjgI1bKhUbL06au
qOXxx/LHdwfJu4tbjPks2rB5y5VaPy647ot0eCcWsMcSrVNk6O5rcTAyXdN4QPDiIAfaJfjelBxl
r1Wy5wkeAiLesZv119XASti1Bbd1ADSokU/0YNgViNFXqcZW/ScLTWL8aa4GfeNMvn3Xsg29pdha
yHybosFpWXruYvvKyq3ByXgPDBr+fpIaOds64vMLhGbNIGA+r4+MvLXdDEspMGKpSjPZz+MfKkIJ
3MlfLDenrrKLXVsF6etRancMkx7TLg7XBERGCEs3S1O+ZyR5EGSqaYXe491iAtA+DDTmTBh16OzJ
bZVfgn7QdPPLItbEuIIk/qpd9zJvklpvpKKV46QeTduzz6GBbEWjcRWLDHQoHEH+VJ1gQm6KsQrI
aufO1HRSIC0xM6snXx3a8vRzLec6XYbyqWsL4VhV/FzTOgXytVMEfRhDY/kCEKIaqWfvxjyXQlYO
NH/JjdjfsPpBkbvlaYWf/I+bEqoETNJKZKGs5zE//oNftcl8TEejk7w3D6SSmwwbVfDJgeWcvnxe
Yvel90LNCZeLYqAzSGbPiK5haG0uu6JMLOYX+wD+1Py/RLGxV3tUi9iCeBMH4PBkFtd8WvTGIEZL
A5BuzcCxWoiI+wy/1ETh/XzVdNI/XCtt5sfbZrcFXBBLvipnM/nVAE3wJ0+MMkyP74jbH3bSRgIP
tafmqDwVU7/LwQ/dV6SW68e5ljjJzJgroDNqn2W1Plk7v3yopckBt6zzO5gEn9QS0pGOLA13ms0w
MWDt4SgZcW/1+jxTWITMn8mucggryBNejD6JxD1MqLlJToxrKSt30jbnqERorF7sjaQkV6VFZwdK
Vtp8t6fXzFXD7q58LpHEgiRZ+eJcomoRcBo2Y9uJyBXYN+LYHLbpIeQ8Ekwky0w3rqD8DxXGqbD1
NklzcjCr5z8Q3zQHR4O80a3NLEuhl9fL2p13fMBG0eW0ZqtS3bTbDy068PNnDgbE8Sb0R59+t3Xv
0Fgi1GeG5bpbttyrMxWSI6PIdC9nCzMFugUHMkwY/HbPtkq+oUwd/2ywK1GnZApVkL9IibfeH0Qc
0btPtp97AVEK/qXT7ZmXgxIGkNbDSVKs6tJeCc0EkWTcq6McwkNbk1KJ6Ik4oigmE6mDtGn87ksY
9sl+zlqlxItF72KKn4+jo2ZtWWWOPtmoavw/ECwLM6RWGBS+CpyC1s6SL2WWalG+ZUqiOOiJpJ26
/NyHxlKj55Z1zP9DJzLJX/RGbGz8irTIv2vllLT8F7eb3QtQlBolBMTBYX0d19oeEUWP8ys8mmFA
R5n5UoVaGQpb9DkFyk22vp7zHyZaR3N52fdBpALXxbuFUMjyVfiiLggE2l99CxDVVwiuuWOKhnHe
aGjmtqqoWxrCjbHxx2p+JBSJLpBq9+sUY8w8tyNIjYnqH5mu+e+NK7kN91vlGQERUj5RFz88Jx/h
iIJ+ttm75JE/MtAXiRh2iBOuNF5UR+06NXDCJZzoCrsY4/bIP20QoaG/Q8GXbTQ8NsH3MxN9P8El
JHg2V5heiDBHirclJdyQ2pjFalFXCx9D30hUcYFb4D07x1ooC1neDREn0JbjZ5OBeGVUHXkgNeqB
OK4K8kunbV3+yxKjEV5w145KHg0JWd3DgPsowOa+dkLXIiJpTSXQpb0HXDbcql/7WpRRYmtyzkGB
YDbUD2vBEeuctB2RrOf8ilMvEsl0X9HdWp1VS+5RqSeBjyqzXuyeGmdCc6AgR2upEx7/JvfmK87Q
T1Tq53ZX/JBc9EJ0ZZbGG2qo4/24/Joo49FzkAuLaNVcoMN+ndUL6dSJ8hGFmanenirgbIRBt52e
l4vxGC0bu2JpaB3MyU6UtFJCSRb2so/yWKQlDmntq2TQCR7LPC0OMzLN7p2wzr24bC9owLFzISTL
rlwgGOIFThyOJU9vOy3WuRQIsErOcg4Ul8vLD3uxzTBX58As21HxIJT0IFhyJHX1Lkh3mSn6ZsZ4
JBgA/9PoX514DVjh2+oSAzzWyYYV0qXkspP1kZAHbrBy6NgP2Ye04uM3VLqZVcCtC5sfUcxOt6YZ
YGt/MIyTB9b7KC1Fi5oumWsw395neeAdVQf5eOcNbcfMRwTbmKM8qEhwQVQDIiM9dN8PtnCyJYWR
p7/32+ZBWefOXb/Yv7do9j1zlhTnyJzFQYkGBVF07vEEgCgcx1Q2kCtSZCyO7xKrQIPXJEYxrdJU
aGTymCL8rBSgs5SbIIO0v/q/noEuLEYv/40M3k1jJV+knsUyDKoCoqUuOaCmx51noCdxrlLxTPFV
x3KU686qx0zh6ruD6FEBEvfEl3qRSQt1SNRGHgkDjIAsU4o1gpG0JPhtqgDAO3T5vDgtvf+3AZc/
HljfkWb5RzD3mJEf2FQfiAf4oenJSt4o6pQdzekX87zWqmPTlWUZFtKD1Z4JUIA/oOU5fK5UZgoE
WWG/3UNI/XYnWLamUlbwgcVUxyZ3/WWaInKV0LgvV6IUQ2pCNqq+itezjTycWizCxmaF3o526wus
zyxKh/4VtEQaqDMLxz1ZwiKiRjfRjQZ7pLPFps0+O6qaFfG4wVGV3fw7F4PppIuHUah0JIvjeEDN
2fhb3QnPLMV+eOG3hkd0I/M0i9niUjQis5ThF01cpc9E3iVlXKmxCVrJyuXd8A7POg3xZ3SFmw/h
r64q3tVWhdV4wAv+zO7Ui1FY4sumGOGE8qUEKwfA45vCOencgaPfxuWaUflLZDVxuTLh0X6/5imD
DGkRds9vdC9nE5tuv/T0WZjybk91di9nvEjt0mbU7vXsbjwFFwB0JbA0dzl06nkhxIj0v3j1jY+d
zrofbIBb6Jts3nYyOU6u8UiWHOIsJDVcJECHbDsQ4LJCq6A5S5DwMDaO1oWfrIpj1qig/mrkEkPt
gKivoJbiKe0raGTIno3bLiKPc6yMs1AmEv6VHXP+3JavNlGdNP4X2dxZxx8fD4Y04YuNkZ87KI5x
f08QC2SlCDtJFjnxZOWPh2BvK5SlJCj3jjlDMNmt8ZKvSZObD1n8Zm8ljuDnKBzKlihFrpo+hK77
aS7vhHbnWJyiiguoutmMjkUv/yNzS8T5NcMitdxDQgqbBT/QOOha0cdjDZdrZY48j/IzlYIcwzLb
SHS2l6T9pAIPYUSWh+sN6Hc3e2U7J0dkVR+AUqst+kTcnXLYREfB9YOEXo6ZwpTl96pg/KDrjKUi
Y/BwStroiZyAKyL1CcG1rz6HIabZPvxPJAgLsqnYfe8W9N2BXWq/zH1+jKGGjj3bQBkbjLyiUNN3
3LIlkAvx9dsOeoWi/gIJJ3QfGfBsgqAZNPhQBdu0Gv0x3Fktlfjt/+TVJ1b1R4UZfJiVeDQ2vFHa
HPVdV/sIPdCE7IhMNbD6w7ACZEjfKy1umfI1unATEOPfbKkmlJhpTIWMX/GNji9DiGL7Bytqzvug
4V/p1KDoc/FQxsKSMFN+1scq1OJKs1H1e1MlIbcne46tic/n9ej4bzflDqZl22wb6CmDRwOkTSHu
S/735C+vmur2B1MqP4pgcyKB7tgtTDWkEcz65y/aPzigETJ+A+L1sesA1m0MZmu2c5S4TPJkICnB
kgxOVkdUBymi4UA3EP36VN+vs966XJ6JmLbmCb+oOr1udk0QG6ZNFKg7DdqY7jdTutdF2fNJeXKj
XUoGe9yGMvMcJi5AW/zB0vlOR46cDLwK58BJwd0tg8AZCzKIZSuTXdsmpVrFKUBzBCFHm0KSMzGi
TTvb58Mw91nPSwGMwJ305J1/SoxrjOH6/YTJZ/D1wwX9+wh+okzT+i4OMnpX75Er1gSSJam4vV6g
3mutZlfQruLCve7jQEuTzjqTKjiLOeRJHOCVNv80lBbNpInTNYPsiTTlp8t1pwFkxl+NRJ5zd0aE
6Wajit4oG4Psy22ChAOvEsk6AybWo+VOPUD90MET57zbnIfeuTQ/qhXiQBTchfJGZkX6ISNTKuTd
ojWbE8BT6XZ3s2F3nTyoIewq93/PUt2iNdeADI28CISmhaNZw5zQDtcvwaGfuDmNk3D1SE9zP00A
uSeTU5KFkUIFG24iPAABMnud30NimbqXRKmlngyHNyoNNjWu0N+72Sr1GWKTEwsQxntjGEov3w/s
JsidZ7i1zjF0aKn9PX85bUlLthpSNZeEpKK2dNxlKCNg9xjEbGfsYDxG4F6Nc2qLHFjfSvzVH6cr
R3OzKDXwK6WbL4+I4ET0mFpfYF4iin64v5n/Q9VjQtPdSQuh2A85nuazGJropPDy0QOz1xJTTfjf
r/03+msZmRIM9obSc+IsMnh4aMGdW7IoJqNMneHIn+SUCprzkjyt7f6iuc6mZdyuaFZ7BR7u6ksa
VnSZ1fjfTL4xOHqkK0kFOX4RHtezFAogAanXk5Gp2MLYuWyVWWZrHddCHqgKUYaZxzXT/nLxK2tR
K29XXMtphzQa6e+UFz6Qj5uc8QM5t4/OGduHpNTOILsrbJ4Lfb+k3t4cypiyhEt+hDAmFHiV60zi
hKdwjyC1DDJbjBKnIXHZAN2g87r9YUlKHhfqVSpyHhh3XHi16uN1pXKGKXZOjwQTsepk0kO5l0Ql
KEurSAQ8b+HV1Ne3O1iV4oq9uh9YjGobYLr0RZJca+aaJ52gJ2KMK/lN45osTUeB16gzOLoR3eUS
tVIQhsNItCWBYsVTqSS6KJPl61Fc2KKR1bM+kVZrMuxl+K/00BJtEIf3JFiF6vXPNGe4e++0xKoV
Wrho2wjTwzjITmZVKCWZiuzoIZBg+Qe9+/PK4Q6eiorkKb3Y6F5fugDIyPyTYMNcNqngx2LQJg6T
Raksb1u4f2rUQf7aQ8EX+W6BZ9gcFTgItgX0GyMQoW/ShzrH5fcqW91153rF2V9btqewNtxDodyE
FdJnsdO+LcxI0VuepwgPpAGv8fPYhNkNnuvNRRAm+LvmM8bKaPYcYgX6BhvkYDs0po/c5J3eRqUA
O0U527Vd1El3bzDoxzx5bPzc+UPozgZJMwLl5TJnwcwEKszDLLuRfdc3t4FjO2JIBBQPPbOr7Ixh
Cgsceg0/LAaPM1xE1dod5ZSCM7UT7MNLB4qgeH5D/0ONAMY2vecWcZ/Bc9Hjy6hhnHsRfEjtbux0
qukIK5aYO6QKKleTX5qdICySk0GEsraF1Jauqstzoh1IGTFNx21tn+ul7DztfjxMqgxUb5FbTUcQ
p0oH9g+DSucYNffot3rRFeCkyqGkMUBcmv8wtnWPX2z9FZbBF9bCmbL0q/458hx8gZNXtK4wZqs8
2c3t2fK3EpkSnSfjtnfNyJdW5Ay4p7uF4Ozeo+w71yQpD6RiZciL2/LFn/iaIvtm3gzfcb3pg9qc
H0QqJfyzUq4mxDwfHpv6tb84qoGsHm8/JFzwAOVYsGFdyiwEO/518GwH//JQWfMlp7Hg/3yHmLgy
aHw5vnlHdJ8cBvdCQrqrkTXuUlywFkkrLBsT1PqTCIw+cxdRTkzMlBdwv9k47R7+vbTRSzBg5Uli
dZKstGk5HsrDDuEohie4YlqIbB5lFuIVyWIldQjCT+3kgdwKuYJ+suSR6Uw3rnq80KFwWalhaCyC
jmJvfp/TxfCxjOXalHT4UqjMsSxmacjhWB5TdZAb61ggq+cXMnms1wmzepwjLmoXMChrMP/6bPbn
N307GhrAoCWx02ELRrpFDoca485v+DGkGyvdpi2zfLmpln+O+W4lKRh9hYycbbFBSE6qoxhhmWPK
FLs+4h5pNwmHhlKS7cBhy12JgtY0mUDVuRc+3tm0/+pw+G3/ImPtW1vq8yp3iaDrjYoVR34xTMdn
0J7Gr02b4TxGHl5CCgDlYrME4j4Wxs583oaB+X9BLUi50P16PiVHLZMfqCg0H6uDui7zfdGIcZ9G
lqZDLyqXbdDSlulLeS4rD3plV/R+xVMNoHGRYXY27Cy9XkmiamqCunrz5X/YUHYG5BT0YkB9LyMs
Daf2CZai0tKqA3Kv1LB2qxwepJ5mEQKjUKrwstouVQScLMfnj6gKYoIzbXLJC3iOLF4Y3yT/6b/p
8KHlVZ4dem1+th5f7hU+Dd+xxQ+0TEzOBc5EWue5u5Wflvz2B3Tu+Y1qVas1I00rUR2gZwI75HIG
qqa6oINrv1JJ5O2s8lo64ZhtovRuUjvO+OeZZE9sA7XvnMzSgQ+oQ5qCXGwkY3tkgo+y1gvIGT0q
jqM6Z9Bfr8GnEmVQOdhYed6/DARcZ59a4C5p2FvzMX+aghyHPYscRFYCCdsfJoASf6aZAeWqh6Nz
fwGr5JTreMtqKMU0SqL2jZN+p1mpDoiIAtvm1vu984rxE96MUbCz2OljNjqEbA2DjN2Yah9Iwa1t
mSOVPnmI08dK52SfzDyaBEHO0aqkuae+X6kabT4A5kK07xWspBg6hLyF3/ixTbZF15A+X8bdovsX
B1+6tR+dRYnQVHsHsIzZx1pgW5wcEsD3w955aYwhj6c+5JHsR6wkQLtfnOYBIaZz1cQvhnTo6jiO
DUp86Cq0R4uJx3CCDOf+DR3qDr473QFAL6OsiuhFGtVYi3k6ahA5CWzoBCB/0ZqcLAupf+CA+ShQ
cfe+NezEGR7ng351BnqnWTh4HUrzZoQeEOZcttNkW8GZ+812hEnOJGm4a93nayWBiAUcwCb+mV6F
YmXhumJV2fC06mOA2fFSem4Y5yRJTG2pigtgveBr9sGvBPbAHyOBGX6Zm+pg/G9s1PMUtkyN/urc
y9QuAglz1SoufBJrsAhkJhw9My5o0PKE65oM1umatjUBxiqqkCAsMfLL8n/bDWeZmjdmL62BY1qv
cuWFrVoQpHosYGE0J0pu+3IpQ1xbpzFfNVB6UHzfVYG4n/1xLnrH6jhW40CVO34D608w1reSCVzM
2APiTyMXbNq4pjjwxMD1gO0Dq8qyjZ+PsBrrYZqBzMMVeWxL96+ZjS9XhplSvNDTgtFk5X15+PRw
OLVUszCHRm3257BRjY6tX8pOpdimhWVY81nKXC5Z09uxpni7zSMkG4hatuylUsvRr4Rkavz/LOxF
d1YHRaFZkhln+CxkeLAlFCpfwCShwXRezSFVK9TH6ZMnxLxglHtqLOj4BGU4gCbjhoHh+gnA0+gN
6xtBEWXOZEd+g5VYeGSaSmBI2HeqEZaRXSxuGalVExt2tWLb95c2iMzzFPgtmvf5R4ECJH1ytqjM
yeppHDBeVTChzSRSWO+DZ+okdScCNZ1IIok45A9RACcE7Lm9wYe7gCz7bVossXlT3BrRgtIiUQT+
lxHLB8f/Hhpg2tml5fbgOFDD5nOqAuABMxU/NuNRwDd5dppuxj4VRgMZQwQ6NhUA4L9i1dBfv19N
VglLk8vmBPjVv0iY6XgsYTF/AIQfrw5G9U0cKxJpF63pRWI5MFbMXktwqPz9TyJNeOvV7l02mYI7
fOPEKSynwVMVAbC1yQ7jLjJowAOT0P1i56wkbM8RICetd+AXtRkIO9kC/PDJqZziOOiPIlt/m16v
/RVfRSKOx2cbpE9EbLsrnJk6QlfO2V5X8SxGpYrKatfBRGHgimych6OxvqvlEKW/TgDJpcGQeVdd
wyimLbeV99zVNtE07VCSsolntp5Ly930YBKyUTpN9yDw8SQwYfaaWq9+CVjGTejUlBHJ+xp8pe93
/ZQbe/FR97lwxupECc8G5ijRCkWqNP9QNVEnLuGL6AwEYklU1owdlM0cq9v78D7vYu+VD7iJdm7Z
PEfAnv0sw1MeDituRs/4tvAxTS3TxvjojcxHODUvlXvlR9OWXK1/O1US5Rw8ckDKvqIEsamgp31Y
hrpzmFIa7N67qmnslGO4eyRMilfsvJ41JZgjtZHeKT2y9ZiQaVU+GDMEN8UJiFeFKAhQJ+uap2tl
zTYzR6mePUrRG3G/1ZU2lT7YPDlvzIWyU/AbYcBfwQ+XRKjB/k8uhpX1fzo+0CjXJAqVx3Lsnavl
rYxVeQ2RMGoEb/k9lVwPUHNu+DYDmiOYUCZHIDvHS6X/7QyBMwCU0YCIW3cJtY0MiOzIXvOz0vhK
x3BW/TbhF0NKPVPNZXY9JKtxNCB3lX/CMkT9de2NtzyzVwUby3kHRsMQ83+QktoSzG21dhG5mFXn
JSc1KXcrIu96UrzpxbZsnlvdImxuJQ9kDsDjAsz6ZTxSgs5fDJv+on7nTSjK6ZSYiqwZLmqKcFsB
NOyQehtmUalOFNs7RSgYJVKMP6t3pVHI28WzMoBp7/FGI1YliE+5GRtlNuc5gKDyX0EZHvEAromv
PhTnfCnbpaUpGCxJRCN5rLegfObl9n4TiL0HbA9LfNKt/MDpAy4lApyW99+Z05HjpKvx0yBiEFoi
h6aIH+kizypAWxheFkMagjzPD0Jz1Ap1RjDbMJxF2EOBRkQNEwr66OfCr34iy03mIQo5dREcRc/j
a0UJleF6l5svEtUbAUSOrtYl6Ksg+5xt4IBO9zE6yEBX0GYVuLuB0oAKUeu4o8q3Rv359kU8tBx6
PTej3sHZpmOa0IqpdEACKiZlEGc4qmAX346kXKOKA5zhleYuyp80in957HAvjTLsuuX7N8buwLvz
kWZPFld2eD9mLuBH8T1RHfAYLhDl6tTS0ehjUqaQb3GFTBVQ1H9DcAAXyOZdS5nmVtvuIpZR7+gq
RNgFcrq1wAux6WwdO5drnG7RvSNFObCrahQQxtkjih7iKV/2LqevScVdhRtoiSuGt2TdvRY6yK+J
c39I9K1wYNaswbSV/OwMORN8eBsXy19tt5o2s6H2bDB3xWVPMYojZrakyw7syh+qwn51U7qYrPdF
MXj1xqqv6Op9JUvva43M9+fIom0dY9cjLr6b2b3ffi2B1hsMYSId2KsruR1GWRAkFo/BLW4rWeSW
ljrfNisi0leXWZAzPgkNtR1wiNjFfPNzkJcxhwcLA0FYWWjjEzjlBaBPYBUn9hhjz4bFyqTyd6i9
o3uQHQvr8SG/gB58/ygV6kRt9N7UJcyNOEGVOEa9lDgFQBeACx1k/JcbtbpkJOXdHY1+u4FVn3cQ
Ex9/cwXJoh+XggtzWO/W5owQsag0LUiaGgtaekefSLIJs/lnxsSpLplqgOwSb1kVMVZj/cBffOAR
3HrMck512HNoX5bS6DXRF92fY9O6mEcG6RacwgSJNB05m+bQoXZwCmGjAb9E9AnOGZmYb2+gRGGJ
hQjVf96yYc7+enugutYeEL7/JLlvyLCyOu9Vy9F6k5eukaqo3W9whrS2XcZdyCCXXNOgBDAT0kkB
BmP3rQGl1mEZmrrKQ0NUMmitls9Xn02vQNgYW3QzmHaEQfyr6zPqr2qgNQtUvNGI0OTenp8moiWC
fIIgvEVqjOfYLhGEwxVed0sAK74iv8pMgMnrsvyuAbQ/aHjlkRl1Om21464v3drNw4cE0dsv0x9D
Yn+UiKwZAhWr7hcb3b3jlb7KTQaysF14Xb0Cm4cVW1H5t+7iEh47U4vjfBajP+Dp4+2yvNUz6U67
dLKWB11aalHwCtPV8EEboLvPVTMNv37UxvxkJDezcj4hP4aajbqM5+vEuZ1TIKIOcePJsBUtNCiq
zqTQU9iOaFxxU40lKMhZgOZjOQI14JTgazW6srWCQ3k4BK5aMvVnu8SIDeHwOGHj5qZHeuNNeVqF
OeoWMAE5axRF9F+QbkeJtkyDn7FvJL73FmCROHu0drLHXn4cySuVoYCQ58yMwOX1KUSsYWREssZW
4HwLllu8dZ8nNN1moQBsgsjnDUbrpfTnAw9BCIKGmg0JhgdIaanAu7p5N3ty4V3xzpHRplkXSCMg
mG1Vwsw9GrQJW5I54QvvHKEqMltzVhgx6UifSod1tsoAhTDuSyPTw/06+d+vzMkc+6YLJQ8JOE4z
PHsg/NwmoBCGAPLIOAkPZH7kuyjfsV4E0YcQRAnlYZtyp9adyBxolXW0kkP+n1BTjj9AFhit9Jdu
qQPnxt2rQ2iAP06d3iGUJMzuwQ/QVLGsVGnbZORLIVkO6/tlSXRCwZcCGgy7mdIh056Np/g9cP17
MqniAR+1k7KcZg5UnOrqOmSaYYZLHJF2INy5ldQQ97tbWTVHycJPcWIybh5CCzZrd4LDGMEUXu5/
AIUurQ3XU5csfGGHEigH/BwrKf2SKRr78QMHKQYPE4SlRNUTL8hiyPBjTf+tXMGoRie1lSh3r59C
qKX8nr1fK+/qB7lYG5ikqlU+zYuKynyj3MXkuB6AXEtsruyrh8QiiK5WUP+jxfmZSY0YW/Ltvn1l
4z8/5BTWMx0+kdOvDDnkTRqZz/Zw9+8PDTiP96eqflcUWC2AuzKow7ON3/1KyOfO6zrNagISTbNG
VaSoL0odiokoOIKkEd0QrX69HE1JxUajtBaGa4Eeh/dpD+9mGZV4QhgFnUmYJgvfLoDLX8fuKFq1
GVJ+zMq3jK1Q/h/kcAaSZFMgallpOV8PO7Ao0sXt83D47xj5xU70UwbayWSrdW9WUeLnW3kOaf+k
mCmoPUrvsyiSqsubHaokcQmPOw5UvO4yEdDUI9at/sTcSq+Yz1o1lENCs9PVWTVJIGNsmzqZ8kdQ
6pUe37u6Nt0A+bVQdH8Y/L4VPpTT92Zq/McADDBuG64hGUy3UyAUvWM1XiFeoTa+jHpylNpX3H7D
oGBAOJEBiM0pBYYqW+XVO9i6a92m1aLPRq3OHilgw+0zYFcKYz7mD3fTfVTgpNX0GszNWsap8UuC
0zpwfhv0xCNEIpZTpPbAJchCdYFWVL9IQuHXhK+MdDJcBknaP/EQGeV7tYKYckx/grULi48Lj+Ft
eCVOzzaq6W6Tln5UwlY+NkIpe1BnGzDId0xzQJrttGtCptsj7XplgEGd9a9+wzZz4PJkAssEQc1J
GH8B2Q357PF046XvU+PfLhMDOSN4Kd7BsM9Ja/u+Cg+aIiU/x4AXrDe93X0fZNat8pvgFhch0Kv9
iOyOsckInn50Zbg+lu+5Q/I+OtC7OAvp+unZLtINyCy481jtxWCd9+CYxY6oOfAPYIkd53t8CDIx
MebAy5aMQL6V1hgjKg14stQ8J+PleAte12/1COQCYG6+4s0B75PlZFwjLywHsYreXsJHgYwIKMgD
4CP2buZua1qRDX+RQCE9symCNmXoKvF3R8oA3VFVM9Zpzvyv/KWed/mssFsjtb3nuvGR6XtcD8U1
uRcSdJewqU5pQHarSaAze9JiP+fFYueibEu/2bNLcVWWn+gSQtKvMWsvXPwEzk4lZf8tMKuZZuV3
j4XHi1/Y2csCyzj9L//psUNg2ePIc4+7BMiUvIo9pxPkqvERG3zG4W8WW7aNRNMOXXdz+UqJj5h1
9ILyf76tKBcbbPj0LowpRV3Cu+IrGrUOYAEpf987b43Mks68mPfW7MLaQIELYyewpQEOy1UTRyEd
pDyqsY+1W0WFjj75n85PMZDqs666VojXqSZuvC1LDVqDLTGOlEAX5UuXx0bqgmZiJiEYJloLcToe
glosFugrTuTyZeARRvZ1SKjEeFdL/V2ZVcWdizhgXFGyWr7G7B0eb2Hbu0Kqt/qGd1O8ZUPyn+Hk
Jo0lzKtNNLDiJLgGZ2uR7fC+oSE0ZU8g2fFzx2QdyIeXJZwETdnNWvTP6wQWxDQfLOtDa0dJiguy
EzOV9YFMmVV61XdPL+gguuHpFLwQzPnURYq1ShBuvzvC8rK2KJu3yDFJWEDiaVNiXWypvJae64+z
D5dN5lGhX1WgMk7ZodLi3mSrCZJfVRzA7AoN5hN9CHj2pjKhCI69lVdsfrWOkSZFl0+alCm29FK6
eTkSRRJog/L1PsbNySkg3vpUmShr6GN8zG9s6RBblrwl646K+cpKwSEA8tq2pS5PMvOKo3dkAtf8
ZwfV/+SYb+3hyxgbwIOeemiq8qv2vyj3RFuA5pxezTWypCQXGICgd+pzjRj/aupNngZVi2Cc8lT7
C34vqVMNqLGeYj/RbIKWYHKMTkUXZdPtUgqusxki58LHSencAIMV+rCTrgooAdZBFLcihRghiA53
Uw9a6Fn8s0z6VMzE+GVHXGtpgyX0xoO8SqNn5l0QxZ5NVLHYAq1WvGL/e8W7cV9PpJfd3z9vnWxq
okkw5jP1kyXGNkWSgc2jqU9IJX+BRPb8bh+dXncydi422oAAmAxBCG6m5ovQjE3QzqeT8Wz6zG3j
aGoVV2aIUpx/7dwBI6O4x+aVouPjRTrKfN84lJNZuNhUC79/WlU5GYehsd54tDr2LFNw18frTkjY
rmtP3C+XeoRlbGxyqGbEXC4rmSOT/yo07Om+zCdOVNJlyMCVKYC3sg1vLBpDs6rOtzkXQ5+76SGM
Odc32VLC2vVHoFB2sAmXsv2sBnk6TIgK73y39IIdMezO1Zuv2UIWOJpXAaIG69HicMh0v/uMc5MA
cEhxCz+uUZip73Z0Q9sX9g413vfR3lMNoF/ZP7ppRhM/HAEQNYrAKA5oypI0LxM6IWTRDFeQ/qJg
M14M8oghHU9k+FT6W4c5PqGMczzB+DANdDOEau/SUC1stBT2Pg6MuD9iUK1TF8UHkdoKT7wN1+ub
H2FcPaP21vHduARsFZVd3POHT728TQRx+LiZpWlr2eHOEfM3pRTYCJN0oW1Xbf/Ee1Cby4sicYDd
B7UqNOM3QTVsHV6lDEPcdKjwyGGQkymuzKyZMcZq0p3HLyQ66HmVwC16RzCkYoLtMdDKWU/SV8GF
7VvCiUj13LKDiAgRSEew+Vorcja5XTR/kN2iy6AG+K3jKlvX+sqyH1BE9kgfPHtofeqjCz2KkGSh
4s0PLZgOJHGdTMoUw6fPlGdQX/uEbWKzhhJTpiWHS0I212QSgcYoWJZFMTAQWd/oFsnTqjHrKfrX
/7/bK/6b9wkCJauDpuyxMggIAd7FlLdBtb/eDFmrVWwnp8cqY+Rfi8qB3TDWdfbAlqRHvWjWGBlg
FQJXBnzU+XCuKxxQkbpLev8TUeXYP51Ukx5aa9Pucv/0pZhoNlbIEBOhxHezRnI8w8z7hbnvK66B
UurelF4lbQV8CO7YHHLmfPnXPE3HjdXghnUVgjfO5G3uFMBXq8vDJ+ixz+ztAtrSzQrofKNXy92W
tUcSwmOhECaFuGBWWM0B5gV81KVMVouogIOtwrfeA/qTGq+C5WwFN62sfkA+sGpi6s+t0LRJ33z3
hRBMrR7y8NS2Ja9zLV+unX5tbBi5k4U8Nm2/SxcXcRoN22IWM06eoR9EPPXLKpQDyyQoEcvXtUDq
NhHqXIPeqa4VbctQFyffEH3/wYkugl+LwfWX9tTwBVJn9D7GkIKp9nfF1wTAtCtip9dxGVNJ7W9s
wEClk749FK88fjm879lJWPgyknd3f8FNSibYBFSlTeAlz/3Upi28/l10oH0SOzAn6x6T8G0EiMt5
JspRsgytjYDF3EYYV6ELLackQl+UeOYjoZpdcnnSo2p6cpMBLqtAPqaKe0FqA1At5c2vgsdhPUjS
ogaGUmmi4pflGcH1IQol8JlRoNgq/SrdQGYwjWKkWVbG85MONgLCRsVMKVrE723I/TGK72eSr4Hx
yM649n55rEhIcQcIhdqJTuK4mGYrB1xAFjQa3HKeIp4aVhL5CLz+QsAX5bckUJlSa4iFEaMLBCzi
u5J1JLH47+Ukjme5/ekASxvn6qvfpz//feD6hWJuvtCCMxGfhHHLRaUIHTnKepjw41jm8CbJZs9q
L5dKGzNlSLgknzdEv3pzH52gmJJSgB/iR01oqEIc6/Fq4rp9ACJVnJsD3DfBOZsuuvRg58jSsc3w
Yr6SbuxxyNyJ9yHbwa4jvz+YO78BGBTy5n6RSFKLQzTC+x1F1CsjpHFfKocJuRRFcMAZwpqepASy
lAmgardIDxve9dyRVInrgosdO8aR/7FYpnyxQbG0fL4h8P9OqXeNdK7KEZ6lo1avOdE7+7LmKLla
BF0RLDEoWocX9YJISvbLoJOxDiVUIkfbD2QgMcv16FIBP7sGVRmDvISo4Xa1HgkL9pNvif6p/aFN
Wzt8OuAVV1ODtePHE3ZCuQyKcSBO2wvZx4YIT+idPNwoLikBNKc82BbSGNAUZdVDoUkqzgRvXBAx
L9+ocJ2XX10INsujTRvhAMFOr92tCyCHeB4tzt1dsOp2I63pCsjsIsmY25JEwCiYpszHyuYK7WkN
EpmaBJVrYzvratLVO2wzDjHaZTKYjd0aCaQfC6icEI3gD94/ySW3Sb510mwsYQL1mH5lmL1d6G5o
8DEw1zDSZIzXht5ilzJ7gONb1mgsmEHYQVhqkYrOKiAKImmpXcFQnMsBJ7wF7HH+N97N+Ng7ioKn
y23rv2zya0qLEogtEwmp6/4kb0lE/sNzp5GM2ynNGpUt/SDCayl4Zn3JDsnZ0JjZJ8NT75jauyvg
8UowbEMCMbJtmsCmvl6ZmSGY6EXo3BB7rZ+/NnXUPD2iSI4hsAdN//E+8AxRvQ52Qx5TkQaanHhH
CBZgCPY2tW5RNaqJwRzHA6REXzP/fJ7g+wwEtys7VGQBD05VyzErdmIulmU9cDP71YgA39yzs8Kz
SreIds0uODVWktNFEtB572M5LocUo5oJucOvsWMNHkDZ8lMQ0KRtOaWLNc0Qvut7nlP9wxSS2Wra
gZgBc+TRuJtK+kOasUzKW3A42ehkfoA2PlA3jA2TRvp3SAOFqhxbu3upY4b+icuILy4obT24QB0c
zipwjs1S6y3jpZKjzWjpYvAbhw50ZBpx3cPtp0xt70XE9h5cuG9tnKRTt8FJkmBFr/PZe8Cr0Px7
BOoNb/vkcEwhlrIERMKMAwlzMdkeal7/kp7dDd4ESLEPJuDYjWC8YhncQw9JqWWvggjFnbamkDPM
fjFrSLWfImfc6cx0NWGojjNYALA0j6xG8J9jXo4bcx3fsm5JpbX6cVQFzNhC+q74GQ15LaSo1w1q
D4KviN+8AqZDNofb7oZ7pRmdi9N0Oj63IROo7VhrZyaB3mGI6ef41Ix5Kedr5VUfg6ZPWu2rH2nk
ngStee/PWfEmEIBlYKpT8OJbh1HSZXjsdTlHEICmC+6Yyw9U6Ki8qeklJbDCDCVcyvlqG6ErQLVX
VDAJGj1/trlHNr9tJTeP7me23JnvqTq+36hpEdILNvk0zYY1sDm5GCcqlsJb0GoPVnOTPlBeGbC1
hB9V9etCoPAwafoCCAjbdGaLjpsniPxH5IhKVSGhNThvEjIsE8jjb2Yl2yg+Zk3Z2W/qWC7MVVF+
klC5yXuHDomBKiJV/lQVZsoPkgNtQZuKH2enzqly7GbjE6Bdrs5dDjKLqg2S6M1OR1/HqeHaNqL/
R0M1Jc2NkiWaHsstsVouBZDBVWFRt0oN7V81KJ9M8Q4qeIm0vBhpymRLKFidKWa7EQZgZnEna78D
ySivGMwtlw3yeJjpIo5oilpQg678oh96fpZVE/i/prrPzqUawtU+2MtdP3ImKXIl1V+YBWHQ2Vsn
eCKWD+mA2TS/BwkfjLuUeo8hzbwsvw3GBsG9ryKap9DHljcKRYRT+R9RI41uh6lWEIFwV2FBvsd7
4ZyWncRHnovuUDrjHfHv3avb7SilpCaDCfaCGDYZzkjlQpQQsZbe++x5LeOpMLepOsp47APB/nB1
rf1kp6sJVXfVvCq6yvk02qH5u7I1W8vqu1kQ1xRLG8riEvL9J+zMBkJZmWgE61pNlHJpfwiLwVsm
SFGQc4x3T+P7uFAI8RnewvSsai6HUWdEH3ZiSEkok7Qmve188FtSRcOiq4dXR30qSGiXY0P/Uu3J
wVdihIJ8UBwhv5a5A22CoLq2Uqw3LL7G0s1cTCkN4XVFN9CY5/5mUVatgLL13Hq1i4NJW6YmvM2v
5TrI/HIPvAp1sbBhnTXTCA3gDGPbdMrqCPj0bVahYSIf8pZJC7L7xTsesXWZMHROi+eNUjRdIfzy
sUJOnqgdTs/wQAYXLZai3hNsILIPjwH6R4CMFQUjcH7kzllnv71w/5yhs/VciTKGd2slY1u7jiOZ
ETD7w0kjb49s80tUxMYm4hevUhIui4rAj4gYjHMA9VIW3kMxmhB09lNaZ5/7DnvxChGIjgSqsrmu
TORjYmWQVlVetBbhYRIF/H0AsZuvWK/DvaVz2abTl2uWqB0ox2c73DW5M97JDvl6eBCa43QK4OsJ
Q7moxzSUXVBXljKeZ8/1XryeKhXruqDrJM+VyeXKxPb0nsMpVIGVJiJPtHLrQ1+h6CWMKbpq5tex
+pPvSMBnzun3uMTfu8zJo/NbiWv3oly/Qo+hbpw7fpNEARrb9Y3koYZn9QYvaJEtwYjV5o1lwhsK
KRLfBEtuf6NEFdur7QwvLp61ARAHdbwpfeR/87PECUG2kZRRYXY8Wckyl/IfXZ0wHaGZ+paEBH1Z
yYS2fZIjCOTriAiTlLyUhYinrrmPr5cCQblGyj3DZqEioLe+zg+4V1c744o/hq+vti5HxYAfHvEr
XFnEMtT8ZZKYFOcr3h/zz1LknxkGNohsNhTgqkTgEU6+WaKeD6EcjieLmvWvhmsDETPKl3QTHiMH
DekEYZ1QQ/p6s7V1NO/Yre1Im+uaTPo5wcrbzFC8nBqeNIUKg93TlwDEdqG6sY/sIjbZS/AiKURk
PfQokYMlxQXIccCCa5YxrhuvT3mz7XVvXF70jpMOHAs4hPkZ8+zHKUVQ8vgUyp5W+WtKAnjiV9h9
AUhVb1KK9EGT+VJXcvJn9NzZmLRviwSDE3tBWEyQf61yExhIBbVLKgcwEPivQLFR9NTSaQYmn8MD
yMVEsd/avX1aIIFOubSCnyqYLmQN9Zrna5m8wnJmnggJbSeTYh2e1L/WtSntsEObXWPo6YfwbaXU
MeOVMyyp/Gug8VRqVCCfZfqfwuskiDoCB8c0eGAlt1/+hPkofRcx6+hNEGFxbVeqU/zM3HzuE63L
ye4SxT4gqfXNSHCLhLrhXdWhg1dYQJxCnCZkpnmusWlLDiZo2SSmlwaFdzGtIJf/tQlgv+W90ks3
L/SfxSKDTDN4/lY0tsqI1MuUEYAO/5VCy51a/eAMp57jb/lO6xeZjWaQmUDY9nmBus/IRG+EdSj7
jlEMOEpBiXLrDZTKKhaHoXhzIS/pL9IWOdqbx5CyEqXAtaK8CjyNiz18EVhyYXSr5SlDcuwKUOcd
039xoZWJWTrH5dIAbTX3DoAQZ/vVGeMrFYzYHm5WtXNNdI++qy0FuGWvRf1/AXedm4qFDWhIiKe6
fjp9VfER9N4u4xWFz627ApN5isBS5O7ZvrnbnYv0U+9yF0d6QeqG8EHnh5hc74tjxsUan2QXiem+
eDpVLU46VD0HwSjTbSn4Br+lqK5F6EgmhAJJ27ZDQb86J4zRkhlt9uCz5jmVTG1beYky6z3EPRer
QpO7kOLCt8G4x6eLTB0IRVc3FDooqPdJN0tOmiM5HdVcRQ5DuL/cFcG3uzsw3AOLFreN6dueCR7o
lbipd6+Iy7rk2jDqGs01JZ47MEDue3jL37NcSipUpx9d397yjn2q+DHZZiy6FQst8/mB1fLFTNdK
sxr6VsU/LI/S+ZDkBD9UjbczUFsy6rsVlQrC1rFbmV0ZkG1ITOAELrOEJ4BvOoKyGezDatoiL7GW
kKZteVuANIilwta8YYRYiUyQhb/2PIRYQL1awSy78WYnJgpvpPpxAr2eEi2gV6ehJHsm2EHZf/m1
vArm+fRT7QsR86F3jftBW4f0o+xqP6u+uEfwRBjlWm9w4gHAb1D3MazJGDE3lQ1GF3IMTc8q01Rn
j01VVW5vEeMT1np+qPaDB14wqteWh/mpxaLGRLIHhgTQKWA2Zf4I5euPoEczLySJlYzEIcBqjqRG
YIQjIfPcBUAkMT+xXoQklCEafpKKqBrjrw0rFpy0Cfnt3PGTt5N1iuX/Ll+1h+wp5ArM54sT72Xh
MhhemPP6RWFfLR1YoIunl7kcgZtIoO34/YdFYACDUU4GA9s/fDCqse2KF3d6qTFgFI8IePbAZW6P
4BqNza5/zAhoKiCJBgXYIaBBdUsnFa7UiHiQ5Il/PJKyP7SAUt//Q0ckogoaruo064z/N74Ja2Lx
tkHL8eNxkq/if+75AtkGS3igS5NhN6O7WIFQGsXsDruWnamg0lXK4hTN4j8VGd36x7Wpqwr1AnR8
rnLwgbPaOB7ZH8HAocAojBq/GjxA6+N+OLiuQnPzGRG3zWmFOWl/dp2cUBST8ms313mpiLPWO6ka
TcnIGiMuX6fV7aPTtvcp5ddi69lF5rXoolU5yNg3wUPlcUQem3IjEn//CgpBzD9caT4Mzkj+Qj66
L9gvaScpK6bZNLmN04BLyKbEtuZsZToDqaHHG20Zg3CR4O7JMqW7WBIb03qBi0j7FVB7tp/X5sw3
i8g8O6vpKVIPL/Lc2mTySbDA3YHQGGCD6lgMy26x3pGo52KItNEPOWj/JdVtEnM7ppNrS6uDEBjv
fKrt8Sr1B4dUGpYpZKvCpY2BSX0CcKTTh/AppsxxIgBcYyfcHp1X8Avr3qjTf1iOkUBB+SN38yPh
7YQoCKktRBlMx4tlY9mKKP9d0X8arKTbXLsi+0uXIGx4KICwzCdjiYKldpaapJqWpTC8UN/faEad
yCiWsfh86JRvMpkvlbjC1Mgt2L0BXlLnGmUhmMDniad8yW89yWLCaik75MgyOHoZrVqJ8KkG+AUW
me43+yehMayXHLjgGQzJnkCUgaRg9ir/43UTrn9bTKe8Ql7MahTg7SFreEHGP2MrI/wAkyWBlpEo
RW0x0IvBOSTq5Fj6mB1Ur40Lr7sVUjp2+G70cVfbE3UvvUo+I/PsMVWRtbZJjz6WL1BzuIZGuXA8
qUpAw3q4GiRmb9ARsE8wdbNtbUINXNqbV5tkCjAFaw7tfInOnAdCiaBoMvfl1rh7apPVMhsFqZGV
jwmX5muPTZ3D1ilKOZqDnkMxp029lTEXBjgNcqJ6qXStjg4Vbm3xlxnClBaJVo2wXnJqwPPcyXjZ
jnwvxSUoOX2gIv3LwhC54LqW+mOZYNxxlvQOBqke4qj4fPwPBg2VddwdJZpe8PDjFzM0aELRwUY0
OF2ZoqmT0+PBOe6ogbI9ooZ5KwYOLmgh7rvVin6k3trLOWAkx0ZuXJPMsIMjpHVl2TgebMmKn0e9
5bWlIiNcGtGr3Y/O5x/w1It64KMLDJgnd9POufsw2xzpq2ELj98TUxMsO0uq9uVhwtNZbxK8k3Ji
aG1BrQyUI9tDuOvC2SRln69efOR8ZguXHyDv7nzhS8J7AbJ8R3EUfQ6DYG/AscC+UephksvGHCzH
4yx9uP6mh2LG51E2wgggLFu67+Lur6E57PZ4Mk0o7kMyDIjn2PH3m1KDzuSmBp01z+pKfmJyBYPM
cdO2+7NvDELhiLbStdD3q8WKQwR52RoRRFtj5jV+khlYOHHjDMechOPX71MwjGeLFKoE1ZCiZsYE
paRdZX5rQpfTTwdMbhhryaWQffe4L5fjc0jXSQmES6NDhUdLd9uuXLH+0bJTYNHeGDbDxZ+VELML
ZTK1U+J3bekooN6z+eyu9aOTWNIzasECrUVGxeBAMs+41eT3PklIvmx2jw9mzLW55zyssYc5rkCo
xQYzQxAGtaNCXItUlDlYPVfRpn9afcRuCk4jM5yavcDtn7K8vmhvRzsdK/D8MJGOhi9K1RANqxZq
h1kCSa+e36en8kGAocfQAzA51wRO1eW3/db0g4kxQrni60Hag8LaniQw0aCoOh0SECzWXVb+Am+D
56kl1cfonxiMMRzaK4oPmwKWPhPRO5C+R18EsMqC+e/IORTUXTHkeqGuRb4vTGZhKk90yFv6+Qbt
cYInDeVAa+QF96Z8pyZWfpk/AujichJ/gwwRKROMTTkOCGKowI5Xh2iMqr5M3fUFgnAtlkojtB2c
C618B3huUAhV/A1ASg/nZKYchedQ/kzofDUxaFeepZvOpBCwTsRp01tmdDJ8pEtREa2n3eZXMoue
P1OAqMCKXI5ERkIN9BWgOlP84epe6+nVzEFGaiYaysclQw/+0WboMMCTTs+ckXq1Vt8wzMKJruNB
1vfScAzwCNmS+WF3iNzHplbuQBvoQB58qKj/aEULYJHaieZkK+NDzGN0whROQIhol81Jh1Bic3xO
Gui08lVXX2zVK4COi3sc1ajocqxz58WBQpOkoflADrFyKMKToCXVT6I+RVGX63Qjlp75DpRlC+od
2igPXaBQrDIk5AHKX51pocjVP5wrrF4UYglzET6ut54m6n+aqxDJaJawTWYH7cYi6mJZH8bshj7K
uCrc7MN6CiYl/jHsSeYevDQctm4+CzOp9WVUzuHfNNtwDo1p1Fw7X/wEWkARbN9PZUaczbGTy+3p
AzzLpXOcxc79mAKF3XNeNtImJZqHbjV/nqI67AtKg1JrMZktykOAbewsInacoIIvHf29YlOfHFdL
gdFNbNqIaK/lBzrOr2wBEcGz60hKZGFk5iKe/ugbl6rMg1iJPuBv+6BVCD/uZUwos2P5fKUPqGzD
udyxcdHzzZTLqvktKGpTsvdZVuU854eaFfo0PGChLlcH7sGv0+wDApcLgfLTKMLOJtPcyKmkHLSy
HlAc2em6BIOb3aQDZhKsbXJbr83CmM8Xc+GFF+e1A7ME1GM4wYT9vwf+OFPAohueFPfsW5oglLZO
DoG49kjov8zRdX6o3r8E90jqaJA1I9Pwhua3o/BL/EiYNMyVbI5SMz/lThLDOObmAbdwqrZrHVTx
EjT+bJqv9dIv/T61gOrvAeW3pj61ljB4gwHBH7NwdOs6i6U4VZk6Hm3WhXMnHONqNm9PZhZoIxR7
PeXI8KEN0JkIhN2qF1WqyPxQVyd24OXdyO33Ujsg5XLVWbUSFebsTolA0J1ZdSWfNPS42VHu2fZs
eLrvRUQ7MDo77Gaos9umeImjJhkEPnvIdQQgYqrmUXi7GzK59Y0D7q4TtSs2CQpVkZAQh+gnAClv
6kurTRWdedrkwdSqqgn7JvAchObiekMXQRONteGg69r1yxlM8A76E0JUhxvHPEFHY2AWHfTBwvKU
1AIKTcOAL1XSsQRWWX0grjrmyWg26eAi/Tfkxx+8ib8ZQpEZq1pcGZvGEUxaMOiuqo8gRCIcNi9W
PpRP/Ng89VyY3hCJTGiikU3VX4ifgIa4vocK92hs5k/DGLK/4yoY1ExR6zKbEL0lqGGPhaOCYNGm
1XPrhZVsOQFG+42KIE0F63sW7e4Tyx2hruUtogsylQ0WokwUKfDAbXlKy0IvhU1jeX+JJsOoucll
5UMnFwOxO4FsD1iczyZQZkH/A4TINdPzhpT4n+1vN+03ByA4dUKvhRBnsSmWzWxbtJ/37jtNR5Ay
FeFbMtIewl5HtRS9Im/GXt0ON7sIROul72aVutIE4U5RdbeNnBuQUfox0LRYBTGp2kl74Uay6dYI
1BgUnaS61Di5Q3Pnanz6Alahup9cEraCqDGNZd6DMjHIMKbb2o+aNcKXn1xCiVpeLM6HdKiNk99u
+uuD4tJFm10TYXbZWYBg/Zs55za6vTViDUhfx74xBXobPXUBoBcM/TRoIzx9jm1gGrSzCKggCTTZ
0r8T+RwTbUwQBFgZDFS5GHaHs+2waV17EhwMkBafrwQ4uYrBrn4NR0VpjQ2C8+YiaZGXlS16qyCK
XK5fY0IXq9KTn36kdwUvPiMFdV2BVz9ChgJbBBHU/FqXtnn3HQrltdUIazqZ2G48vyte4B0dxG6W
bTudDg/a1y46e2k3D8wWgW+BPiHZ8vhlRF0YH0KPMtbirK4gcdnB6MNQ67Kz33E0sIJZYS+g4Jk7
hmrLZFH3AUf6iSv4GEvVO9hPOx340xDx0NxpZupsFdg5SQIAD2FuWxhGcTg6B3NhalBbOPqZb5Y7
loOVMmNEZHOyyNkFTIteRyNzFQWI5SnbRqL+uEhHsDgVoNedrkTY9jGK/7IvVg5oT8zILF2DR8lb
RxClkaXWVDGBOUwCncjcHb5WWwLnWJ6qlj4s2hgg1yiAgLgvgC/fMeClmc5QDKzUVUVs44MWSN7J
2Wb8zX6eh0ewctkOOmBCqDd7DirzQYNfAUvBsgjd89ShSzekLdqjqp5oXD8I8f3N/GwTuPEUIylB
hrt9bwL3kQJsOIKg/xlHgXxHqvsL6As/6OPb9q9ZaLmbAO+RkbbLAntJteO9AGYJB9CADrj+BjLz
i+VTNeoo3metwIEhVxC88ykLCRnK7ziXFoZR3RuygKs+xwvc/MESLY1JrugOivXJUDGPSJ1ofnhk
Dwb/rd9I0sFPE8iTSlYSDe3vJDXinvQX6KPtpR/az6pYSVz/+1p9845HNae6Hfgqa4gHGCfdWVD6
3pB4QneDq+XgQbOtuklLMMpPGlizGWdaN5bh65PyGt7OVbHWBbTRN5GtfuNEFc8mMpv1a1nQQj4+
shWcRq1sOrxN4hd1iRDginbrn+yIAXJuq68BS6TeXoQHrw3ycqLhOT/BD/OSIbm1oqSJzECiryVd
qgrrMa8G0F6PSmn5BOCQ3lu8kS2ZRL4/8RWYTntijtc9GY5k3Hu4ko0alun9lvoiAtS0FEYrAxJd
xRer3jZAxQ1R9zfVX2DiP+5x1kwM2WorkMD1/QxNrLwAR2BNX88uvYvHFLqQu27I0xsrzJLBsBNc
+iKaDfom06NIM7XB514S1/WD3bp3Rmc+pmxLY6fHLWmJ+zKmTZrMdpupSc5Hzd7mxxsThtCzBa7U
oOnsvvVs9WMZGOzbkImJpUs/O8sKcpwP3AiiyWgyek5skaPOzez9P0f1YAR9E0R3cYSuiIXGnQXt
A188HGZq+f4LYd+HKa3PrdXzNCi7YrbJZZvapkOMCpn742rNQDawP5Je7tSJKgYFgTwDWDZjPcp/
MlOF7V2HX9ojxGotiyAFRbHr5hudg6wOkja8e+ukKmoveSKYMN0iH7i5u/FN5x+7rdpAVMWgc4i+
zLVCZ/U9fhBHr1PWAgkoZjXUigwBfPkcyVVHcG7JzwFgG5HGMXdp3V1RULD+ZYos6oDfho9E44tn
XkbvsE9kJOYxDklAe9M5yshWf6j2yfHmJPa/Ix3ZfgnWGfrvwrD2BK3XXmOEnfjCrChMcHdL7e9B
z6wdp48UqV2PTO5ee+9jNygVl7NuSi8MDVEpN/5kq463xrfVvFowPEoKzUP/u08fAIT9q+DasO62
WW/tkhjm9mqBebbOHAtaKWy359KCec4jPgo7XhltTroBBZcE1N5dwsSNOsAbfxscVoMjx6RkPTwq
4GuhxvtuRdK9uVL5B+rr+8saTxZyxwunisWeFeNVGGpmOHcO8QX63mMQaSvQ2jRXC6vYfVX9AJls
pXT1etVlfTlC0AbGDT6UA3khBH1MCyQLB5OLEQckf8eQwUR3JqqMGkNPajiPds7TRkO7oMvTbB6e
xrVzcGZBw7NKMzcYD5rgjo7aIiubD8BloEqL9ncJqyaL5QwChlk5qcRJIbicZzTwBkH86SMwO4Ti
ddWM4VQYzj36nK+/cmdx978+8mNzFi+nc9qARDZhcYS15YIwKiB1Ep4aFoAFKTIgwmSqWfCQl7yR
gCNVtKYrQ3ygIBfzC9bT9YleWY4yeMqzWe0+bKhxAT1HPe0yTijrl8pJQGYFpsvrIdRuHMhl56Ju
g4Jb13DEuSbJvlT8of/ZZk6s3yNw1MELytbyFPJudPGCcEyaIkwyYxjW7wCLAm8/LaFGCA6XEKFa
of8CocVkS5cMa6w5RtUFpR2Lcq4k/DYIbs+yJfT5z1QnCS+iDx7MSnrR0K/tehOqZl+FBls+Y5Ly
vnoSxvsHX2fbfZ3ZY48d/agf/SCWgddL2vFGOHQRIyridRxNlgpy+vWAPW7weuIy3GhnTy+TyEc5
gATPYk6GqHAdRhdJgwliJrPBSKlpoBdzbRt+cUJv/QwdWP7IjayUJ/BwHZ20vQtqvK4m/wDn6Wnv
PgB9qdRGjos9gLbuTIGGRU/veb3XynJ396skCUeFjxIVi0mDHN51E4z7A+DNvgCR4SmduWuoVFcR
leWqesTlb71EfYAj/usRVTWbx06RfcRzF0QUd9TLmE2FFS0YpsW/VshZOApnspSPKA2AxNnNtULp
KIWpA8icw3mD8B52crR3wJyTOvOgpsFpxvkUWofCH0rGp5ObvApcQ49T2MlI6FX3z77IHPUyia0/
Rcyi2GeCE/nSkgld85c+3IzE/BFefUS7QoeOCg0OZB1mWtJMPxwxNi4AEw4aQUqS1FJSWb74/oTa
iVRwaZNB1Ucmz7l7Ihm4uFQrJdIeitQxExKoDjJeszUkv/r5rDGFft6JsuCavxkq4RBX2H3wbCr0
A7ou66BCaBqku9gt/JGTcc+WBfLfZO3UeaLPkwn9ksnp2VRAj4T4Rog3X7wR8GIjJ083+0c9wBte
toWcaZcCYbLryDnaWqS6ctwvECT66g/cR5Jex8x7rGh5zIcaH7Rl8CH8XUNpSng6pby7+7pAHQgs
xBvtDBg4+KX8T3Q1SQRBTD5K+zcgXl/wAMYzWR2bIn1VGJFw3BSwgaJjcVlnjrAR9E+Mpqf2rar3
fmPmwUQ9Dy56+rNTvSUM7VZKpVB3U45/c28lj//rWhXWcx0XUmvwxEv6pvs1pAFFTEr72LT0llVl
/k/eObT1mwBxa86hmpmNJjIqklKCqehKwuAQwjUhN7e+XKEFk/3fX2sN7CJb26aulb0kfKbksOoV
sbPh0P0o+TWFkJS+00kjc/GQy0hXBCT7pgiQ+Po1sCWLJxNFhziB+GaINUVRh7/OXxvZY8EwH3Uc
Lb3kz5QMApzxWVNvACVAlD5ORVjrPtVR7gKryMd47zwd1JrR/tb2nEW+iwWTSQUYBkEt2KaxDmp6
EglfpxgZy8iQKfI4DhUw3BIkgDJc4A/Am31rHmzXIfip3qmt/Pix5psNeWMUEIz31RVYvopshRgX
seyWpxOCksJa1PiTGgnoJ6OMMzu/G78KgFoyd54fWQ2Ml4Os58HqZvl/+a4upQOOic4NH7HAMqpc
C1S6Budmi0Bs9Vtzl7aLnTO6VYN7ks/MtPY4/2d8JHVLVhhmnOUii2iawc2SoVFqVH8zlk5+Twt+
yObYM8cMP+6i7SuHFkapOqrD9JJLy7naCtWrlrr7mUJiyUeePn5JKvBp50OCRNDL/iDwzkhB6A8b
kLFkhe1FDRmr6fbUcf0tCZt15PSK5Yb9dlTLzID8Vh15KaDHU1nUAuoTxpB3NqlWhx/R0Bmq0ghT
5fEhdIeiUK/KhNvwxKjOEuSY2hAkXE9Aqe1exnAwyycbzC92qUSui2/Buuu+Z82GiXHfKq3CX98g
3/7hbCcKQJpTEDaow0x8dSeKpYp/fN71LNSATybCdCnVGMEvKHxxQ+7ND1x8OPlWu4gixn2eIgm0
tlWibDoTDhhbMHTmcb9H1OVHZ/KAW6NXve86uMiL7mSBjyuZRlptMdbgKav8no0NGAV4E2nk6yUX
cFQaUv1nEKKmha5a/y8vAAa7hwSI1tvm/vcHa7yetqIPrcmpoJx87xlXDfgI60AiEjOQ34FAAdso
R89Q2uDkhZZ2UcezOsO6ZsBQJOlOez+QirjcBqQ4fQECD6NDFMNRga915/AxVjGSIVTUI2tfLBUP
W9OlBXkWY+a1mC11SQ4dCW1xTEyC3N63GVnyRP0QY8sDemDWQ9smIaloMhaaAhMTBHPXKK+Hp2Zt
DQAYDdcXhlPW90gA9tmbfgzEBPHBjk69xJyhPBt/uVOYNlA+rR8AFLSygmZkJXYHruVpCXcB4z3T
Gva80bkAyxJ1AbTpDb+lvXBBF8NOJfjuwS33UvjEZopEgsbxsNWXd5he10GsrzIgvQ+Zc/t2EbuX
CuR8k+PruqFCsA4D9WavJRQf+0WKPbfwAOCwx44TQjnZwoF7qsekF5WnLP8iSd6dHkzr6B3tvDLg
NEiLAr8pxIbpwTqwgBiD0cH5LoPkVhJhWNWk0pheEWzbh6Tz4NAiac77VTF4jRQ5fOjOvcZ02p6I
s1MMleKIjilkI2w94dgBNFtq1QntikYEVIXOkI4RM0lV6xW5tMCy+Gozhl6O2ktCIDsFkL85/2Vf
yA/3sGllHIqZ8vqjMzA9rvqNURIKreMDv0UC0rimLx1EKEhgprSwHS2eeKJxg1RsXxqFfCgImJoK
0JvaTtbQhHiOvZVgxvn4+mwQL6TqpEkSZlEbd/922unzldmOuQj9bP3G+3mNeznCsew51TDEskrq
9sO8j7rdxUD0Y8aZCRCGBG4LpA3xmyo61alHqSk94ApCqMCwGrRnfBklZ6vP8+kshcjuCUWr6hRR
n1CN9vitSbGZiiPylGUgfARR+JYsf3gb0n7Ise/Ctp2HxWT7H30ySwQuEBZOGBJHbguYXwv0jYVB
GJL8J/okTjZYfbT95Ipg6+vGoZnxctvLesnpSGGwVrYXzA8TFu0cKaPXNaRguvdzn4bFuY/QnIvz
98K7G8bge0lKomIOh0xnPqLjttheCMITGxv5G7umfjuv197ZI+CN6Uabmy1tjJHRcdX9DwqB8UGO
ICEA4hwIJak17GsKyuzjEY2JkVQYZxBNLegSm15IbaML9dmVToVyRSzJ99ydhxZ6ei9KFyz1y0oV
81BaHN6FtO1W4PH3Vz39+QmhvObBGasG7+rB8Yz3Km9WHq2yZegXjpNS4pwdIDpQ4XKaM949TRTW
L1t/A+g48POHioY4wlh92PhJA+mdGY7pTZ+N8UMKlxrHzzZ09dS9V3/mwQ8v4XhsKnPE1/pySFrj
GmT6pTq42xuwqkd19vy7XPJwqvGUNIl5yhJgnVL3hOpSGsJuBnecVorjoDSHTbyByCXNfUSaOuHU
FThXSTJFybDKEYX/UKoiNJ+RB5cnpEwpO1t60dPgqNe6jy4MagIKBv2eMQS46ndN2t/vzp14U4yH
7E3fYZT7WNYY/h/5GVdX471Ag3On+f+9qbg1Z80hSusIem8zxiUiq04LEZ5/Saqa6iPwu5r5vJB+
OGfHCiN49v6HUy9y1IIqQbKlHIdW++wWO0alxGKMUZDMZxPoI43wnCekIKNim0WndqSDPyGDVTK1
cVAcJbd20UkkZe8ZhoBSWz2EAIaaIeAhKO8tHvc1fXXe1aJe5l5YkCI9WKo60Br6D/zXwghBBqil
lSc2j3Has79uDlBLiaBiswXlWP9LL9r5yDe9hZMWC0BlacfbO5K9QAYnjmDLNm465tGYugS3eSc8
DVndVcfKf4J+CxGNj30jUKRjKs1Rw2xqrdLQE0I/3087giBt5sfMiqIjIVILbmsTiNsnGBwn8GZ0
HAmYTSLVbP3Zf5QmyAkAkLihUG3DYv4RIkiIlqRNomTENtf3e+G6eZp5seRGzblFgdkgFICkDtA7
yJTOEQCM/SKNKrQYiSymUGE4FanJpWAlrzby/0l/I/srNNK0NkslFDezQsnK9mcZELi7oIwctjhI
6+JMx62LtSsLjzf6AWD8Ulcs91+6lRebolMokYvQjkzxox8UCTtYufJhQa2xI5GpA0gRDrYNpiUo
bTbq9j7oAZizzJ9hgnSzdKHpQcf6Ao5ntPOGpUjglC0jzHYrIsoa3N5xsju7fJX/onWDjt8oZAB4
pX33i6m8YlJcxqJILjuZy8Td45WueUjp/eZfa/e7vFo7J3DBOQ6LETIufL0dbS5l/YXEIJ/pY/cT
f3UlzpkWD/6mCGRt/6Dbn1yhFJI2nSnAJZ1FM+qpSfCYZ6aqCy+SwtWD3NVSGEKaOMElIpaxAlQW
wE8OdR+nRGMtJW5IoSQf0JMlwlLhDrcVzaNnZY+BNpIysjMnoxd7Lj37ZoNuFS0pxlHaVr4/YV1S
oEq5V7xm32ITcQVsO9fVuz8wC7wJytVfuXegCMgahV7TUv4SKnZ0yFRwAS3NrCwguNvbOoPw2b63
C88wSxcA29ggWMpvTXI8J0DGn4qsl7LW5k0abotypJu5ZIb032YvlWtl+Q+lF1dwzP+wTpyRo8gq
jaTdzPW1I1hFGeVD9xuoJfxk29wgc/XTcBAMvvG3FR6xcXWXwuy2/fsu8VkVwY2McdcCOtv6XeKZ
sWYy7cvTWv0mqDkVaImQsoFjzhikBnYx9DrQT+k3ewK7Q4/yHSHwI1fH5sm6zlqXsuPmdyOJ1asa
uNhJwb0VSCkzO5sxvSILqK9dlWI1NlqN6JGhkMUja8xg2wU4M/Rxp8qrBwcM0Z8OBLgCk4f4QGyC
BSkFNYVvoPt/Vixwvxti4JC/KvMJ86+VS2CeMzvoiwYr3L40oCxStgOKEP8ON6kjdju1m3fRlbpl
ztJbmB1zsavBqnwHzuQNpodiQ79AgMgB4VHSctBCYPXwnGAninRC28vIhkAbiC5x3yjWsyJ3q8hL
wwcTgSSC1IchlnDWSjw6fXd2Z9Vu2GGWkqFYp3ed71NB+CRGgJ7UyliHrpKjsmmB2K6OTaGjhpNs
XhWwIIKCBfG11/rlyCSpwS1MPd4yJkXlRaBV2qJ02a2B1O3u07Ay5CFFkRQYI956WR1o1y3S7Kqg
9mabY8oQFUFcuTJlytGrePeprLmBReYUlIpuxh8+AqvUseeVZhTVLDmgVe3ep953fXdhBZwHfm+W
RWjY5MbkhbYv/dQutPqFw5UMbSwDNyU0DISRxloe8nlkAHK2P1ww6TlmvdHjh29wJ3hXmhfisCQO
H7xSLiAXOvy4+948M0CaR0jpDvF7RQUdr//lezhgbHWeDN8FwxBt/pO/C4MJ8a7o5tWdhyGoUZUW
MWItJNt91IcjOq6d32//nYaMeNagO3rQos9oIFCYrolWINUtXk4KGTXySZ91tcioW0n9ibxila8t
b2TjJu1pJjpd2a9tjq5H7QH32TsaNLxtseG9WNO4OBwEbosXeNZZ2gr0ISBRkzbb9yg8FAViEps+
TYKKukpVOZNiKbuH4EK54FW6v6jJKY06JAAkzoTBTNSzJQjShmwV+s4U02sJ4ysGapQGbNBURJ+P
Bbtt4F/in2PSG1C05nWUxsRieCzaZabTlDMh4SImdmg3pHwEGAcY3zwBBpRTmKys0uDeNAYEUfp8
gfhayACthjwS7TsNoVLfVTvKL9qSjcIYvd3w1g+zhEv6o0UXJQnmbc+sG2yAxu1c0m5BTl/rlmmG
WkHYWkQKd99B+yRa8Ge3Qw+tS6WH1TQxKS39X26A68B9FNdi2AcenOGOcnKz2OPIvpRHVX1raU+h
K41VApmA2MfwLC0jJr5itbWS6AEPO69SjpshBuQQdjrnMI3vnUw0M+n5Ml2RMHHXBXSPdHsuqSDj
jA+7yiq04b40EUXyzGZiuFCnqORSzCNlnz9r58Wy+ZnzDYCFnZ7IXRDitSUjvKjp8uKh57Kwoj/W
3qWtWTac04QbsSnuI17VmVUCz6u8W9sTRcK5k7z1wJVn+wbOh2427lJaNkEvmBzx4p3AOWdMNvpH
qlgyG5N+Z1+Xp/Z0xDnqErwVyU775NydlDV9nO8Pokd15tiq4KllXzX1+rkIFqvWZzIrsMxGxaxc
zKm61My7DkcBLA3KHnH9G3fK/2Cai4Kr2ofp4lbZt0Q88OH7SvFGs7LsUXw6dDvl8YfAizFEpBsn
lu1w4HoZeQjRDQjoO2YX/9YLHI1eLN+64dwjNdjNBu2kqPOOWN3HM2RJT0BNLCM/9nWgq/pPAjfi
xcGq58zisdthsJ8fUsX/1zfyqHOqF256ZJ0onllNEwGmFRnP1tO0HM7KaZlxEwf7wx+IsmTnaQfq
wLtVh+SPZCv134EjslUAa3M0Mj8f9GSsxmEp4eoVpIt9K7usf5R6rlqWxzm+GcPLjDtG6+Q8y+u4
NZxv1G9+JlyADjzKlDyY1/bt395iqllbmgnrxcenTg4seftA/HUubt2KmATjwndQ8ZGJkFO1K54t
83K9LsTFnDxOfGuyasn8r73cjgsz8df0kCcJJQ/Tl1HwhxLjNbZaQgoLwPJlcuVyMRjn3SO305zn
ypOXPe+cL+SsvMQPw4HLzMRG//nnLY8Du12SCNsV6lQUqIfznWN5iRLHamNgXtmuGEE8w5G7PToY
ogGjJ28XGFZO7kNk//gq31iC9zauLJXjq9bZF4A/jmXZmd7vWXiCEmwXEYf2MWwP7rB0p1g6m/Co
ajVoUd9lqkA6bkdfbO7yPV/tEKf1/SASHKOLWzD8rWxt4zxdM+YwUK503IFC7iJQMyqc3natQAP0
FGiN8f19OG447ypWhEaf5tByQbkBbNfHPQQPIXlGBbAQNg7ZDHWUB6pxKeCjy3aPLLZLLDgmsUjT
gc/vX7Ly/BLXb64qZgmt+zUTcvEfL1bhr0et24LkN9Q+DTWeEZ+CeSKGXtw38EIPUdDUA3l2Wnay
7oCWCyrR8ctxFZsdAnwBu4NuMNKujAY1SFZ2PqzHTNeVTTdgjcJQUQZhfhIDcjUPWQebecXhSzue
tqTPsZSEJ9UlHDQqPPqF2sGD6ZEY+qpxBx/satwznLsT44B0xObSrfE9DQT/zQqxgebjYl8buAGn
gG+RHeey6Me+ukBbTPrOYkFGJa6NUDwjudggy+NW3vGQKfm31YbPj/87raGkirrHaT3DUxabzhds
+Se15gusaO4AySKP+tQBaM9oLJT1lcW6GSEgLjlh17Ac8Gk4Pzu6KxUetuZEp2WhL/SzZ7hdeJ7D
ovRH142S1ZAeLas5IcoaEqNUVM654WPaZL0KXunWXVV96ELsSUuVbfOeoFFMRPCGBA5IhyS41pSr
MMnJ/mMlRvcox2j+J/otRm4dKebKYqoqqCdQtJ09s6dyE13jwBhbT2q3iOPdKw1KIvfxy1t3J+tK
IkHRoPpwTxhinxe0wS3kI7W3wTdfnw1I83h1KFdo9/PpXYa3aF/6QET3HP0qzIXsrU/FMwvZPIA5
OpaUbrCdiXwDUpeFoEnOUVPBQtTPZB1JQCKETu5eKi69BvxluyHYex4P9vGBa0lRumc/nzsE7eSS
vgvs8U/sw4Gf1NyIQ0sLByx1maHM+94OF/a6Q2/SXJbKYhK3qPaSePYxzC7OZd5j59Hy6b/yCfB+
NoiU3UJsfPCtn8I6k1L6eN7ukl3ATb7oUK3rUXxU55ky4pgxre6LDJPAQUhZdvyFIuOi/OsFgtU7
mz+iRqbV/s+WPtX9yGWzQ2fi3ugxfbFE8ANWp7lMBBTkHKGq/Y9BTQ8Q46BjWPBC324E5neNvHbG
q2kwATLlpo2lpeQJCvyXapFaAd1UwN9HlhbgIPfWhVDme0xca4PbMmWaAqW4wD0XgG0G+SKLwy0y
I7IjtWaBkrNXeTVyVOfLQMUDG0MGUCkW5QJNtHjAPX3yb7U2RgA+9laXsQMl+zvxi1aiomMdCG5I
o7PnQM7iDnnhGK/aZ3H6YpbP27KmYAbp6kFa+89dX40hEDWT7vg6sCEJbtipfIoEyVGXEzC+3X7B
eYj46ThFEGmIH6Ai6HjINChJGdB7Uw8AsnDz0q/56TbXoZ4T3lesEXqkz1mQ0+kHCTceL5V7T3pE
Amm9QAJ1lfy2FYAlCFAHKWhDL7QlmuLOGYs3AZLVug4gfLH/+AtlGDBvO202VCpIdUbnK7xMKCR/
MNbz6S1FmvIMMZSTviPM/7C7H5OQ0rp7dSdStSyG4BCLTej/JTNT8t7TDzexlzwkuHMqvjuPrjte
6oO4XsMLaGct6HZC2FamnyzjuZBEGnZWF4f4xLEMBL9jzMQDE+lrcR96ZUx0ahQzEndIn6esH9ho
k8uzuvbdbTda8URKdmtLJCtDm79pIjR+hqvl+OYsBOwy9IYLryLpCZ2RFAmaGAgJ6Bu8ZKlJoyWy
CRFT8QJJJSyKW7/A0KjIgFOrbQVFEZcFqIAWiaVQZEpoGyzy0GYVUwVWOFdxrFIpdQx+1veqj4QA
kSAQkggGR53TbdY42y4R2+gnJHdP+pQlx9N/5jnIuXh0FGGIkMan9psycm4nkcJPgG4Buv2xzK1A
4u5bJDQ303ZMib1pgVt2+kEa4U33EZplWUbkVoSW4p7Q8ux48MKiiCRfinqz4Vk0Et+vf9Tzgfb9
JwIU6tKjMtTYdtUk58U0l9Cdyi/ppbrIdVDIltAk/xCFcFIe0j3J3MQGlnHbMMP/6UwrJerF6X6O
sKOIUEyRa+q8tioaeZ8HoiPG195017vN3yKQihwITtnOccrd4/92ceNDrdM+Eym9p38h15XaOBhW
XiEfxOKJKm7KpQ+6Zm8um7A7BQhf5B2X2LxKh9pFfqdV1te/WP/jeFMI9ewoSmgTCu2r0P6MXSoR
wLcdGGT8iD6/tjaXHBelqZ9AQ1YYhAO49FS48BwZaCcgOZ8W3Hrv9QPDUhynX3fwearYJxVgfbWU
DegP9NClPpU4P4l5+5S1B/64RT1L230aa/DYIvwV8BFxL9uXvDw2dBzh73UYp/6TDP25Ka2bcwq8
6L/sxshKDjitoyIY3amiG6mB81qkZ4lN6/BQvo08374j+1/GmzAE1lWbe9Mj9ZMrGaTZIU8Uccd2
LTpV3OoJzmH53BmNfGFfExrk8/x7r7KmAlPWzCzV9WQYM1MC5kk+Y+aA9zbZu4i1TKhyahpjIYpt
C5KPy4uOgzKrOBCfJq01I+N+uP41k48nKFvQlUtO+DFjoL7Qpb+vPMzk4zU6yYTKGoJHhbkbstyG
XF4vWimz3Ggr4CYYearHlEswb6Y2OiyEyfwL8Rj9RyxvBIwrbO9Gc4xajGtXo7Mjishx5ALFvX2n
/l3tVDR9DgRGmpMSOtXJqaxa9nPyKlQkYb1ivosuy+EaittMHDe2fWlRVQLWQ5YViWA8F7NJjMQI
QN+3oPgQcQXJsrYVdKCQ0xoaH90BTatAYAYDCLVbO+V2DAOZXW3yRscWt0MlO1Fp/tv0ll7E6Iis
fMdJkWeKYYCLXye0jFsZqW2PzdiKzIhJ+0/RPx5u4KsKoSqQKxTSK0VniPYzvR8JrriP8M63ZUdZ
DqV464LhmolvziqpECFLLPyaGQs1R1ew7P4A9otxN/A5DuEiE036Srr+R3cuCDYeK2wfCzXHUCKe
jvPQCE3+rWtltK8t7EKfBCvRwkivq1qaQ2yqLmiOnczEMYgNsc4VZulF06/Jo5ZuRzgU6hAWmLKW
43My5Ql/4+/ftADfn0uHxTscBBwFbBFfU+GVQJqgogH79o2VDAg8mFvOXXlbbLtqBEAoLKT4DbyM
cyHhMasmOhIpsDcKjKrKVm7+TDBZbaPl644S13HjFhh51fVd9qX9oZGR4WQaTpARWMYmht0EohAC
jvFqnZBsDmfgh0gdMMoW4v+Z/lmPRrMsU3kX5fHE6kaDXff7JL7hX/H0zHv2pdTTJpiEvTLhRV+z
45FOpmldm2SvvK5fTTl3FItSDobnr9F+MUXEuOYNwngU5lNC0GFLAI2BL13U+8Kivzv8W5LZ7hjB
R21Fi0PpDAvgoi97oNkhU/Vv8F2SElQc0xtGdJAIsiXj/Y4Qz83Lg0NgOYQmfTHX7goEVdODyhlR
XmTOZszlHEFypAKNSBrjYge+7e1bl5ewB9m4GoGpUJAKa7a1hti25eQrjcO/c50NuXvsd92eAu/A
jsXguvLNixU6WGWsuSwb4XobbIStQbtO1IVdRYXAgtzNacbMGrvbV1xV8FA7wbJbH+9mnvcDYGMo
ln3FroAnFY4EIylH3n+YcBwL8tUpYgRqsRnB4Rp/dm7Pyw7qP3fpXRBqd0bXj5OYzbwYZIenKH2O
OsniuF+0AIkMFytZjBnfjT8IOIKPKp2tKVwRRuINMc2hNguG+ww++xVAQZ44jKhD38BHjM039p8j
bNvVp9uckh+a2GR2iRQCa3dQCK2vGnvlgG/HHVINvai+8KpiBETn8vwNVvcmQL9yKjnq4cfGOWik
D+gOQ0PpJoCafdX+Lnw/wNQEpQztfc0EOpB39xqDYwEitswcmZOg8gmE02JrvYufS3kSMklLxTvA
Gmt4ikYslO4rkvcM1eqTi0Rbhp+kjERNYRQfcyJXHsH6+jBWDoTBy2r8T7cbQEUWTqJ8ceS57pMT
F3qgiATur7oCjtVkn7TnOY+IVhWYZbQTvA7/m/YyUU4/oYHxC/u8pF7OhFjC9KxNJ2NHUN9k6f5o
LrFK2c0KTdxXRP7eu9nko+kOSKLBb0Ng3fddIwkj38VuCyXLzcVNa13aw+Rwe8tNNpEdFDu2YBUc
qe/ymHX1nuwZo8ijYp89Fds11/MVvxZZfzZYcVPIURq3a1xw1+GJb3wRijKjD1V/I2f1grU8uA/9
VZbadiaZnYy2zeDMdfFifeVly6NHVpBW9hjZss4UJyEHKAzY9brtCXuNNaE4GSdnYmsQk7M0JtVo
NK/FRedFg2Ssem4/DiC4R3P8h+o+CuHRSO23dlK5pLUxsfXTnRupkRlIsQn83rnJwvj3nbdH/fdq
JgSRXAMeoa2wBAXGZYEjxbB9kDec2qBxxhNnadxUC2kxSULwhjCwxXZMcRxnFOE+3YdRUz0IOuJH
vM2+aUZILz7gEY6ZVmYAdFHGLZ/9jSWuwHg7h0m92rY9hciZ4F/hz9EhFLhBdABjVMGPPVKT/x3O
whSxcQXtXO4WgNJUuYcdvtRc+JpK97B5FbJb5u3DnKYF2JmfuU1eXniA3YgAJkrmgJSl1e9p1v2r
WCQ72wwQCm/ZfEpSPVloBlYOgVeGGw2w7orsU+pvnFLu+Mu781sq0B5hXYFn716mHZVsAo2ZdBAU
D+cSFvyIG6GJfb5Vbur0C1QChLbA16kksNqyKMcAPRRnwddTXebAUv4vX06t/QbzL48/GbqejL9y
aeYJICke3GG6/9i/eQ+H1JS5WFo5vE67nrla39VYYnpj+s1eNv6Kg7dLW1IMIyELzRRt6MbErpkb
9Mny0RzWvVnfvye7t9ELQorrwe06tDLW7Q9xM2x7eea9c9lX5hV3yrSQHwIDYJ1KZ4a536IW6wpf
F/gP1US+Ri7qkYaKl7fVhx2kBx1cMIzI1EWBgmmYiCKVMve/da5tA34VtjLogCNrJprQh6/EQdB+
oqxCoKv7GTG0VHOhzqQxWKT/sE+mOXJn9fpspLKry+/ZabRovW07e4qgeLgy44Kb57XOk1+z4kC8
6qj49b5lc59WVti25LfYWiBMEIlZhRycD4YQh/yLAiQYdNibfkXJl+ygZkOLTgDcnCEJEI9XHsXX
0Ma4xsTj3fdp91Vh46gKSZ2+8jVrtK+fPPqJcs/COnFu1CZhUbsbZo1SVea4Q3bOytUpsYD+UrJ2
ok00P9s8ImdLxNX32sY+HrU0unYGJKbx4/F3aqQNQnvEAoZWZw0cdtGabhrC9rcB0Uhjq7ZSgZLm
SeqNUR7deY5McTgfFVwEzoka0dvzYGtb9p1qpE8OWHtlp/6PFYLE2kgz+J4NTkx1o8LEYa8FCTSq
/XO5yEXNw4QxtohvlFEfM08vuk32QIf/En+/QnwUWwofTyNhGwOvfnhNdSgYiljAQ56PUDIhHCef
QaIqGodCXoBzjk0aOjpYwNI0NhmZRxrlPOSzunVwa/fNsBY5VCnUaRoXmEhsfXROxwFlOW0tjnmR
hynO5vhROgeytPU2QnlQGsVvi8V3BvSzIqqqE5nFYd+KPBlYXt3Jmj8Fp4ZhRLfpjQHXZ3wG0P/b
snCO9grjWx0UGuZyz50icYCZZ4S3UdrW/lDgb9J02ZRB+A6xgNB6xem0eg5Prv1SWLDG8X0wv6na
oiVQZX2DP1N4H3bpapP/IDOtQBxL7bvHd2DAt8ykmA6DDsyUCOYWEnBBAJ/oBx1dFYKVdZRaeMj0
PxPLfPGB+GhGxfC55AIBhjqrloQwaVEbtDufCSmpvjh4UssPGgxvYPRjl7Q5oeYDaYcut7IFVQMt
xuKavf3j6sDd6CWYCN7AtYfew3IsTXQRDxXKgUNQ3GPE3U/dOXWuD4/pp+xyhBSNm2VPhbVSf0yB
38ryVyd5hSjqSxGrqT3je0o72xSdVZW1x+mWWfr/QzWyPz2rs5n+WL3DqQClAzAyNuxKzXMkATkz
8P00agCxHyYSd/gj6VzRJLuImNL433/QdUINrl9WJNltA/3rh36qwLliRJ6iCkhMQ3slE6OkMR0n
R/IrUkEqsb14FDF5NPpGg+dBs46xIfos2wdpMYNdnRu9CZC2c4FVJ1x/MhbVb3/pdWacRgod9UUh
hHzHOMTxss3k3cB9QFbUYhUTj5wJxHogrpx/CwwVRbZO7f31L6sscyzfqxyGmlZanlLk30et5+Hb
t1/xc+UfeSdCV2WirXuURF74q9h2r9mDF4TpLndqjo4mYHPcxXp2kE/eE7euNRQtSQHVWS3VhyyQ
4N4Jz20WSIqlTRqtTlya74bl4EkH/YwuglhUZn2Ifq8GumsRq8DIlLoNz1kO0Fu25DSNNu9vGAsO
kv8lDnBq8iRhTI045PC7KXMBovgVbeHtTo8bEwvnZteZ8EHJW0Jm40yfC8dvtVAU2kSIr5pllAeW
uxUqip2ivXhgCUL/ZnpLbJusWXmcikYFyL/AYvynyMlZRlYGKrSVzxc1eALIGBFTo0PGt+VP+UdE
EIRIt8bzVdhAwElLFkrPugYXJ9eCiN6Rp4EJg89Rlm8BOmzmM2mEEWLXsVf3wVn/LEyy8bb49lBH
59PbfRRPfg8rBmJglc8WwC+FeJ2h2KlgJYADEhJfm7uW4nk+teqj/7RBRO/S97I2nM52emQFhsdZ
bx+GuFAKHNzYtLWHwus5AhWe/hqHxtUd/gDRpFHoovCacRm6qH9jPv5ZcSjCYDkV1ITpSV9+N2wP
vBxKbrTkFSS+BnlyvHjP9Chqwtm30y1O+Y5zypC+ruZmd1hZJt3UI0i4F7IPQKjwndOdqQPPfqzY
TuGKwraexhMl9XseZnPnURyU8NyJGyQE3agL1oPJHt9KceLjAWrymJfOGTq0oZE8qZIyLxeg7Lb5
aRGwtdHKo5YVTEROlmIFAquTbHXKB41tKWz0R9RT/9Rs1J2WvkFaxtbV0lmm57yDTtOsVyswHhbf
9Xk79ZlGdE68hGW746A9DjbJGXWY9IFjbgNG5HzYA0uTLDvNbSR6lTAlMTJHvXMDKcekYvVm2ooH
ETyFWxKQ/TI91SQNUomfFhnaEaPV7VXPjuH8f3G+2sQeeDLXMk/2ZuvGMfwgiRAVS91fQVSDR7oh
izIZFs7eUefRbAzRDrQbp+TIVUcd5772MCv8avRuUjrLNvNuo5WFjf5Hp+J2+S2IP/MX+Gw2ZQ1V
ddjBS5c3SKJaJrgGi/BXE895geUo7OrL2FEbEkpD3M8m7vqMSqcDDIo/aF/KuxmemzigOe0X8G1m
N+A6XUgnRtp2Vb/A58l6I4s0+BdxrNos9/E+v5D0Uc1yOW7U+pKf1HpNdlZXV8Bm5/3XxBDXTACx
AAgTn74+QpZIcXjAYSfP1nQoYFQu6l97se0Doc6HfN2b3R8bwoZba0QjyYtXyohoKDnTNjthNZpu
vbpc6E4bVZLhjCJbd028EGaK2AzOsA2+HNNEpW2QIeJCBknQ95E16PwLUst/GGpOl9tPr0XuDy8k
u+R1b89/d2TP80Qxy0S2MxxUZXjF3sw6HjsAkaueDhMJq2UWgSPmneDEdK3gBup6D7GKlJvYZsg1
glh0t0AlzOx2JkbvPO3DYyMnrtbGXv73Wl6BBLr6SR5jScQlEkitcD4ZpmN0hP+XkncWQAnZJbu+
0GeH+RjcAFNXnwRlU6PVrGCVeyzI5ZeUf8qNQ9slSdZsxt9mpWKnU5gG2mdEVOxl0fi05o5Mr53L
DJaxi+2648InjFecQ2wd6mzyqa+I8zt2Zrre9TBJQRn7Uu8TGygrOaQo2P7pNEAA7zecuV4Dah66
2CbN6rhpu68buMdK0rwoKJoZS2o4oKYasStsEMwr407Vbml0mVcbQMIufbXz2JfSoCyDkImmJnGU
ggWyv59TgV+sxJ3Mc4S3GrDEg66X+qZeKOIAhwsyW7Sw4+PoNyYxjHrkAsBIFZfBids1ivMiGi1+
Gv8DxbULYC5zG90nqlB26rB1Lp6g1Alv2578nFlTNy1UJcy4/jUsGdIoBcVU0ZaZH3iC8krcbMcx
30pJcbbi6MxelGXA+kn+71RvU15cyiv1BkuHQS2V0z3o6WTuRd2B7L2FRe9jH697691VfCMNc42X
RcwE10crdfaVvLL3JWnbtk+tPyYZFTA7kIQ9gr+eZjNjqvT+lN9o1uDdoFpzJn+IXSIsNlryzmXu
IPBVSGt4njbc7z4CSY4HlMK4nsYxnf3dDftmgJBROYwlFAtmqwyH3jLr9AVZlD5y4RztlA66pUC4
UqGctAHAiopZaDb0kSHaK9AijRBUd6DrY6IwWpqWoYpMDEvJuNZ7Hv7VuDu7GjsdccvXQK+1GEUD
xnriBiuSegGIx7cGBp7ImH2Z8QO49U8hoVG+JGLDaHG6R4Jv+LfFa8E3rdoJ3XXtKvZZbXIiykap
BlW5JZREv0c3VBkoPR1FQLXPZnu8Khm2nlc7JuhQHQ/F77Gj0DHIqSsBOjn1HRECXQa4gB+qjL1W
Nq6IQsHMm1l6BIDkhnCBstlJdWvShCYnn06YJbJwGxksCTdAW+LuMVZdVtYKNiXixo38OPGfmOeh
eQtznbwbpgnL6u6FD0G8lX/2tq1gMJkSD6KhQ7J5zq3hYv8sGcYWaxUq7pN4klSZgbnbO+fstWky
kWFjdxpRuam2t/EL1Y7T4Z4lVagqglNuFX53hqHk+Tu+oyyK+L6SY5wWH6be8Gf/FQmwgBP2qKqk
R15TK7aCHbGEMF7lqCBgwFBQ+KVwPOxChpalIxivASZBMNc7hWCjq77PadlQOtR0r1wRR6szZqDY
vtOGq7bJ0VI+uvspjU1xAuKYW5kdxfMuG7N+u8wznA7uXEH81s3/Cp/vCzegb6yJ9b6BrNo2u+IT
q3yd6lZUhTZg6mM7MFz708AZDOeXDnxQQTMls3TfOm9kOadwbxBTwhdBW5kL7YiA6fpAA1mFIzeE
ELX6CPVrqFBNnX7N2CI6MTF9R5zONoCQEWKP5Cr7NUU/vTrXh3C0EwLa4zEIGpZdKf7m6AdvCJgT
+m4Gwwv/U2+uVkaOVCrGF+HwyIBtsWAXafAVftpapBmpYUQNgS8j/TkazXHCaHsz0ykIXztZNpzE
kSAxpUZAxFhWJ0vnhWUr9UHfFx8CZo7fiH2xJPTHw4K1PobCLBv9YaqrkNljTfDB+jC+SBeMo+HD
17ActqgMxnDQrx89FiCrFSr1AbKcZibipRDdezLJEukStzGXR3aC1xO9sqQODykmZ0gqEQ3loSMH
RJtRuAfOHkonpgsbCrH0h9se2EQKO6tegLQCQKKR9Vl22WcoSdH+eD/tlwIZsvY27MYFUB4BWAL5
PVtyT1Ff/6Z1wS7C1cfR21E9f6bBP/0L2uIHzFEprPIWc8w1j8Cws1EEXVrGRUZ1e7U0qizSFvli
JUXLbB0Xfoi7F1ll7tz7JTmKirAo+i4zrE7u+A48QuH4uw8F2cu2QejHb6UQvC5S2ZjEmnZQWZL/
HvFSMz4YsHvwMIeHzgKEDblfwTAkQQLnkkVvD82DWpxLp41BnSLWERc9/oRFtXTeL1fxke3ANxGM
7By8bx2/ZBJF889Yik0m/H76VF4uNF1wlRicv1fe+PlWfFKNx86n5LWdFAVqpWvD3YkVgpPPcpMV
fvV0hvltJzqAFw3Bl0BCe3qmEmIs9CMWg1mV8bUHQnECFgXfCk4p0N9Y5kKxAM0q07S4MtLn6abo
eNxscPq5k1SMGhizEa8pWT/zalO7W+4WyIAt7JGPjDyCzIZVSpufSdpuZUFAzFqFyeEbCZT4PDNl
N+8E92AIj/cKOwu7NSomUk1B2ptSLj2ng7pWNsGqH5htJkd5WSjCaFZYuyTGezCqiE+3aioGQ9gR
OJs4wrxz0ymZUBZ9BOESZcG9PFrccb0U6x2A9k1Ob2hAduHAiIXJN5KUCSnHZfQQok/WS6OYayN3
jP9idWRv3hoyYUY/zkg+6PlNLnZwO/vPQPyFMot1qmqZcEL/p7B5Xy1p+eAE26INPnUwB0/rLFLF
2nWQVy/gQ+0r5qQ7Wo/BJRob1U+JaVQRHlzu2qQFkHUVInkpNrOFXiPwxJrK39f58ybwjUyZUeSi
ZC9/X3OBj0s2y07zLWr2TDWWBIdfYLIXFgl8sjDdlkZgN4fNoHGC/kLQwuHd+k3MBQMyo7LYgRtc
A3Z/ZBryIslUIsnDRw/z2dXcD6sfZxP5B/Rylj23WGZ6IGsNxZ+HWs8j0BafRYuWPKnf5W/9mvjM
oYSBi3fKkJMeLD+qFr75H6I5DPZL4USs8rqFwAXOrsPcnyVsjrswoDUUg5oe9P/Z7We+EylCnk6n
gRfXVAXbVJXHu/ZKQb3yoOc0YJ0o6wXJ+dsEITyHrToNBpZWqWSehmliDl/+tbBKnIu8fkOex1rg
QI19r0YFFBPdacjsMiZfm864Sb+MQgsDi0uXLJL7rgLEt7ay908BbRTCJDuUez2xyiuytl+X+b6L
yvOSd2daEksTHMWRK7q+TZORNDCIIyt2WFbX5bHplIyWki5t/S3wUHT38zBOOXviWt83+x4je3Rf
V9jRTiD16Lz7xqQE8TWYvz1lqztMlg0GkIAnItmJ23LrzLS4EWbdOK2X1alCzYXbj+4qgY+0pXko
u8t7ZgJ36suZI+3GAReiPO/wvF/bTx/qCh+eAPWiyeoWslXT9nfAdod+AzykvjZBnkhz2+HFENVt
tV0dYQ6gG4q59Cj45VX2MbinQhZ02Emp0RWAQxAuIo75lcYBF65NVD7TFnX01TYn5nMox6qB97zc
TVzH2sQm6+byodF4xfUjYNiVliZwrhRj78SM7l6WaLpxpHCDwEIuDDrS+oLQngh1Ebo0eKbu2O3z
Ig6Cfdp5xIdDWz5JB3gA6qpE25gXuuTRwD7Z21gJPb5FjiCZaSq5Od5nO14fwVzmlK2rX2iR7/09
3QM5oykxapDf+F2lBxS9IrL9DwfrYG4ZmwmVveoS8V5seliB/Zyz1vtjU/Q/0gvy/WVrIKllh4L6
9yj585Tklf3DnTyEIL0YuMHQS8jeX1SS1nFkzaiT59Fnfh7GXcbSars2Ms+FQVd0YPQe7MlkYcn4
LpPiMm3lvrP+U69Q9No1htWDIrTTYqq97sk0so8ciPVzkymr4T/Vcc6+vcUuLNVLVQZFUZI2Y+8A
eE17g1sWNudnFXodMnrGw+I31ql36jlKoPPcREswT+UglXngKekc9f7C3zgIgChVU9uirLAOVR2F
klsLGEG+1KLY9NHjX4zhsWfoUSzH9UmIOa5iyvpJ34w4h9eik6F/S0xtZG9DWDAcFXTHz+PU2KLJ
LpCQ3Jj/ZklC5qHHGbRQ9qizIRR8uThsI0diQf3dsCmdPX/N6R0oqNS4hFntUDNWEcJ6qb+eQ0zV
7pvW+AQ1iaxGEyit4cEAgn7Le4WELIklZIefU26nS61Xy51Kh+O+HxOSpxtpQTTPDCBoF89TBlEb
MkFyWkmyuEwiFKPudukD43g8fOrST2EzI+ahxGS/NYwfmj8sTmxqI0QiaMfVWFYydQd9tQkyCIRP
+jmvMyp2m2pr5+h8smPEdoPRF/ls4vbGTtlCB/sapzasS5n0MWkNthqGngUGAMdWQ2efbykFHG3U
ZYoYpgLgJTg2pgK9BWYZ2Q4Q/wFPOHIMwiQHny6DSEuOya1dx7/KujJrpLcyYwbcV/my2tIAzHex
1vXpF3T8lmByvLM6+s0h9BlO1M0V/1GCv9bAMP/WDtRUD5yWZCQf9bqoYSG0X3FMjVt5jyEldiAR
OzstkXahpFdWsp1aOeUslBfSq/a12q9wN6DFMd22OMGec/1SL+GD7nr3dDpFiPsYkwHAmcUssVkD
twvnZjV30FXLUtnipb3RuXjGvVxDBWatJ2JoDcrZ1BXdHMuJVd+AKBy1cUtsQqVu3zWsDd0kvWOn
Sn64P8tOHgroYS4V6tcb1KASjd7B/W2VztEjtChLuoz427Jtwust1GQsgom1s7axvmCrKKvJh4Wt
EJ3pd3pvzQwMQJu/Hs4GFbwuWGmEd5YACdXbx8kb9/IxqhkGlN4xIcbhVahcGBA0UlM8KAsvwZJi
hpa5fnxZRqSHNTet16P76BAAEAHnaJRAlB6Klvfii2umttFeoheDUbFwKYG1i7p9j1O8HncaT6BT
YqcXGcTVXEBYzoFtpVVfqxWciJvseyNLb0CoPBFAqXd5WWid9R9ac1DGyI+9IgPcq9SmjbRZe880
mYgI066PWNEwA5UrfEFsSdRyEdozN+1GwqZmeWMSJxY7urKm7IZ+eAwN8GfxHk72Z8HG3JOi/6Aj
jmVDVa6yJGpIx4f/wxQwHToKGr59zUHgEFfvTRAgHhd4mCHh12zcIAZG1UtelxoSseT8mF1/DSRZ
h1KYO1dKHoBQ+a9bCdZp7GpfpyDvsW1QasiM8wJw1Cawd7n972/lA0ZDHk+gqy5j5ExkRzSpOlDD
5jgch6oTGO4dSbgJyH2YnYiilXWkQ8QNsFNvDBLQJhUxlc8H8Aft5JrXJftd3XxsdnYwy3FJ0xjk
0aHOvhkb9wY8FDoXTkOXT/eKUOFQXQCBKa9NRGbdHE2j+KFSmIFqtOb3hixKARIWt4nqoblEBxxO
pRPfV1gbg6Q9zCEsPZoV43K9otZo4r2ljFaAU80aLpvkoI+zVLcNAOOEJH8XzzLECXjpLakvukYX
iTsSLqHQMbUrO2DZJuPBy7gFatTL4a/sOkUh9dV+V38XqvQKLlkRJsb6MP5gdAeZPvnsqj0Ix2n3
RuU+HqxRCI4vkdlaegmjAJnfYoD0AO518mCNGLTVUwJUECkXzCKsFhMVvKXPBeBzgug0ZJYiP6I7
eHS/08UpIcO9T7uUGxQHQz2886qbTr4LTX+Hs55+1MYouvpnIPL2bXIBjaOAHNVhL8UjbRvfkE80
OybTwcB/BOya8dW5P0aYXgLWe5mHW3xJtvObsWysHFz19WTNPw8sIJ7U0uC++gmH5hVLgrBMj4rd
8+bJ4zlnjXA7j8nvxtpekAo6oKzSJecKH7sQwHAtqkgq8eSShdBXbAiBhzqP/BQG3nM2/FnRyrUu
ERO2oWpqQSIlNfCLoF/EfVb1IdaU9gcUWJGYxCz8Pu2ptxpUOiAFr16HzYLVD6vmLewNYijwt6Ol
BExbGnIVGR5Zq1NRnv6VKaMGOINIG5NcIO/TkzirAX5W49sB147K5XGtEOs0pFmId2bjvFij4tPq
U0XMWcXAH6mDLUiNd1V2/1zE80ln3tJW5qmDZO5hjLDMzOvwXhbL5+IxVewc4lrll575aQwo7foX
+ECUakoGFeNutQYPo4Y0VwOxNJP5ge3gaGT8LpFFoZTSkgpphyEwfJut+XRwZU8UW/1YxF0NeRUI
sMkWqG4NwnKXU+U9CWLHkQFngwpYobNwjRHYouVA/vo9n9HyX4RV+h8CYT1wkYBI3TaomwnlXdsS
bK74BIKWCzKzJ8Aue37/5IcUVpTbxTTR8GPdXz+GZHDdFEPRxkQmFjrTvibZbnF7vn7+S3KAoUpL
Fc5XWGJkDuxbgrO8knGjXn/iW0HpVDjc2Kb8d07R07RJCzQ/4CR/lm6d1A/OtiXZAagyPbwikgE5
/xg2NE9hJxjwgRKF/NkkeggKZgkEEJLfNdDAhXacPjSVzEl6jDVOV9U5MJtB31EK3O6KZ/EwY1oi
vCJJZmCplxXKyoVo7EMdSekNUtKC53pY0THxkC0cXmtuJ6Rk4/IjTHV7HKvjVsuPM4JA/0fnFyT4
3RMLJsB2QrE/WeRvb3mvEVIZq6gX98jBjY1OUM14hDnVd7g28SROJSJYn6OY9Uco2QAjJ+Jp3nlN
0oWuWOF8/SL1zVkhBYW1tHleOy+xc3lN9gl0RTYQoN1RG7HBY6DoC5JGxYElnTtADBrz+WsTv1Li
ZJRBr227iuq173+/8gy4rAbZSBeffBOdZmtC313k0ZZyQfROuStMMuUlOCdu2Rof7ipxngRSPjtS
bcSRcnBE94ykITN2UGgHsZhKSmUIV+iI7Y+GIPLcn6MYeaGwEniua0IEg6LMeI9mO5FqNZikWb5e
izVbRnmdMMX0z5BYhuvWp+9UVuVAIMYAqlycLqnGUON2ZIDwXXxHudT/Esu4w2H89U3pOvPjIsYn
/H8DoUPu+Zk3VOHiv37fEAaCfWjDqNaV7qsHQ0cajsAAMBGsgV9iVneRIQg1IpGPKxYG1qCW3zET
VZ+6Oa3zGg9cxr0paZVKFzM1X61HW3T0Tm5p9QgMNGFE4RudfiBydVwaged0XjGR4HfFovDbWVmy
wIXlHm2u0rti7RXWMCKdDSK1Yjm+iu8MuMIecXYwB9MFBCVaB0osw+VIX/jsGPKz1B+H/6a5Dypm
GrWH5+EBiSKW73gUOYTEyk1woP8TQL/PzVrX1vpjMRoJVgTK4AfLqyoXUtJFFGV+Aorxxw2rYcUR
S4IpyrBLJmacqrk6c/+9PEnEzXB8XiWzwR2OyvG44ItP/GXC+8VevgJLZ4UBGUtW3YyaORVkiyjt
El9AqJcV953irCMQaqN5qFGsaLJWW9wSZOvrhQb/wG1o9WCWFG2jPb4VhEKdvrAHPNj2ucKoyyBz
9zEiYfiQ3o73Cggm/TUpggSxixgri6lFVwcrccL7bH9GMhO2CPhBu4K08Va7y1dIzyX6uNOl0uec
88RtHWuQlXUsmnkG2QjQajTiBq3SuJdElqbK0ayVME7dZy7DJxUfcCShHFx0lrBsyGHS/GdggnWa
kas71mr4ejuRBK/HMicketN0s9SzIeBQvCKYoqOTiKEED8aSLswVkQSAKZ3yDtxldT6FA6oNtNBj
tXmi0kEltk1aBXxNI813SPa+hXfkoW1xGg/nBB26uxip+dqCz/AKBqv36efxZ6bdml5PvKrm7H/9
cHRB+7TsV84RC8jk96JlUej1A6fYx7epj7KZ7/jWIBZOLpvXabDb9HDq8N3MQmMilz6iDFCrMPSl
z0cK7lQC4p8uFsSO48oegTXIquR6q0hFGliQ2/co419cSbvD31tu2BZZJzu22QKOlbfMwoSyw3a0
gKKdQbg4TidMAN2L0WJkpDn9MhhTj8DGjDPV6cgLz4J7sdC8kMvXrQ52cZFLWL74HSMEjGbJATDq
uiWv/PNupEYa1Xan7/JmjWxC4Tx7wDbz0iX51+x9vd5LvnjRnvfqc2xrXy6YrsJRo52Er80VJVDB
oqhkq0xLN2Us6h3KneiaIHT4vh1O0RIJDLUYdDaHRE5lU3qPYoVGfc0KqsYsCbNz0sP7zYoc82XC
eKnu4nvynnnsA65mKjodcfUi7f9tpwFu3N+76skCb2RVhhyqL7dJ12ukqz0rCBmuDnVsr325jO2f
JNDlcGPTuoSMFqvWsNLkIxZ+h+MSYzxfsK/NQILev6QlnwRv1H94cmaW2fvw8ap9LZOxQMSnYT+E
lRk+Hh03sFwluHGCi1mcvkiulh7SNWxwIT8ppt5PwcodS2CCWv2oBylAIWPJ7A9lsUW3Y9FmIVXW
ZqB+y/pdpxfvt6YkfMAyf12RDBVrh5idmX6kC0K060ZuivnuYoL0ojVXCmyUIZ+qu4hmgyjNoWA/
wDjSGeZoEoJlHlZkajCQhUjej67ug3YajEOfszuXDrrsaiB7FbxA7GN6OmefgBcX2WkIwWGGJ25J
3CHMZfY37vuC1IjlEg3IuSfJIkRe74YZy+CVc9gVXbbJFi3JQ8/NOtyX2EaOBbJFdo0UzimBfJqB
o+GJFTU6O4bwE/8hupCVE2E5I0s70+PBwteBa/I5XLePwO92wlU+pbabzd22oqDuNyRNHbxFP6fT
ymalFx/nJO+Fh0JNhP+nCsKL6AmD431OHNEovgiONc4I+5FBDmUrF3SxSI61mAS/YZy9//utt1ud
TouJyydJSybJe40tup/vPARN81cB+V/6/j4M/Ipw0oQgWPYBK2aKikTdJEiW5W+SZB/8x4y0bqB1
bqqyqZXlgSR+t3jisVk21jQAyUIX3iuJGLLVQxfI8vXqsMI8n5C/Ndo+HUBT4ouB1Nz8lGbcibPW
x8rt3OQqnDiZbAKITDktNu0Hf15vN3DwVKy+rJxaRMV8c6Dp25WY9JUwTKx2J3ykv8Iz0394E2EF
FGrdMAfFTOTQjbu99U84v2dMQ4NvKK8/ty3oL0rLANalIjEU/BIw4K512CSGl0GNtCsDn1fCyd7/
Hy72P/1MnjiRUeRMAYg29M9t8TzTGYsf8DzaH8ei84LKXeHXk8zqbnGYpp9aq2E7ysA885P61zL9
gMPUPO/esZyABfbAfD1E9kUL30GZj5f9NLRqgnAJr7k7dH7Lo0bpyK/VYkPMjUTjpgdyy1Y2sF3Y
HHs/dQktpgkc8ZIqysRbBz0ABndfwgdfXn3VJy7uxF3UdJdStYhrOcwntXQvcHSW6q8O2t6j+7DE
dUlS8jd3kAxu2oTF7hwvd4Y22A0DjOJTcTxPuC9zhQTFBvH/rjNypnzu7oKaKYmBkhJI7AnayoNL
pjeSq98LfaRdpkNwl4KP/eVgjSQLWcOqLAFLs1TRwJRFlnV3YvNT6BSH6roJFgsJhNkyP4OS85Hh
FlJ+bLSCdklGXwRn40jrlxZloO7NOE0CBwGrrrEFO8SUrNcZ+qY6poybX9Wfego1DbZGWPT5Yit/
W+oRj509EM7f0/mQpewoKUi09ALwBh9QR8b/zOnVTHarHhCMqa6Xn/L6sP6uztB+EU7t+EkMgM3m
5nerJMTx+nglohpaJvMHsCBaL56576JfgVovgSPshT2H3rZfv6gZkogeqqitOlq658tMiN1zbQ2z
MwCs2mrf56zciMtKoBWoDRl992QRolqOMnpb8KbtujtjJedkSJIk5431oKn7UiTk6nQ1cSZWOgVt
n9AelKRQiZNp0wYbxsUUdjVepg+7Bl1KX68AwEpN24bzhhS7G/tGblOPUTBkaklz1vinNYyFEMPU
hEGNQVMKUSJ6mzcaI5qerKElgV8LlV1tcNRKNo3ZeTXZCNIHrJolWa0P89xvhyNtHi+/vLIPKKLa
3el864WQ07OoJUefW4057xCgNQvHtSrhsjBoHKsCg1bmwOjmEHnipbCdatR9YvGOxgCdoxt6WQ9i
YxpAhSuuGgX1xd6zw2VG9PCbxuX7/6gMoEC5bkvYEbHkjuzu1kJdvYnv+LHXIZjoQkvIj+iyS9l9
2QVWbSvr7I1nsAkU4tZkq9ssLrj6rK/wZyPBgdGnAKrwCuEOWLBMNzKZcoK2BdX82Xv/Buh3vClz
mllgxi8S39TYcQIh2i8llszK1Jb0VfsU0hK/B7FnmTtajxCL8gkAmj9hP+X2KEA602ewV8GFQpBN
4zB0+OLIUflVzqX3UZbRdJWrdmnH6HOPobcCdALbg4emxwkq2x1H04r/0bpL+nEe3sZvSARDncjm
ZjPh2TMJ3qGjmR/m/lZ15vjFaUPAdUnsNYPW6Hzk2CtO7K1V/nquzehXzUdTuxgbAxYXgPI8R/8+
cSF18sw9DuSbFOiybCl/7prL7ZjS5X17rdVm1m0GjWoQ+w2XfUrJvq7LpHeg74My5Q0Rkpqj9189
IjNaDbVwBmgwo8ARi4y6qFY4N9Hf8+CihbLKvgeT5FtSOEXdFFx8ww54NDQKku2vro2IHEK5uHnf
jQDEXZfJmonRa7vGJ6+U2kRVD7jtthBJT+Yue32d/6wbpTxbkSLAX0IP2dI9Phz9wONM4s467wGp
5fhdlmXpZnniR76eJNIR/90fqNy8igEvwkh/XB1KxAa0QUV84ITUKTZLecFVrhpQ3TsicOO2W75i
1/iXH7z0dMUTxKkN+bqfGiqsSIOy17d4QwCv3QHv3YptI37GjO3cW3EUe9NBA6X6qhZQAAGjIMhL
q5MAnlqhs/M+Iercjsk8ptVHq+dH3hdVRxAnd4WNPidyko/zHH+zASbPrWH+ObHiqHuBQz8O4+il
c0rgXmtCpOTJf0lnups6gSj2duNa9IyPbKyW46BTGXVE+5+JznHWQj+TaqKPozJPzB+9B+8eCnEH
656SEQ//MCxjCLD7HPEy/jZnqKMK/ja/qnbsM+elqcKUYHjBNnSt3/rNtI2cl+em7tISoNGgtEl7
tHf9HocdPxaEgWdKhMCV6pkngg2ebfOjEZqqZN9Iax8LbS1iIOylGb7xz5UFAKBojmtzUkuLnHnJ
4rflLjTnmBIw73xG3YPmWCXKvbaA7wLB9kHBzJ0EIkr49R0nD/cyzS6mRADW01xGo1LkNa/uRE9m
LTgEvQHc8FjiTrtwf8IhGFeoISiiOWckiNTiJg8NGaSEBnV1xx40fUuy8OTRIN2QVeCrbEihrIWJ
ck7056/aAQiRVnXiSHeX0hH9Wosj/OryiP2rZd3es9zv4pb3ThWyLGAGoOzAehlkaLF1CgQ7DmU8
GvTow8oP0A9xfEmFCU+jDFw46d6qsAmCWzs7aZV7C+dWOJxsBPch8TKN6wSJbabHW4sqHU8KlCo/
vd7yoD2YJJnk2ha9LKrD1cRO22aSq4lcy7NuO2YaiHwacJMvEdXbyWBcwj4WXPvswot1WpsS8QmZ
NVseogR18ez7N7dM5KTaF2fri0TxeDra7QMN7y6+F+aj0Ker8tdO8sEII5EwSp+o8Zjhne+t7yin
WeXGbnB6e1SaSDKnRxBNHbnPtUORmbrLIV8jKiU2pfQ8OQQTX+BrTJwBd2w6F1LyMZZD5cxeXy/B
vxqGxR4LWusXFCgu6bzAoIdoQ0riqzzqM4fX/4nUNjXibgIEDtiSuF9UUZu0XHv/bEogNd5OnK1v
DfHmZha2q9p5tGtbUGIR7Cayzsmgie8XcecloRPIDoD6bIH0MWXTrGWztKoaKvO0eBoEBSuE3aTt
M5CXZw7eLbzHuMQ94RWaUQTwiav6m2enH63xvl2em6b3jangqHVT2f/yfUrw829qdXtHPlhUFo5D
X2j8RvtgGpcbumKtoHbx+oj7hUDM4Mr/QWSL/ZozRenhbhFfz9hKbqCRe0XXp7D2EVSyr4tYFf7t
AYZ2xlk3p8kvr+aBqtS9NlYhukaSAnbUYTff9ajRm/+UyxCA+HsVnCTncs8LDyFdomlpwGPWPTup
+3i3QVGrDrSNc/8arS4zxza0rJ0ZhIe12UCPqmC3dq/wHq3DfAyPaVh2kPm4iebOAvp3yNDUF8QI
/9Hu5hBEX5Y/ApfZvOSlmwPgkN5PeTC+XbBtO2zff0rKB9pjMClTCcsKsUkm+UMRXbCdbKGpcUob
fSqEKv/mnV0VJ4rPAgLsVKwIFvkopjSY65wVcJWPH3kmPv3qeUkicKwOuQW9jFq3POgOdK6ymHG8
rZ9BeNTJI/INEg8EuFF5xs58CnkB9GFwEJWtuugWdthblBAW4x9R9ZQFZzXW2uM/Zot7JszQWpzI
Cvu4XAXtcUV+Djb5spoinSCLOzu/1GmWY5OYDTkxolexG87klbTGg99SCbQ4F6Q7KCDkL6U/y5ux
c+0hxV5XOHsvvGU/XdFe7mvpSRRb4QE5TdL5vCi8rw3u5+h+mp/4tlLijoi5E/dwjNIvH906bLZ/
0z5oykhZlt1uH8sFAF1gSpweCUZ3hjlrWjAb41kNqNPwl6c5cuGHGUbpGWrdU0GL848WQnbfhwSz
BNNoS9SYqEcvZA0FfjO8mKKV/avFWsaN5lv/qvqZzwIvcBDTxGuZyA63X6GPGEeZHMD4kVAdN19m
9B44CQfMqohacyBFja1UBWtB2hxtPPuS0H/9QOJk+HK3+v9r4ULmaJGhFd878UxJljLeVEfspILr
95vMdjiZGvbJXiwqA1ZhzxgaRaH5NBxjHSQDwFqu2/FnxeT0R2jaMr3qKkJg91p3zT96UAba7KEk
+6v6/bh4+i71OcUHZ68qQ94Lia3YzZL8R3uaIdHsNNY2eN0xmDVjQtEB7Hs0Qz2URrtyJgKeLnCw
IoNbRxI94NPZg6+VeQ5W6w3XkJvKn55jVnmj07UeYYpaEF9ORqv3QDTqk0OV0B8LJCRs83vikIiL
ct7D8ysgsnD1+UwReOjRqPDMosotre+f5KAuZgQpCwL4fO6ESeFr9Fp7I6UfjeSJkx4NhivFons2
wzXzhNJ+biPqTanS9seroj7ifrZr54owQNi/M6n1Y49Aw9UuYuUYt1Vvj7hMQyBHxpndj1WUxz0v
JMZ87/hrxtxObqVrd+SAqxnstyQ0tGmeqwR+Kd+OA0/9VdaDwfc70Asy1u58b3KmNJ6qy+CDm4/R
Vuqj9pjtAYtGUMG1vgrZyE2LdUgvnIsjEQbHj4jQG0rTmShalig9o/4mNJNXJvAstsPtgZWeCPE/
umCB6T4vjQGl860Aa+zmQ7YVKTm1vwrKd6lUHZMRZpd67MU9vecW2LSFn9JYKBuVgOMtAxh9i6By
Lhmd0IAA7BkAGAmbtJyAnukHunY+FjJsjqkZdmnwZWjRtVPGYis8ngAAoV49/AhDqMR8pCql2Nkp
odMmWW3Gox46yUoPqxlWDGVU3beDD5lGh7r6poFOENsGeRj/5swV0ECMPftsZ8zE9MW5sxMDiYk0
LyLzArbn+D+eMAeINtcYbgQOgLYLx5RYwnt/q1n6XWtrQWH00g6/aN8NR4SREsCxf2AGG0nt2GuD
B9P+qUbVWF9UzgV4y1rYOHMgGO9b5YhrvSpmtvom1/UoMbtH8tj6w1cXgcsDum0RJo5g17ITV/I6
mhqXznVpCSzUhq8cgYt5zwXT++eeSRKedxaloKtPnBx1czEOpLDLGgplnSMsPv/R1Nm2kq1UPJz+
i0JjllGI1EUWU20G6Y/9OH5XTN3U9dT1ATNIf0GuX0A88lPu/0gHvRh0g1Tbg82Ha/hI15JOuKA1
uDYDRpzwPfrhkK9L0iR9aK7nBNjrGZ32KhR/E/GC6V9RHNEF5rt5PC/hLNiUWGWD9Orbqywe0nPz
YaNcCgjzkVlSpod0EDF4r9AEnTQX8L44mu7hp+pt7ccaKsRhLIofIRGdAqgsfcERMH5XetaKBK38
HDvQWUgZAZMT//rf5cfEwp6CWa+4otJNS1HvJjqNnohtph/v3ESh9bJfp+jjrlfhHmCbUmsdeeak
1qyyjo9j7FQdGEmH0c4FfN1h9o1PWjA9P6biTAr/Efl9+tfAMbTAdQ09GRD0onSb84YeHq5tHVII
PLF50GwWw1VMjq77kk2Kd1WuMUFOsfd6pu6LeMhspzhpHBKrNFntJAotRaWJf8qSoUEH08XZDaL2
f15UeAqFhNy85I9aLl0kKlVVi7y1Kaiic0rwo38iOrAc58IpDoSkfGfPyREatxdn/iVrQ6nYfV1v
jFwrvGuTLJGYHQ6+Awoo/4S5BZdZdP7XZYv4yp7VX8+01DzCuQ+nbZIAku82WEOQ/UNu9x4buOo9
WfoMpThJxcs3tsbXrgyeWfqxj2lg+mA4QiJ1SuOxDx5xG+bdMqcLJ5DSsftWLhMrn+r5ouXwOSGJ
q2tthZjT/TKQX761Yw0Ux2t2t0jTuJ5Oer6DYt6zQ4Tj7BH4XZYnsWGZNuTqCJo5RTN9YBHRtwm8
BIWUoPoQovNf6XYmvLJdEj3Eh1Nb9FB6sbp7jeJtH/W/gUhb9HCGLjJttU+kZlDmez4NeQ2Gunfd
dzKoa7xhitV3jmV3gDVK4yR3PH8sozLKjYZAYaLjSv9JHvFpvj0OeRRZUJmqZ0I9COXm+FNxgCI1
9bAft0w29EWQr9Kx11w5b+rjaW7Xy7Gki2/4/czE9DbV0u15uiU5FkdWvddksDe1u3WYE7lwmNie
4i9+BEoGDUGgaJC/FlRULfJmjbP9zURE0sB9xq3nRA5zzQscC4f/OdqZ31Xf9wDYwoOaQGYHeSD/
NS2aTU6M4jFzR8MQUVIIP7N+i9jcHWW38yiPKFcH1Exp+FdDbftWVNw7np6tThxnefWv56c2QnT/
eiHI5C2Bc2AX6aiqtPSuBpsltQmDenW3GFlIOrJQK9ZuH4eRPXNcttPeqoBanPYdGnw69BMoFy+o
eYNk1mKFX5/opzjN47FxZhxVlq+2YVph76jv7ZMA0YiJSW5B5jmUe2iRl9xw7dFPvl700w0a0e+c
0InVweZTVnadOTzC+tTvwraFEe2ekmqF8BY1DEy3dTEEhZNXLkLBGLd8ziROgOXgQsSbeDCLAW3K
XhpBujczc5WnIyHZZlJseky1g0Vp/nvVSzA+J657hAAMTdtzW/ASthfaBkzHrGklTdIFm6Z9LNU9
XkNMECuaNO8VWkBS6LaPVpdXnhiqN870eY0ibacZUUWeLVjdIs7MQHdxXg35SahzV9d8E2/NhYaQ
PpIyThF1qQCtjvjKdMdJsbYMw3WCAtkSVyeBtfQayPhUVjNh32OviLSePB8GMIUCW8cvpP8+GtYo
eZ6a2lyeHvXqhhtsxOdjyNVerpVo/AGnMy79nSU5R0HAH915YqLkUX70800T1FIABLBvfn5C56PY
ej7UlQ1QKHdTFgvWSAA1+fn11jCDm1ffkN/xm8aiDiV9/9JjjctuuIqwQFZZXz3hgAjXs0RPC24q
uetrbuDVAPnKlwQ6l39UDEblOImzxffB3JM0k3+i5uMepmrmtlU2Yu4V3Z6RWq5x/UMZcSkZ3AIM
1B/aeng243ZEICjmiuIqz9QZfKOOMuf1sqxmWpHyUwIKU0hfhANHAUQirMzCQKa/TZffUyhPGsdY
7Bbf6Hwcj+XiyIJ+8ClLxHp8CbAHYqISg87MIvYI25hdtrablZZefSqeINN0QjNJVjXdtVDuvHJ9
iXM5MK6JYe7Q+R4/NzVKTIMwntBNUkg7wU7CppNKnbrqoXklM7PYHUL8k9lXIer9pYVeKl+GakrX
HkFeJ0uQLsMja5wAspK4W6EgEZJRjIGDgCg2RyeEvFaFRGvTGAAXXGWtHsB8RwYevAidmp1SMBcY
PHBRV+9Iv8TwOwzoCiY7QK10iYQe/7M1ATKDI5EE6TuKy3CNV7t+tc7wcm4fZztV5qx5fUE+Pceq
qnvyFqGozZ/oY/h1bfGZDRAsOu/g1hbKmp5nie5Kmshw98SU4Aq/mqV9I8lJb1sJwteL/H5CGEGT
Q5ePyU+Mzr6x5wAqchNhAe6nVzZC9IEmmk7inCHytZjJ4MI2/mOO/c6Ywv5epSaXzt3cEwt88nKo
xMJVV91bs3as19TP+K4YWLUx5RJj97wf1hB2jtP8IEln6FjjFO7OmPtNT81awEnYiGl4oDnaNKsM
EyajnvrMZLJKNMnlYKGqCtBBDfS/K1Y9dFiDKcDDh0a75ZoByx5SmcFLTMvpVzqt9OvPYqA0ZGlm
LsM82kXyOTaIs63QEQEgIqSafffDGUvZ6Qg2g3b3x1wQSCQDCntDxB6XRLuJlI2viw2UeLKtBkLU
vqTtnjfFEiXL1gVsZd6TbPoCb0Ng9uGkVvtJ/fxEImZcqGZz20Jgxz6HipSfMqpAcH41YXpzqNKV
b9YpVxQPe3bzXXafPW1IgCn0MXofWDzDV7w+e186m2sUAI7u9OtGtOX0FfU4c+OMGagr2a1vmdV8
7qpbVu0Zq801CIywWcErYA2QQwaeWAt3EkilTWPQI6J/piI9mkh2vVuZj6lBVxgaYhJ7amF9iPiF
fRzmUp/Fy6yWoFiDAzAmKmKMBMNfaF/MCV7/JkIIG/zfCBCeRqJk+LUTDgQJdYibckzxeZqU0ZIW
jyHceukxs0AvxPu7dVbyaHC9MaI8UA27XIXAJuFc6snCzkv7SXMPnJ7FWs5nOd6JDe9+QO2LP+en
1o/9MZCTVYR8FS4H1UZ4+hRjKgDiBRMALuJgNAXS/OUCWfVL0UfM6AUalvFxVpi+JHEI2os5Ik7R
VCrPELW44tl+LqkmDdF+DFAzam1xx+qAG6RVf0zsPPXq1ay65lD8LQIUtDgBxgGYOh/mJ14+U1kZ
GLJsIr0xeWCFEDpsXygm77ZlAk91yiOGkkdcROe/uIWzCmYKtxDed6L7pUEICnYZmiugYvQ18fqf
u2+emgJn9TCOLhFvsaajTczY40n+8VC5RVr4NA/JPaM+mwBczM1PbDHzCO1v4xZYC+vlzjKCrLka
VLwFhXKl2Gmlqxi8jrDINB6IMB/rYUSsXMOT01iaVoJzx1jiouWOwjIfc+FR1BbIyyJSNHnD2RWc
2jt2qSiHemeC8UGYfaIgfU5zEzkXpG4ei92Jq5Iez9+WWWgD+MuTEDSKBaOvlKXsMiG75YFWb1TA
vMBfrqE3QBv6D/pdzo5lRvX8Q0ayMp8qHYOBnxWVvDQw7L251JSp6DdHDelNizirfpY3f0yIpeMn
l4U4u0us3OZOaEcclFqRQVLPBJ+Q05hmLgZ18LZEjTzXpsbo+5vzOYgDbmadhpu6HP99nZWJPLUa
qAUDVcB6X7uCFo4krBZGEYXQkG77feo6xaF0uQRWSk7aaufeqo4uzpUFmDPwMqBnmgdi+6y43L0i
k/p498wooAQ/aj8WcsSzay1KWaSEPSP3pjC/y6lskLGrzySiM1aB7ClLq1R9JcqkSNsyeRMD8eIR
HBGZ6AKFiVxPxPqgnAzDaI81+NQbtqjDAsndH/Ee1cVHEPYnrd03yGpEofbKGcUvgR/oSb93t6GR
+jdqX/R7BFgiTGIS5I+BI4HdC3TsfEjwu6wdycdXAnfUJpMknecAqdEh8Ksa8vuXdqKKYdpP0NM+
V92Ask4hTo6u3Da+2LX707kd5qa4GEEOowfJUkLDXRbq18bvLUWRS79MnCizZYUpbpi6EfmPgbYT
XeMStgF4Cx5RwebQTbwuIhzUthiQ/imczWLOgCxLA7CZEH4wCVwFCIJSw07GZTPrlX6D+gaIosad
aijX5MNSqSFuTaTr2xBx6TJwLdQOu6cK1Gdjf0cT+d5yggqapV5ZIAMWikdXona3bCl9BOBLEJvo
3cDPFdc0YFPZxxlPcX0Rfp/y7r9fX3UY6kfyjAIxEDAinJGP/vX96OrMUsRniOwmbpDVGp9g8wb9
S6sZe0kHV5ey6LALdbv5htIMg6EuTR2vs5i0H4RMsDTnPX96f1HV6vPuFBSpbzKE1mQ7eL/gRBvn
8MI8ZJ76HjVrwXRRtfq/QonGIx7l3B/OnZUS5qdULj6Q/uDj9NhUptKFdt8r785dseAXFGBet+ga
Z1BKtEY6tBV5udzmQ/8s4y3bj7puF6CCniYZWxp1ciuaLJcKDj9pFuuFjdrFxwKOqvW2nmeUaOps
vu26RAwMMQIuz3JyDe1XErTyOV0O/EXHI36l7QVaD1HWgrG73oOPaFo3nkzxL6wsqPRkhAEfxOn6
lsTe+DgGqMtwXI2YMdga3bxmmXsyAEtU14ml4Rm2up3ZoNaNScAtHQ1QbeBLdewgg/Cy2wWh1XUz
FuKcrCBU5U3RqgEch03iBj1SjkL3d/4SCh3j/8j6GI726WesIzsAvr5qtkl2Mm1dj9ePw3gNw+5A
IGbvvzfHwrKuu4arSRvX6G82Fd3WtSVtgaqtQiACEdyU1eKIGKmltdOL/c6sPtQbcsCG+lCZgjfL
aisgv71Dwu9T/ncRzxiCPJVfUIW7OGJh9JATTe3YpFKtKw24g3h+h1PraULL33Y8nANtDicBoKfC
oBD58K7PDKU7uEmdOZxAAEML8qHC3mqtSsELR4kdKOE2kDMy1xZI0Bjs8CPMLczgSgdqFf0P11F6
WhKZtRcOV/o3MEWH+sdyIKOkWKZFckgh9G4DvQTx/ycR5oxmwnIIddheCmq+k51pOJwDqJSNxQuJ
gSlw2S6jEZ0PQXc2GMjc6FBXFq/3RiRZdQtJTRXUmd3SVYbUsQwiuTJBioW7RA2Yc4PCeQABm0PC
4gVx0vYgg2ZDIZ7M0Qw3550zMZjaBeCes1DUfJU2ck33gUZk4EuBQgBcI4Z5vdV/6jiYsmcoHv8q
8FSiu5fRFef/Gqsd+NfF4vIdkLRXbFH2DD4PNjOM8VuaY3zYj2qybpyiU+u49XbAuNhsbxINg026
TRd8+CKay5nsu4DC3HgYj44mQHLlWIofDCC4ypQMKfDEm4GbUm++nIXJmCqybEdsfNVe9VAyyz2f
2TaIy4URPShIohjhoC6TzOG+MesTfhR4u/yOcEL2HRFY6dlBvgKYiCCNyzQQ85/2pswOb6NmAaqg
yk3UsIHg8kUT2+pUO6evU+y/UDFHEtMqK+LZSvAJv0tJC+tC64q5P2bvDDqryq9uACwk+KdhRpfR
9A8agft13wgfYfnd+mVd4/1vMPywEJ6hJwx7cWbKGqjykaNm6hZkXssbBn3G5RKffWkDwyv7d7sp
Rtqm4QygyfPOW2Pq/iD5XE7Oo9aFYkgOr8Fxk09+qtNm38dQ5OKDG2scxRO8D0uTWNOIGci5ylEC
e6rChn+EgC3sXPJMIyyFOs1ziAPiIUr36TbIoVknJ4tjp3tr9bqNqp2SNQeLNZ9yygL/tDY3LZL5
pJBdt66pIjcikwjwcux6fkKHOaNGaFfSzxcG/WVadav4e5/Wf0i36fPrl/9GJMO4bd74RS+R+J8a
5FV+dvaTX/9fonp9io6bN/GoEfj3VbrPW8/XFwD2aiecMU8GSCrTuIKYSBkWQX8EnqdqABDCfMn4
eN89K/eTfT2Gwc5yZsB7MhPH0J+yp36nIPOjLPQYFRGnCXb34Q1cdKrPSG/65/QTnBrHR5LhqCU+
8w4v2SQyecaHZ7a0RwhiU67s6OL4Jtt6mSSsldISOr4VXtXc5gvapdTSwIu4nS485lA6lJZuEeeq
iefVpZ06EXrraF00iOqDMxCNyUgDCvffvSaPefZkuv7t23BovrjsL5H9rvzR7uNKjFeHqWrAap3s
wVCX4T3LzaUW68UtNNsdSWRO/3J5PBctfaq9PSYURH3WfNRz6wl1cF9SfUsJO545xcAoR6jW+9oA
ihWlHTrJ9e1JfDtp8E9R+oAa329xHmryDWk+qkK+vMa3TUI4tpl3lpp0EM9nWsWq6rd6jPrfrVDY
4eU98GEvD0ZpwGQMcUwrmOM8qfzrjBMje1vd/YT5fJxCdJXKzg20hKcBxywdJIGCwVInTlu/z/Ny
P63t87F0dcJLo/KLkdwBdmXHtxAYKxSA5+77t104Aul0mS+pKWLAYo9RKjLmc4xaapol9K/yPjMK
kwzvy4Fkvg2pRbIg0VSFLQnm11IEU85JSJ5T/hQyx9vaa62rzK0D+5CcFPYLnQvxIWOdSzGwZj96
4fux6bsv71tZfo3jW8PQdY6kU2FjqJCgI0jT8L1c25sU25LdrwpbTGFmNJ8lTnRtPPv6c6E+FVWl
Mpl7vkQFem3so88O60N22ABn8w0/B+1CJqCmDytSZd+/93d799nasj7TlgkkqOKy+/DrpmzpuMn6
vOeOWnSxasjtgGQLLRhfXGvHS42Mujigtdq+3a4EQzMgqTc7J+hb3VBHGCEp1ETI4pI7XGnvOJEN
Y0UfhGae/WZk4ELMhNu3yPpljLSnafSBLHwgSSX5ZMsn/7dpw82WMh7EkAWSzbt96eThpJVbvCVA
53pAqn3UuVaPdLdcavVHL1oJIx5yOvS11FLijjx3pjo1vJDiQ3K1P/OsCyFFC/FIFB0VNpO1pXC7
kfIXRD5CpBtdfZnlBpLsoD6s7qqrMQ3zrbVz/PR3gkLEN5IUrpYbk8M5PDlPUyw8w9dRfzaADyeQ
//+5ST19M7dFJObhUoVpPU0SD9s3uZssFFUcfez/7VcKv+TwLvTkSweY0m5wOOuRE5ACxveUfV/W
KwQc8FSKMpfXsBcBuplqDY2cscLCD3bAiB9yZZQoIqnNB99Yb8WVzb+Dj6/dczwuAa+Ay3PJd7Bq
Wtlmi+chHHau6Jq5oT9K0uCEtE44Z6c7zw5/z/N5kDWN9Bu+hoBB2M1wvWawxhFTRzRzAypRoXmK
7XusFpgcwqMGopaWy0ZuxkbHdALj9sNAOa8lGpa0ZGYl4QyiA0pMaX+CSigpcTLTqrDvsgVetdXy
AUp4MWk8EL4t0/flCj11ihAYYOBv8ryZ52DRRkreqjc8x9nNaRaRK6Ef5bGnnSK9Fs3cSlCzsoCg
2WwzpQwXLtZPHNLfbiHtEmuGQOnXIgVl+O4fIgB5Y7ijwTFk8QPgI9wr0x5p/Uj2MGF1efCiZ2eJ
N0OPtaUVHatjHEKnVILLsnvOxjCbsZDHAv+6dlBgXVyrAlXvJ8wUerSFWR00osSyxc/tysuVUjuo
s+anTHBU1wcpt9XbztXNX+SZfjfFJIzEgNageFtmBOLOnq30WL5YaD0eJ/ITvGuhdb04cUcCIC6A
Mu2/9oo4je9ImveD5JcgdDu9aQYWOyXVHncAsEPCAuzdv0bKaG43qHcMOBvAXTFGV9zxgs12np9D
+TX61lP/zlMfQ8H5RXysbkmH26iyiTR2XC8FLfWtvZA40pqz8OfJgBA8RJOIcAaYbuu2NVVavxDF
D4Vswv99N2Fxuk3n/GyMPYlo3pVTTDTDtOXVSE+K7lUfzkX5plh7TLCO+F6ucXaRKpzcpix74E6d
sXMQbvMIPvW0CXz5O/A8g7HEB6OIbSJubyGbTduB+1ITHGgWXZG6D2APhS+G0MgK/knkd8yadVMa
mAlzqZI7CaNylW7FGtfRLaCvLTyrcg9z9M/q1081w4QNdPvopOsxtdYRcxICAQ4+jj5VFL5RGxWN
GSciOudb86NLua2PxEJCc4Ja3j0jfapK+/KlnFUSoDIYS3lagmXZDG531Iii9I3PKfcunW9C9cJq
sSgNMb/RkNBXa2W1JdthlCN0TYP9F1Op5s9ff4vnjGtE/3uBZIrG92ZyIWGpGANnVHjkFBT+bc3p
if075vqWwgevtQ9kHqGuGV+VY4IxZ41/vGCxf0HSWxkpwQDZGeTtYBE/FFdCxE2MCRUgb2q7y4HK
g7aaZsk+BTRLqWukDLFXr1kDWrBdMQcEEVQ63zvz+UtZSxqLjiidIbf1lq1JXtdML5Gr4qQioQbM
5AQN4OXWkX8kjqWGr0scEz5XqQAWM8/k6Z5Cu4x0t+nHQ6/jMqPJrOVjqAEYmPLtubA+/YMZBouo
BvGdyUut3vop8ZMrF72v2WjgxaG3sRe6aVZMlJk8VQRWdaj+ZeNthvhav6VqNIv7HgBcahEAMkXd
vn8K0606YGBRPL3/Rab5xMkpBi1vmzlupZ53hueSr/QadFqsy4gtLg2WBikA5WCAyfTVGjgW+0uI
729jeAR1bk5lAUVRQ7Z6MmyDoCUbLxSLZ5MroTA7xQs7QhC1jGNzcCFT8m+aVMxHCwNVC+zUZyLG
j6PgCNd397oQ8z7gMJD1PGkFMaxF6tHJu1L3iTOLWBpii+EUgMNC5LUPG22u9ybbR4O/8FSppQ2u
HlZdj7Sv+lGmMC9JP7hKqMsija7vVqF2ykktXWcE4wkXNxRT9NwWt0mnTlTJ4Sb7nHcMsUyS2lbU
k3Fpl6dCpvRr1kK1kG/zj87My1cjeph+0Pj8fX4gXw6md8eGPeBVPWzD+KmMWDNH7eCRnrx9ecC9
FEOojr5ioXQ6LuDF+Hs2Iv1DOL6pPMMsNP10ZiMIUE5xlV4R03kd5jurS7FFnxSKn0nDtq1VSKSA
PotuxoT8I9QWdaDUB48C3AE/OVeN6erqlzV9vcgf5fSQ0TAU+FIVab8LJq5YyX0fJY14gm+a8cZb
OihDkQbqnt+iP7qVCEb7V49YEixattTnEQmaHxoQHEmIaf1M1fP5cYPNn/SE5PREv4HLbesyf1WG
D4SUDSB2dVwiHs0lxNnC3STvg1TAnNCMj+QtuXzdTLcARHed/m8D8m5zCVYXehnanrQAMz8Ortv/
8HXxahvm3cyDc5ccEyLkeX2EMN/wj6hnkQw/rawLEm4GsabAOmWIT+85EpSsjImI39dMZoaRBoel
4bK4fOLDSd2tyZyEY7jRgS64COtGDTc5/3Wzel7MsPzQJNPoUQvXKNVZzwBMrkur5smtCMatfHtX
iMN7+cDZCTNxFBEXSUevR6cFeKHdb9/OrKGVaRIgMgtJGFjFSqRP1nTqdvdE4W080eyUvu6Gspso
dFr2Zt93fqNTL9Nw7QqXrtQ88gpPilmWEH8masv4rdIdGEUAhaQjcPcweqbUfTGPCag4JhVJBmXN
vbsNOpPAxxKyusmtVBjIrL90O/zJdI08hguMvn4ARREr9A4xI8d3eDfMIxfYQUQ7TpK307gRc6T1
bwgjKfi1qDu+q7sa8pVHvunp3iE3UPcHrcvhroCbmOynnSkI0pWQ53tPGK8FCg0z9vfG7UjBaZIn
dDgDMxU6t1yz5SZrk0v4VD+nORZXcg4CSUwM4JAuae5H14sMd8GoX4EIJj0D1bbAfrnoqEOrFxJc
1rLGZ0lAFHNy+4H/0cMGZHm6NQkEZryzxQaD9B+R5fGQXBxBuTBl/Wa9A6nitHFt23ZEdlUMJExI
FJp4isEv3bmf5PbxtSUgAdi1CsUmUMuliutE++OAUwaj9junQZg1hPjVGdpftMrbCA63ZmSZfTvi
ytKtH7nVLfwYR6phie/rJQTPDPJZwqKURxws0NkoWs0LEGsUJ76tvVzl+YC5odfEHbn2kXiXxFpT
nCMRabIAFbkK6ecVcbWUp/bCEaH1HfNrzuMu4dZvecyc47JPKrSx6UbX3aj1+ncCzll9CBwsZiCS
+YQreZg9Zmd0OTpJBTAzviAmo5WMSUl3lvHGkz6dVxwRogrsS1bogG/DCCzgvM478I06oSU1Vksp
p47lyvEiSPF1/OdCWvfSyRjhQuEsMp0iJkbjKrehMNKI9QGrJXFJcKKyDaXAP8VXCofa9BNonW+H
mYkBHyJU/phHu/HlGPhPQ8MJvXWgc2hII6Yxupych7eKI6IA1+7MMUgFTuUXVv0h+y1pfgaJqEUD
j4CW0mUUiCa6tIr3xmYWnm1RBs/Jd6FwSPTBZTCg8hAPD9Iho9ylBLMWMMOlIfv0FPxAmn5cgLCb
0wUkDOMMugJrL9hRXwwKSdEM+j8oEXHOc7OZ727qtQeEmr0yqZBFHKwCDwfogxTIZ3ztk81dYJhR
g1l9dfK9zkdwclr3dDCWr0yTmwSPZmoOMzTjIF+S2jldyrOpgOA2Omfp11tDAHAfAKwMTjzF6btT
pDXu4/QLJwUJcY910aFLA6al9KBTvX1p24ibLI7nG2zoHWE2u92jy4FtHCQ4OZ4GD3fdUAakZZMp
SYpDHAPsgWZ00VKKwqDIYHXE+G1ZGzjMHpTbMWtZFGUwa7GT231zJXPc98EJIBPMZwiUPbrS1aNg
JJDBbpEDqAU5SdptZpB3Z2Kf01vDzaUPHqNWbOUrDuzQCamFpUzfq925pxyFwhUOanHZ3LueMazE
SVQEjM4KW0C1gwuikgrLoPAi+bA8tIuiL+4spIMCHhHTRsJfLJ1ysk32T6cptMozqJk2waAXwWat
AI2hkGy7G8ngnp6X+3DvEIcWu7ewlBqwXmdaKVX9cC4dKycqomzX+2vGVBFw4GXT/FPPE7+Ke8cN
+RJ6mdLVpS/F6Lbylj9bltYwA1QoWLMvFK2P2XuLoTKJQn7mJJYEGidJn9Ltc96oJxoeQPekuyGs
ZbnU3k0/Ytr5zRfhb4FaNz7lu5MVg0/EQ2Cvbw2M+Y0HeHb3O7NlfTMGz1hOlxpg51IpTH+OcTAN
EAPbF5pT+TOZ31v1Rb0H61vPAA/RdnHRZ1+pc12MxKqzOJ9yMmIRDTt0+IZ4wSw8GT3Oaj7Fqwy+
tTirOhgoCl8Ito29abT91modURWKrxD+QIhosjN8klj5TTalRc/H0t8fOPwEzDjPtfFKB9N/mVJ3
54tCIJ9QDwTlMnnBvx7ND7JclpAAlEluJrlXQ5YJ20lrHWoSEAhGL1VAvGjNT+2U0+8PoUiqasva
mHPZzXP7XBZetlpzZ8oWQ8aH7ZdcH0yh7YeUCH1uhAIPjFYPvg4i6aK7k/H/JcbMHHLe3z/QQ+rC
vz+JBiUpV6pPbhVNyKy26hrC4c8O1P868rSy5O3Ort3IEjO+6m7drih8BwPIjx84IjVKa4ptpoyb
l7UNEa0LNSKe/vHW5iklrErHwpD7a8ZM4HZGj+HUsC1GZd/axarBn+bFYEvoECJscHC7Us18B+DL
X/HPs15ADUkE0iHrhd8EmEtLpc5rHYyhgiKJH8wZ5OVys3CAsLRsat6UN/yk+eXQGXj4kOfddxKc
IK327xniGrJcKk9G7DhnuUdyHVRt/1F/SGCFxMWsAGDEuHioV0aPoe6EQ5tnoFuUDqtQr6pH+IZm
wbKbcFUBoz1NaCSIJ6PLJvj4dk8IwyrT8+NOZAoZp5plD/78MEYyUCcblLqw6vVm9j8070nKJ3AO
CE/RluZZE5WTE1EBdreALwhIReOj6ko2MnXiLlxEbBZk0CGKmP+U5RE8KtpEgQC5yFEcp2gqiMmD
DW/scjfE/xU1aGEJaTWg4O9LYSjzEcNtGOmAj5q9B21q0QdfVQsCZSRQdjhp5s+7WhbL8L9LNhHm
nkqMmcnEOAFx+ew6O0wX3PqWLviGp+lVzolMBe9JoVKDlaRE6o15QIsXMCqq3LJ0WzEI/z2YN5k9
VlVIAisQUv6MHkYpon6ZYQphmzAc8s9tuegXh66xhcdRp++R3lRmD7BQPbrh1kabjHwBm+YFn7Ew
CJs5zPMzLvWpxrkrPAV5gbZbFSurkuTgw484+fpvHblajYDRVFWSRUemxtnE7BFit73kTJbcIExz
bKGASvPtBqE9W8k/Ahg1sQ1+r2NNVGdBg3UUFXjVrLiVFAz1R1hClwd55JvR/nQGdNRSZS0DWWrU
qc/zRCGJf4NDjBZyhY9hxMulp7wnaKsKYjoigByWj5xAuZE7HaGZaTylD/3pFHKcQTb7NwwX/orN
ZthO5PcHtOUJ7nGygdkCTgmk1EXl5nsUF21iiBS+F7tSslh20Y5k7baX2Jzmj2cJos4EIMZEWvB0
nOdvDyJmIib+naGCT2qcWeyji0F12KTzfrf2SPoANsuPDu3wTAScQK8AXq59snNsauOGtbqO+2CH
xH2GPHUaHAFFW3hDO0FyZ1dIB2TZ3SxAVxKs9fizb4KOLLxpwL+h4Ol/xmCGhA63wLEwq/Qqh1YW
PXCfOJO+/slOs+Hl/pbU0jUXiSNeEH3EMzbXuCF+FkeqJS2e9KZYcIH4Kbivr0mZCv96XfLSo8Yv
caYXSXsOhoAhDZd23KJmkg7UT7IEYUio31ljy9jxeLZOyoV32kI3ZID4wgwzNYnXYFFaugM2Xz89
B2C8n2pJLMsT8ZdrSsVXkOJ+Ls1Dmk6XaFKDbOogsH+l4cbNoEJh4XLc7DQllLU0+NzeByx08utf
viBZkBl7WuFCZUSL+7baPzdJxNG+Ioy3mvrT2cAQLgJkg9WsRrH2J8Y7kM4SBr36q1GopcBYnuHG
549fqhbO69xsRCbjtL0MXWxk9mV3tayTmZmuFDCJJaKXUSjAfr8Cij2Zou1CFpEhRSsEKnuSWuBK
slZs3+fRiKplKiVgaoeRQpI8xqjbJHQeqbeNhAzoXcsveQ9qLWFvs4cVM3WLNQoXbm7sNMDm9/Sv
5KOk5lMNUikXR2Ch05g17NBBYpywE/k4xjGN3/bu5Sr4VCrA4z8fdI6ejlUYzpNrwDRvRUWbBENq
0Aod4eeIzbsfhgOhoURYVmQwKLd2duqxqhoCJy+ZOaNPzEGE/FCqL3tYPt95AQrx74EuFQNK60X6
I0L7m9iGNgQYHZvApZGFk+wlFPe3fU44AKFohK0D84/vdlkeNR+pyASPcx82U62MYcy3ErRsxwBd
xezLcwoC4aB7Uf1JznNUSy4KoG083Sw9nVSxp3hqQsnXd3wNorRAKZhM0f2zERPpWr5l9QYS+Ri3
+7+fhdXqLL4Mkhll/PoYw5Yhl0dpYutKXQqwylxbC/fsirkJmgRvoS7t5Zgpfca+4ARHLaAbNZNa
UfA7eZ+KdxlxDleu3OY/1b74vZlHOzMQzUH75yHoj9Law/4mgbjEJ15f+EFiox+Qtz8yUW6/pPjC
NO+v7jOsfVpCFeDnIbANGO/goRnmEO8CfRNLgD8ENgnrsVr2lPJ2AX03Onj56Fvj3Rb/VdqtmwGX
nUVBoUiwc0YQ5Mt0p/fJKDor5At2NQ2AY11DL8RilnxvXP12SX2W2fjv7alVU7k2M1g9g3+cuhh7
vRH9b2Y1+T9Xl3HpK/Vi9kigUhN87rq3J8PvtJGBqX7Up9abKEiSkYYxT45A31PHmjoFXPksU4m5
aZtbACX9P9QxI22/BkIgMVp7Nq1s2fGpXgJwTycxrd1M8qNTL1Bi5tLXsWG4nYjIE0yV8Hwf+51n
92zAMpijPcHmYs83gczDUZDByobGUYH+NQNC3uNnBb8ZREg4OjOx5QR17oy9mA9UDek5LeVwv/nn
HJYlOkWDfs8D6Pj7HkMUlXxxhF3IHxji7cd4nFhesRs51mW9JxThUEhNtVOZArupjcmAOnV8PT4b
okHiiXIcrsUH/XJmhVtU/pnn/MEwwoN6JiCmAo/fAUXmf906gwbbNbl2/Zpq0c+hFgzSuFGim1+q
PFWuqImbmvjJ0JFaNFqpwYLXUzvnEtSs/K57OV75g5I+PuTz5x8rsGbCBnu0cYNEjhaajFDzNr3l
6zvrReAAwtL/YkPc9AgnL8T6Xk8jexqH8I/jzHUksvpTu+H1I4+8dxEhnpUWfIfz9IO8z4vKkQ2B
A0CtOOymjaClG7bvKs6pCyHV3sYJgjfZRz8jZoBHWi77CXs46YWl0dxKwp3MWhXXrB98bAI7ZcrB
TErLO7MufFjo9o0ZkJauJftRINbwPfmY7dHQS/sVOcw4k4AcUoLxuc0ZzCczqrwz4jQ73wUBzVH+
/cBY0L3aRIxIbXf7GsdRy9Q3K97hNSKt0n1yRQnpQJ/yMkmHlssWAqFt+mRVMPQ7BmcFmHK48aWY
DO1Lc01hBgR/9K9KrSif6BcOOvsIB9JWApTKTK9EJpj9yMEBgxmeTc3LPPEDZt7biru2C5DHSheT
Gn2czkIwWkG8XYr1y/AAcXDNlCPp8mg67hp5DrRrQZQpugrYL5jsFu7x6QFqwKNBKwYrl92AkkII
L0JehT3puP5xerY3xfPTHRfk9QGjau7f//pE3seYfkN+qh9pZRVcnCFvpdyGmcl/G7Nbek1Y8Nkq
LoFL+FH4CXs1WvOE6yrtBc3Ys6bisHPXIXVUyy1xad2VRYZ62h1eGqG9hhuhr3FGrX75GuCGhPHu
p3upaTxH5pM/8XKmZN9Z9ENnJXoE3VaI6+aki7nG+Qsms4pgOIUJ9VpRaBfGNJY6jwnVvANwxb40
y6jkZbImwqZKJvVm8a8yjybTLeP1zsd8LsJuAzWg5+HZf5QXd5wl6sH66emgGPWBpQNik+O/rL/r
muNRhb2EzjWuWuBnbllXfnuOx1LUB0rzKtbi6EhQ0G3eONrbA+hSqSfCK89k+y/n8qq9z/24uELP
nmz6GA7iGzB4GtzqqFAf6Va803xFlGcu19NKWIQTbTap44fOzUoyffzImYToVIrItK+YBbbJs0Er
O8OEk5vdtTYnufeRLr6EoX7T+xwLr1lEuyMfHKm9WhIFWg6zjLytXUKYXMPBaRwap1NTO0g+PfE6
AWBpn9mfGOIX8SKukZaAFQGnpbc9wao4ryCSHNw5650zUH3Xl33k3kEbbe4ltipuK61ly0i6QuoN
0mjsC1MX1TgYwpgzK3XHdVx1ySjZ3zmra8RcWGj8EeqZ/N7Fy80wjRq/9vI21sH9wG/kgTITmp31
AALbhPl7ItJyiHtEp0hUoY6VvE6VxdyMgDfock/ZU0GHtJbikEnWIVlgq9bgXBD6D5L5TEVuvhoN
GGnO1H9+Bk+p7UGzefYoIyObzFnvf0sRAA3oFeUa+5oHjLWjuUlEfGtp507TI7NHeZIfx48iKvvK
cRjB340enry8IyTjpmY3DZxuyLBQUKgnOkqImod/tm6rFRXXvx2O7SYcs7rm9++LbXuAnT0S5Gsb
wEdzlYsk0mXWlIX+rTqU7yTfYBKp5QLhC6ytAIcDIx1Dzgwj/PDjEB9jlCxVi7bntWH3rMwA6PMu
T0x0kyPqRdvCk9OiONVrHiE3gm/HXYCGwYZyoGhGofe2k5PYBhl22p1A0UyRarN+Df7c5kNQA6J6
mrp8soTzCxmgWhSUOadoZ/QV7M0xb7Rllr6vIfRYObjnnQWlim0RrkVSqKF0JNIeKYl72H+VKIbR
M61yOrBvRKu//JIf7SQe7fLj5UpSTMkH+nCdz7lgY8/mckYoHtMPPF9DPcEq7MzTjplqmlaJe63m
nUWvHvXoRVfbgEqSAcjsv72tN8QB4Bn9LRR6m7fkuBeFdeCjLoNUvdIntocYmUZa+U6/kWYpsCee
KnTUTXkE9MLmbrTBdeeTG7DBpoXZddXKhfhPloiyKNAjTziK/SswGcDkfYwkSQeeiNnXCpFKvx57
pqGYn4MKrlejE2JFxxx2ZiIa2UwMmoUbdEXgYnEL3eV1GMlVbsse25MxyRhlSOWwd1LgJUcLBIia
8ADZSdY1pTcSKkjByS8fPMGvjngNV/S0np+6Yaf9fmQyQZYQgfUOwcMhYZXFESzF+amofAWWtV4v
0wey4OmCs9X1G+hy6zuNiAiOMTVtupE84BWSm9XalmPnRMrVNH47dNpyWj44cryeStSXu1MExPG1
q1QZaROv7EGFz7LGNabSZrdW17ToHFNQjKI4rCycVcqhZr/aThEQhDvN8Zk1kZ7AM8oB4bn39xIV
20clKN0rchj2Ha9J0DDFrgqoXNIpEf01sVuu+5c5qV3xH50yiOfeWCEH6KI1dy9RoJRBovxDE8i3
sboufQm8rOspjs3XBqwlYkDSaGRpbfV99gjYvy6a01eMzWBXHzXOE0UN2aW4EEYXnmDkOXtTmF0+
+H9AFw0AQ2tvF6RVOQKM55GIrL71NcCwcEItvdIcD0TMWqsVwiuqjDU73w0l4VQLltFY0uKzdfUs
jd2s3ICJyobEArD9ezknomwg76OJy1KEysxMHTqsoPZoX5frjmWhq7ImBrGjFEQBIRhDSIEUKAKb
UGXsix89I06rOzC49tbEcQr1eVxTulM+n4K6VXWMkbcmNDfro1EYBXTdv75XreTtgp1ebkNwXsx/
rI+5iJRRbQ8xTgAPx1oklzXtkVlsax/T0cNZ+DqSFa9uLPtkCmW4lLcO/3GMOkpAvNUEBRyutN0F
3uIJjZDd5Ep7KzUecNvVfQXPaBjHyZtUpDlXT+/4+dy7bTSJ5OMvZQLJ9C7OI6q7LlSbxhyjmTHD
Iaxp12FIPZ2O6lv0BMLyJHXnw6mHfs3NCLiVe+mWL5e/pGQhi0SYXP+MOxSpuUrn4hrGM+ZciXDp
OJeXipFRt5eqTmPyutYCa7JQjtGooWUX8A0LLGVRcgaMrBjT6WyNeeeRobAHaT4+m9Ou1n1GLcrH
xwcXupgsiztzhLGuDlG934vvPHYE8K0vwsusWUH+Ysfl3d2grp57PEAcAfU3fBFdiNH+Aa4FZOas
+SVY3Bmd9GpE33EMXDyhORRYvQpsG9w9jvd1lfruvTwwK766HlSSQTsitlqJkzZvyhBk4dPSxqaq
GIaLFEzQYykJtx8jPUUN6ZFqoGGIznB+crutFiu+qWvfkia2jLsBQaLfIw+Aw48OWVhjqLU3jzQ4
ov/VswrTg00TVNxGGWQAGJ5rNlOkkez5K8bYaF6a8KM8drgunLFD4n3+QJ0xP2Va5YTqaEYS1N2d
4aeKRXmTmUm+2DcoBRWoFjwaPLpdxl/Ivh+OZEFZyJLV76X0ACgV6qACDm2FNHsmSllPAID3BxSc
kNUpTLAaKZJhYtK9au4zYgdQrzwLwR7uVliHjWkOBoiwdOVIpseBbwwduxLVMUIv6LfjX+CfTzhz
gByv+rP02VenIkHUs0Cq79Annr44DkWkqLdBjoF7xNeg6PF7SEPqAI40BKkv0IOT7c9O2/V1wBIl
swLBsJ9vIa0LnfK/eN6GXKZexngizto0xcE/pYXe/XuylexPrvtTb0/UqpH4dgkl2mpLODehFSjP
G1eodvH4xUVoisN7ml2WoEj6bL4wQR0pEw4pBFFV89AvJOaqau/fekf1mNf9qzunNWAIlHQ8dlPd
8A7wOtuJPPHxF0HsIXIRAWGsK9c4mYazsxnHi1Hi3ZHiyHsv+F87el5c7MspjYYayhkBEjJy1WAj
c9a4KynB+heB1Jl5kaXL1/Iay4LaO1hOVxpo5jvY/XeXioIHx2hC+hLBIpOT6JFosXhjogRZkdPO
/d+UiHmyZwbB2B+K7HcUvXsK6D7IRvh/JPiSdAvUBuu4JyEUBaxwqz2qwQpPYSXp9+VtXLXbNhJc
FpE/R4ASxqC8ltvkK6RTfYJvp73WLKyxFuYpZHrx8DbqJSToQnr8Y8O38rS4B14Vc9uiDlNgT8/Z
hQukhyxLr17BILrQ/d9WRJFWgeR+LMHVd7EmvNyVSXSsgfVL+SqMiEy8bM8hvrkKSK7BQDQw8igF
5oJIYVRGRFl1H7+pE+2W46q7smvAYRzidS7j39/K6RCc8C/Th7h5LhjpC746nh0O78CZz+x/xCq1
rr5cRZS+px4WbTLhCcnfVxYiQ1tneDmEZZRThR/Ri04bd8pzCw6OyBem0wGGjBsjCHh79fZEByGL
TTChP0iSYjnb89qlp7VgwnYdK/rLEbtCSvBIfFDQEsw4Z3LHGfW4V6UYpFSKcx3BaaMwEqbGPVkn
V6+d4r4ZnXc+lFz2t0XsH8v2qWdq3HnsUDWvKjfcbdZA53Ubv+0GdLDZvShJZLOt6QN+c5MdlkbM
rEX+Ih6xNUHxsdEcagLQwwfHN4j2+s5OW2tIKtc7sLG/80V3AFmQn6HbEPX81RXZozNIAUbkMbzJ
qqRDxSi6h6sEWd7qld2ha1g5sZfPs+SwAGzimhkEZNM05k74xo17diOia9xFcnqswYshf/eaFIyF
1Ibl08qaFWY0QOajgKsW3y/KI++ySN9q57Drqzd/GKnrxLN9lO7BXvoo0JbQhM1l4/mPHw7gwXDV
i9D3hUFmznrPWGlF+Gfx2saH2rPQ+NHsRiXqhSfFM/Q6COfoESZ6nvg2ZuUH8996mehuPWd6Wqao
VWqdHiEW98RNLxDwGI70HbUJZyNQHQDTxyX9jxer/WajXrL+4F25JrLgohGl5aJOXlH36rxnXush
QVWTarFTbzxDyqfdaeP94r4O76l1Fv5Zdeqp2y/HKA8JhX/wTxoXV2Co50EdJoSZVtRIQOWhAA9i
2gh5Ne0rkWwTXESY+4p1EfmwQkE/zHBGAHGg+B9aon5XV5O+wLhL/S09iq9wVX6PL66+We/B/II9
X0Jg82Z8NFtuhZ2cQVhK56dmvei5ibUF37evwoRYkKei7dg6Ot9CBUbTBZpG7IjDvpzzTLhywXhP
LVgQynRw9T+cZyX3RYW2hKBBw5QV0SpN9fQ+81DlwNqXfVV0J97tCzz4ENbFtakzs1fqCZcK+u8p
9dGJwMahmJ05L0i/LLj6+nvDc6LHqq5sEdC6AB6LxltKiETPiWNSWTqlDR/13J/eBUN4G7AYa9dd
ZIFDkgzBaUH8Lhg2/CnOB3IobQsO+WGRxZJ03EbBYoGv4JNgnal1GWBA7FBctRp/3H6TGnGrhwIq
WVKEo8q3nCAM9b0Do7/YIyOhadyadZwQmDVHhGDbqp9S5XQRVM7ZlHmMqAWp8gyrfSXpqbSR/+7L
CWPcRE/jRvVBriK+7UxhL70ZlpabKSG7xxJsm4JXJHb6nvMe4+zgNUFpBgvAaHCqyjeG1C76q41X
+7Lv2frneqOpgeki48umRfbTAPDVaJQGbWhFu9G7zl+6qkPZl9hC5hoXap8j8eA2Rea7+3iEQeJP
/QNuCtIiWQoYJ90h2zV8vOhH3YF2yoBTj/jB+WGneyoNd+x3HLZ3jkr/QkgmQKYawLCzIrxbyG+S
F58JDS02TRwWxmk/iBqO6yhqX7l2xpgZTc8l9B0pJTiXxWdMAfNRR/1bcX6S+6ZB0RiSNxCI8Mwm
twYZHO893VMl/WPR45SUGI+/i7elXxkpu0WwP+Ws9YJCxFx7A7qAvjRCSRdXYOEAaR2ghq4wNn2j
hLSw5c5K2YjxPwKgMChztGXweFolQHP8E1M/RuHa4XmbXUpmgT25wRXqTIYd0oRXhTir5SDoeZwW
VKmdQEmoHauaeKV4W7PmCdC8cpMawMH6OyEky8yZ1No00yaB3YgeGq0+pcgeozsPzYkSPh4gtywC
DHxc4XYXBuk29/CEsiISSUYyVH/5A4eRdQnFDpuAFL5b5U5/3CfERtkJ6zS2+mvR0VLKRGW1AXwz
/YQ3t2YnRdMDkENJXOj6YplYVhElYutrJv4PNrJ1S8m9kC8Iorzg7088/ytD54oisagNXBGH/uLt
w9uvDhTWzIaAePuXmGyNzVecYkHUdduadjo3CJOHAPBh8b1YSAdoMYbRZEYH0FAMS3kW/ggO75wN
yQ+WFK/jan2ZgcVyIWi6L6Pz7R4XokQGNfya8cxIrF/QznPJl4eU7sP3NLuJRxAwCKZ9BtgSkZjb
h+yxtg7FfjGexciTzkKVX8Ki3gr49RQe/XQeqdRL+U728HmhE2N6jocyL59ixH7m+yntAam6TSGA
XugI/a/3Pu2fctp8d4qJmph52YYWg5sEdp8amHL0K+il4gkoQv8WLZeKhoUs061GNe47yGOjOpf9
+NWCRSdr/1VmKuLqcxUVe6sVLBjSFJXDQIwD+xJXH21+BhgvHBskYhQ1bPOM8l2aV6SFKhitX5WJ
F6agctk7r0VJIVWiGWQ6X8kyGMD3qVo4ljN2nB5QLxEgDpKqGnU7X4+pUy2mUVmLzfff1BsOxYyu
CBS8SCEhs/qXjWpDg6K/el7+fua6pt9C5OmTscFpShi0hV//HBP9SRs+q5CjGfV0IKcCRSNVnOyX
vEtjPE1B6WE6zxXle9Q7kFa5Qde9LWh+9fCf8d7ETUogBifC3MKjgKLm5hmgTsBj8vwZOGpdU3VL
ZEdqTIUYMEQEGQ8TwBiohNQDmcYH3R6QPgS+UOEJU9o82h41ZqD+04GJoBHL/GtIyYmceydS11F5
G7RiXYdNHZri9Ilucg6xCwsjvXmIcwVzLJD85NhpcFO17Xm/gnHBB7xRjYEsTr5acG2SrR+nx2MJ
N4P293D/3tngSgYADnu9sBnmfLye+3jr6cLtp4jGmJdWFonISBJ+lrTQ173nG1vcnOQRA2j5YtWS
+t3czIhj42le6Ntiq9gUmxGL+n+f2bVDKMJT6pl7uSc3uhVyE7OuGi2aTkp3QZxtqnYfw1h+kmr2
SFGzkkCJzkaVmHCx3onQ1Kn56ANPXdcQ6QOdsZI2NEkndvOV6+vhWglg/lh3q2SRUFQ8V6+SDMtc
x/6NeBv8dO8prd6ja7GIqv6efCsTbjIuUc1yHNQkvLxPVlpgpJc1w32uz5RKx4pr+g0ko0vuf5Nf
Ws+1O2aUirHo3DqCVKjvkE+aRfur0pbfpBeg6Edu1WMORcb6krSN2uBobO7t3hLYANZNU/GHn247
MBEO+Wf5B4AJwvGnph++/OFtOzT7b4eXJheaKuJjHqod3h6je4uUgZXGoAnhNO90WRlqq2WMfwl/
qAXbS9VB+BitEwYZumn9P6rasbbqWbXSetZoCBCIrSKgC3MBFrdjPW9vN/yzA5VERRtgNE+AkGut
PgrzBlqufmibeUCeTDNSRkPqEY/XmZdwWjvrdCQnraIOMGb6d7jXB1N9CstrwzrzG8OcpPMhcy5q
Znv3EMhU5hMgK3YWC8lh3UvutidgjjOHoyXNDYMFGYYgjRyjxWg/XtwlO12WDT9MWS3fODvwC3Oa
J1Lw+8l0Vtf+fAkRIy34F1+b67qoKMBSYJr32l45GHrX7VQdduHoencV3R6aQojnRad2KnVTIn2Y
0qz6K4jP7BpWu0ITipeJDd32WU6wK/jLeysgd/kicOcsg1mb4xOezucZq4Ye+NnAf3Y9t1u1EOln
BwB13zyeFnyxE3Sq4Uf9w4zau+JLukrMtM2sXK2+OBxgU0FQ+dHunYg80XYNJnda4CT8wHdcdCDG
c50PO+5Gvlx5WUDRWdqSg3eZkP8ON37RUqbPOrP2rUDPzyDBhwralkHzwCUv4erN8ZaREpVqejsD
8iXsVGA6z+HmFX1mWLo2w5mGL3d/74jB5bzF8r85/Y1icm8GKCumKzy09qiZswZsCIQNbT1fJSM4
EL2LiXlkfPxi925lA6OK9ePnYadatZGbBB5I7tyzUI6yONWr6Qp1RsJdDdxzJKgv/+Rro9eo3a/D
408d8SLsb6wIMxQ4qvZ7N7BbeS29snE8bi9WhpqZ2/99OL3v/5LCXFjv0EBCGuJndirFxi6e6uk7
gcSs3NGElKn7HDGyVZkmYCqWVcHbokA4fcyZqpJnrlef50DAww2FdK6vlCRUHbe808Z3hqtGSI7d
f/G1BCP7gUBTOReaz+zCPZmfBa+SkptGJZXC+8+3j7YLbpDFz2xb6QyGLnlDU3rvUdku5uhtHBw9
GoAZpfCpWw2upLWHoaX2Y6w08nyhFkRDUdOnXPTFLc4OTG92joXMoIYxQaCzxy3NI86JOa3cv9Iq
P7u6OFpY9ajX1Hu2XgUJngeD+eOq7l3RHGY03R7o87vSk/UZ8mOKFWJ2QizMJQgOeTY55edtKQC2
7jA+eVKHzVV+24qMqRK8cFzaoA4yMy1QddWsR7QiNgALzi6SOOMb5VJnPefMjoycyPo1ph16u7wi
MYzE7cD+TYkJMwiRSRnNYF/0zJyZ9tYm09WhSba3+o1Ij4RCs85O8KczgxEfcdu52oq6EuvcDBDX
RZo7V8BDE3/VImexzRcG1U+KTp9C2j08HEeHIdO003/RX69qKav57E7SXutRhgCLSPxMsg48zRw0
J7VOeqD28OYqi/LS/WMB3o9iU5fE8W7pS+wbIcGNgxHrbTne6bmjvA7lo6sMCgRfCkuOW6/DXSLq
4bfRypchBGfb5PqMVhxAMtTCDbYeYHMWtiZlTSh01goj0oeF/Ks2iYUBJet/eiSg3DSSgaJ+GUm0
9bw2jXqznh0l7ldML2Y/OJNcb2oFS3yZ+u9PJzRzjeNRTi3YL05WDwcO35D1orAVV+VI/PTWI3GW
1Tid2GjZTOGPc/SVYinIYQDwMjMbL5MIoDAvkKuJIj79QT5pazV6BFsYeoHL1PoBDTzBWMAk3r5+
fVxjlpVb5ICth/LHY51cyfQtH9HG6zAEfxlX0rauso2UGtG0mHwJI/UojkmsE0d3ZtrDshikJKwj
MW7UbRCMP18kX7t3C83F5afXkjf+8O6FkTBDYiUywl+0DGgplj8o+n2Lchl4pYlMYDCP+dlMNs5B
8BibZXs8o55PGP/djIAYZvGroyFI97Hg7UKP7/toJfmdJlDsDUgQ6jdmJh9I3J47rLi1lkCnwuGi
cCzapx03kyDEqe/SaQ9ND4NkylVBoCj58zClDBM8pw/EONajmguaBz8+JEZjOya4DelcV6EcIUrS
7k4NLllozt4Uo02Hb1gQc3YtRbYBcpjnxwXL2SWb+G3kNx5V0mGsDKDQtrwz3ZbUYm2vkU7vscBN
nKkLcvcIlyaYti0ZSU9xPZB8FzkEt5rt1BheinVIpOHig3G9Q87ZLsxtklH5Oszl4CsA9jLAMB5b
GkidXkzFH1OIdpYZbI9nnxEEBaNDthtucnhgNGMd3w8WP74QGtwxJUB4fNn0/FmU/GUzUAcWzcl3
gVqs+oTeOyomMRUmC0hvMGncUiqxymArXtJ8KjnabhpSphRt1Hm7kMv7N4uJxrCIaDc1vbGABkw1
M1jX1fqjht6AwwBYRhOYwlAlSygQ0SxPCkPPczd2ZVGKWX4Og3J9+OtfkcZk8t97l89kOlXtEgZ5
VcIMGp9J9s2LJwKzMBLnayV36Sltw6fqc+g/V8xPZaLuPU9eOTk4VcdmUC8WFch0/CNlUqes8fV8
1wzFTkgj2zYiTeGW4fd8XCxZdBLt1ZzQVTTqw8RN8vHDxYJNSAy6XDr/RKwJp8VMYjcmEkV56Y3v
GvVPPef8Z8a2auMvVfoYLISIHi4PYAzUEeerBai6RroEH82DF3tHkCLRtZZ2shykbTeaQW/Uf6Os
EXOskYrvGVFqvVkfWIfE/i4AgIi9fRT/ZvDN8uybZ+tJ/yYfPkbNObR9VT/loitiVxDNP6MK5aO0
99/QwV6RHIOR0d250pIJA3vs0MQPkRoqVRa7JApD33uvpZIw8vPXbSfuhPHgcQ+mdzoKDlYRVPIJ
cL0rcFnNm66Rnh2QHs2erkzUTeinvhkiISrkVMePxVnGrjJlTxOPtY0UNXdzy8Eyyzwv7GC3tp4S
E6ApGkkAupswUlUwhFYoRjXriseKCWj+STIeNGXvUR6O7SnYr1bmq0c7Q92He1sf4384Igyt3web
NVKdFk6au8vuy6aPTAj5nqtesfUB2NmOXAh7BHNu3kPdACV00x0xbb6LQsRveYBRcPtIS39nxVq4
velUmuzvodcmrBsQ9om9DB9ojYM0f6QDke9O1w1+bT9UDLYr1LVNC6SS8PT5jGlWf9YrlpEwBjbo
Aco46/IYZRvfGNdG/VpT/ecN9f03lyXxQQVl/kDwz+0+WxUXtH5++NgGK6OT1oIOqJs0wBDaw3AF
0J8CISFlejdvm4tT/dCylUrUoeiS3OMvjin7zWwd746BEHPX2SVwgctLBas/HsrVIfd1Ag5acy2n
q/KQ7wiyjB33LSs2q1D92K94qENYGu9u0Z4tm6J3+YiXaEVjPoCD00MRoRsB4H67jvVobO1CkGfv
D3wfAUCMrtFdYA8zVic5fZoYkaeEVmgESC93txrIWrUOrz0DVKoxwVob843g/+C0+8wMIcvfVgux
I/1Du3coquAFDZQIiF6IpJAEGk/QG20oBivBt6JpO2PPHR/ufvg0jpNaD98MuB+/jJPfT6i5Re8N
TXzrqK8OzamaMOBIIJHITmB20EAKDIHneTT2TO0/mo+4P0q/OjyzdoHRohFKzGKvdkJ4pb9sUd7o
amxbllraNneixLRAywawz8deIxM3SsP5O8OHHq0eBgMEayAZbkcBaWNKpCnOx03NWjE9/Oj5FpTQ
OQ4JYHtjhCl26KHGyIO9HP2NYh5PMXP4jCeA8LobIjytI8icg9TRENa2WA14koOqfLvCFEixveWl
1pyPNhOCrapMP+TRZCyuQY0ywl/RUsPEcZjaYPEkUkGqdKpG9frH7SNTJVHrCsbzxnsJdiyeFJnW
lg2BN4Ji+ssiCjfXAP2lR0UyXZGx3bCqLVwl74yZuldmxG95UodV7ooHwSPXwp5lktdZ93J8UfVk
wxEYFZ85ZTR1cLSw5R3DFpHkNsmwxsLPWhI8R5aIGawhf1GhOsGutGFrohhxxXpwRSjx5OH64AQ7
MEXmERMQBNFqHmaqtl6e8qbIe+2zl2c/XYqDJ9/iZc60QATLcRicHYi7zvKlJyE1ZIYIl0CgBNCN
fe+vI6wE/Kef3Zs9cGmFtOXx7NOGJuQiTOMwCGY9whmrkt4gDtPLV/lrNhXOJqCpWivzNdSCSbAU
pHomGgmNSJhH/e7uQll8qNeZmN1JzZEREjHkSiUl5aR2v1RmTjeP/zvKbcYUoHMsKl6vSstzMkxH
Q5ObNmdWODEK6OOrXddcYSVf/K1kRcYf+lvMxWzKyk2akKnemTNeySMzHLFsnqe//+ZbXggBuk30
WHlEQiuDU5Hqh9iXWjvoAjyOVwqrwrrmQy44XxnsZlcQh1iLquD+Qi6HWny4WuHvfpuPfGa2USHp
6hi4Ji3bglre3iXZ/bbMP91FBSm9MkLUkuwhoYIZRBF9xLJneilQiJVO36TcoHOAVlSMiuRgwZhR
k5q+dz2TIarxcBvCJ1awkU2qbxeB2KaL7ZBLScsu9DfXZZyOSlcHVPqqtVHByS2GkwJU4fX1/F1M
Z35oO6qA7QG8eLFu3wb2Mz4jBwyastUJv3nZgCAXVmiASw864nHKRwLOP9cJU3sOtUDK61rzZGAs
lntekHxBUxnVvgD8IcP9c8uryL+FJfL7kezqXFxftV8r43Ryt1BjXS9ZQcNCgiIP+RkT3jK3IM44
/njjURiRwDElFHtSJYLt2H73RQ7uBthHEwNbUETNMDkQbnphvWVtxFJ+LG6iSwtoxcpYvLXwlTXI
lzLmrNanAjBQcneZ1fTcIoWMaTb0wCTGMA9jkvqLQxIxEibgbqqyaV6RKv5U42djaHaJXwlq2qwG
JlOyBzBwwkwWPCukak/N4h+ZQG/Ty3s0QxE6LYtDTeQ55UnE2xrTqLy9sCxaFNG5NbTU/XVPD29A
V1oGSzv2h2sQL6eT9QXmzbrIU/ftUC42nxuTNwyjgrk7uIVD4reK2bfoogqh5PVGX2mjRg/G/MQs
NPNeaorJ2/fUh0lmjdLIOUQXRhRzDA7THPEOy/+txhFNo09QwxQ8M1NFEG3xC4y6yEufHPj5bxZj
HqSnNrQ7jidfpBMbLAtFn1t5acn6c1WEaUb7jg8Tj44a27JZ+HV5qeHuZe1CpTF4bqXI9xkdKgdJ
Kr2RYgmNrTV7HGloXyk53hKqQnFRAPCGdlfu6i1S7a2OX5ZINUdyR2IkPZ50IWfYIGk0eT5qIadI
2fo0bwNT4IOFqKpw4tcqHcG1KWAqWIEwXlNPuXPZuWWtFjwB7i+6+MPcvj+Ba//8e8aAhoW272lM
AWUyCP2Qbaj3xwYpnI6xmOfrJHITrHtqggMWUMcmcYMJu8vcWt0NPYW230u1eA5xgPnqiNIekIWq
BCXHXT9r5/Tya8nt+09cmmPKhjdJsVDGn2gFbvAGb8Q+dUG7/NrAFoKwu2DhtDPGKcnyc2QVTk9r
AZPXI1YnTuvW1/tfQgFKG7q5Bwy4NhhC7Aybmh9eTPDC2rpnrPc4GRTt0vfpBdRa6HRl4Kib/3PX
OClNLZoxlQIc16NP5ZMpdvxCiZj80NQ/qRN0QQR8PRxtdifPjBsEulT9hoqTYoI52H/jFFmR7a24
2iCiACUmBnmv7NyS/wJrJ2lYBYq1pw7G9MW3kRqX1HXWvrp2keHg53AofePl7PazJcD/BYKaVVUO
u+8AazzIl3gDKaQkELZ4GlMpk1okchdRT4hKcUeBjezjvgJzEQuyRrQhBC3wHoTd1xxGAsxnb9UL
8SnNGtr06CVyBfQVC0bGzAFSBH46FDGWg5WGj14IfunDb2rBHRbof0bnGAC1cqz6Tbr5lkGetHri
oD4xwUT9lT/5YHqM7BwAPig7WYI/I5l74xKMdJDJOSOw3ZogaU3qZmYaDfsyX+/r10uuIvWROQM5
1JCeS3RICMqNAjykIe0oYS2DYJti/lD7XD5hT/4xMYJ6QAq3ceDYsme8XLBBYv5GEEbyKa/afYCg
UIqlFVGr7Xl3WRF3MXvZTFB/FUmAM79yUsncS2eBTn0TLwA63zIWmbquZEfn/wQQmFpBKytJjR1H
1+ydWZKFKwmuAWOHD5ODMmZT5alRJ6e7l8MOWXcugKyBEPqYxKVtnbQb4Eyf/o79Oz62jHLkzlf6
J/TWEdU40IALtwUphgGX0xR6YZGq83RAWuN4p8zxaTfPtzrXLVCWidBaUEMYJQTBDfkNZor+FIGv
rOX/xpe3P25KGNwNMtQo8WK1SPHeOa5l4GYCVXbpUzfz/O0TedrWTP0YNNz1mKPRyYB0uYijFBYI
hjHLiV0mqhXCgkuZ/vOsDGOAWSSJ9C6SzXJc1WRnEH1kPL2DORb0XIxW2tArI8dEgEFr+qIlGIGs
ENOyjTXHtgr00gQSR55JMJNA+0eiAms6uYiTZ2lgCbIpG20hQ57zamz9eDfEUL5k/KOodrIbmiWf
xEIEo8lyGT102J1YWjBzwi1DMYgNI2SsLvXKjcoY2zp/UDVAcBZh80R67NvLfYi9TKYASgXXnNQN
YMeapL/+ae6u86fDn8A80XlwXuhaPwwe6aA5PFgm7MoxrlGC82aBsgd/kH75+3rmHsn/V1+aH2l2
REmrCSjtEuBG0a4GjO/NoNDAh/48FEJSWJLWrBdwbMxfkIr+wng9GpB8mZiwZvc9871r+qqhybtX
FFJ1lEvWTxuFqF8CfL4IB/hI0g3UvQVSdClVL5tO/YUPLhc99lFqVtAMoMcpiA7UqIU2jEWFzRWM
NRiQU7MuXXOgwJuazUtX//cOpXWFQa8ZWsm7+zayl3hck1ose7RMyRXXnnPc2Pmzto0MyqfuUoRd
oc4oKHmgPOxHYodZiV9aLO9OuYtCUzk76OE0QN+tkMFaMnxS/Ns0pZfTDc+e2ZNG9Wciw2R4cnQ1
4OLoa2act8Suj0HvNavdXElRrOkOICDwIPQ9tOV6jbYySSGHjrCU+ESX0WauEQLqLRNlViFB6UB8
oKmF3Ft1GIhV3HJ2Po/csl1ushI4bwJ8UO6MKf4I+Y+wID4P/0660fPRqqWgRu7mLeYHEn+XPLsk
XnUMu35EHxP6I566qMONFOPxKb+2xUhJo8c4F3HVr0YwaYi+eAi1tyo8a2G+psLwX3lGtBjpcol2
3YptP+h3tIZq7hxMdpJ71jGvylQeoG0yMMGbNNx0kWsVht+nrUGBncRj4RV91gVUgnPW1Z2SB5T+
9A//9HaNGQNLJ/mVA0fH3eREz+bNEu9gfYdcqAzs+Z9Zy2+4rFBBVz+ZFpi6F1FQFGt0bTF3cw2p
2JI4u8uCB0Wj2l578+vBJMVGs3Ko9TGa82b2Y+WNz6Dcp87lhSn6AyxOcJRi0P/aoxRk9xaY0jZ5
y30/FB7bkb+pkVwRB2tCxmjPAC5s4oHR/JQL80EzNRY3lP3zWW+NW0dHCpcZywS6yNBlFhZ1FJP0
LByjrsYeqc1farGHURUZ/CarHp+yAC5MDtGspXVPyKGeNNiZjk3C7hmCyJ2+J4JiBY34mCF4D6Rt
utlXf1+fiBJuQ7gtqXz/WrlmbXlkhYd2qhtFRcx9dQjh7n1FAIdsDEWocjLDySpmjhEYlBNQ1ojz
Jtk8vldVIPOtMp3zLyUV+/nTrev5/YurX9wnny+5yNETTY/WfxGZRc0wFAqY1bz0r1sJNElFOFvn
CzBbJvhBN+MTdKkgjeZ+3swWHmgkH2AV+3WBoKJ0cIH/gsUsi8ISqu/0ybQO2VMbR80gvzsdiPQe
q9DdDiOLnlGNn2rzTrBa6jJFtNplTncxKOAIHcyTqByuxIwqntbNnWpbOoo76D5yjNhseQ81C8eb
xohMv+/mORekFsOb3He0w5ovvRPuWjM5x/IFqlIp0kx0MZuwak0TX7eel64teDGCtEWzD7umUF+a
w3dvDvsNo94RulZZ0AkYitTUTKJHrkWNNjrG444Lhoc6IaypAHvp/4CO47dpdJI7+m9YrB8u1gXu
Znn1ZP3/2FK2gf4wOd+ikXWflQOAKOTGxdIk5JqgwWrsPisgHYm3+QZqOXoHI9t1mvRu0Moykrvd
EK9EiAOXp12/hIXxo1iGabT7m/WXuYYOUgJoh23+QXbvgVHwpUQ7MgumINHz6eANK/Y+RsZXXdBg
9zYNwlwHIcV4TzGQFPvabLDQcY/GFk2949zLrKyc3U/o/ibRYVuqxcmYDXnDPaW+I5sQAOL1ypAH
NSKhVULYH3u43+IunAsO0pWTxqx7ePnkqdgzFptLm9pb0rLlvG75RF/pANbeAJZLIWRxU/xQKsio
ojzkMaNZkthfQJjinspHwaFxajUJLZgynoJOClVAH4/u/igVN66tuTFHRXB/vNCbIpznzGUC/hzQ
c1dWvHdVYKugp8j3BSYHPDPk8TH4R32CZmSBYRj6A7uCR+tfkMn5MNRE+oerCCTvQusV/pRgitbz
5ESH/Cb8tDaxSQ7uCyX0D/C9vUPDIEoAawJwyg2QiGFB3eeLTx+BZ/hjCQmz/LRrS6QbjnI0Dcoj
V3wa03YwG7E5r6s2Fl8hRm1uQY6/ymMYR4KgeK+zquuHGadCSLK/9NevGqhq3D0JlvxUNevr7Goq
hb4bpAcHuW9lw3KJqcTQTcnXSt+wdtZ1ou817SYENxfTBJlOt4ZH9hjvE9PjSzIEBLmfVDdTgdNr
Eccvelc/fjW2/kZBlsa4HxuJwbMkMibA1ox8Jdw/PHzI8evq6xzn0IJBzN8AJA37KyDvwWyTzuTw
IIuxyykxvPpFVs2UfSNIFFPhCVdsM+CIsiuNOuTfuYqkSBygRuv3hn3YIgc+wLbheJENMWx/Q6rP
DMHdvYYt1roVxvU3NKwvHDijlmmoZ0OgYPjJjgnUsy6oaAGecwPRMv8MpKtu0T47VBp4CznaGGEE
Pv5weIfuiuf04ftihEfDE4kuUaRXCNbDkcJFcLf/r7RB01DQHU4gLn36eWeKy+VLH11VjFPYtQGI
ZqJhx062PaITyj1l5NOkZ017lUCqLj7gEZn0dknL34qRY2Z7+0f2koIpCL8NUk4GUY8kr4Zlu75w
s4rETPjpJc1R+APkQzxGk9HyHZdgoVGcSWfIJVTmAbtfaGdcF5i9g87dzyKhgZfH8f8XDAaO6463
Tz8YVPtgnPm4EethHTmhRTofBtsI3aIE/wUt5wKhO/Kr1pJA6S6xPFGeoFKIWoSPjGgwMDShOXbF
eeZ6xUBMwO1FmEf5PrqHi35TZ7DwatzDxYcFNc8NFOUuf+RIrWwWjjreku06RzzLC+mindSVqGJH
+UcLgMmo8kI92bVDpH/O606r2tC1ulVN6Uk5+kjSBMIS5GWRo2rLHNOE8HXLkJzuQ2tm1UCwRJt6
N+6C1UA12GMStBKxrNVMKtF1IKNvlON3uYeuqAUz0NOKSvTHPNWP2xYbJWP6NpJ4WqiP5TtXv35K
ZbWNcc3WgEZ0oB1JErsuOWhsucmpeZq8wpvfM4fgpzZy98huoEpBo4gOF/yUhs0hujzp1w1irRL5
HL6BRu/ZA270bSpFmAsjz2q1C0KBFKCU/ihz3u1o7Ho3Bnr1BtAr6Je+qvDTzYy2p4GUKwVMsT5G
vDHeaSm1GnwxwZtBUJ/5xAopILUsCB1NOKkNLwhetS4se/h74l7/CF1SocZfPP7vRALOrQP8bcoA
yEZcG9jT+6H1OUr/k+uyrbIlGE5lZ9CyMhch22eZVnkDi2hiOT01lYr816W4wOX5aP3LyPATqU+U
XmxkC0Y2eYz+4w5njW9f74D3ULzRxwwbCMRSBuecPpawwFoBk+ZxMJTelAoS5uyBqMQ5KajMyHlq
MRTnUxkl5G3cwGMHwmdHSo/nKpgedoHjb6h/M+4YD8w7Y4ze/KwpDMfliGhr+q9O240TN19cHqbu
5TzLKbwDWLnvXN/x2ERUAeDj9yBpv3s/mNh/T3Pu/gJVBdhxIMDpqU0kIlyEc5/ZXnrFKgsASU43
FTYv/zpLbUjq2Ibc6j2CPUo8BT9h0GYGD+qaYkeV1mmPePmjuzPWUNPFTUib92lz9XrWffnfdGkR
FT85lVonAetRDpjk+ZFhPAcsmrwq/Eud4Sw0qpU6CkLcHYa02raQJfuGCE8IqW53BBisM8KxBJRb
0k6HQXht9erqK8CF+DYEndaBpg2CvNlG+l+VCV/LvFK2XiOcs4yMaKy9zOpAH9fxRlFDPnILEESX
4GY/fA8swZbxzdwi4yQSRdnX5ArraXssCOgmdh8Htfh63jxM3jP7Jz03oW62+E/RPdiIeLv5PGd5
kvYwNi6QdQkF+Wqjgy2f8kgVlHTgWzpIdwWcYYhphrYzF/GQ9Q/Z26Oor/59NreObOmb5fVSYW97
8pDXGy05ftG6cArGgdyAL7TIJ4nFrAFaJ5NSQUHIjyuH1WwQ4jybp7asDLWeTDVh+NThaxA/uWCs
DTfvjZV41JbRFt7drRO4i5lY91G0JJhHKXybtejmTM9hgx48vSxxOxaJodjbymguijdkom0P6HAN
m5DkkZokC6KrBnNhCpUp68XgBbAsNjP+8WUYyXIO2qbQWPHlF4S+teC0+fX9tOmPjEqr4suj7bOp
zd/CI5a2jyIlXlzPk+hOktq5b59yk6YnyZmQN7guK7c3pYWd+eLVlBIIJep605JXER1Kusu/4Zsw
j7yij62lzmgUl7PIvs2QmNoCYBop5FgMc+N7wjze6EizF4OH8ozXd0WkTU4oI7Pv9Kfk9tuJQJ21
gKWZRUENEc7cDBysvw8P90s8M2ZcsoVks41XrYHDhrt9lRnLPalFjMfRKGXKR6shvrINHX8o7eqP
Kx9ofIhqFCpKAWltSuTAbe4qybA8kvlemRY8JuWzNyTgevcgG1igLzLstzPyO380pZxX7G+bjHLp
6rxolpBNbwyFtma+XoZv4ZEyMJqyR17qMDpPo2+5jiKPSr3h36+Y3HT2P7+bFhRZ1lb+eLo7JVBm
sPPTV56g4wtCdva74tU2IqFpBtjXa2/VnDVfzK51zu+tOUFF6YUmwpeE1fjPo5egXIuLFIFVRE7x
Lr8xjRBIPXfqn2EMmpiGulokqX+IMhVqoXsq8U6277LLuBaUESoFaDrGACYYE0jmEmmwYBMbGDu7
9jZlcj7VZVCVl7Dfnu+OIRDf5OHhDo5vv8klvBWyGqnHRi10o2qFiyK0BrAYwO0GzzcFLWtdetln
r+vJ0ved6XxC5HTRanuQyM4LMhhf8OZcGAZp8Jvno249OPgeB/2ThUPdfJuzhxNL6hz+NA2ban9n
BgeBvqKldg4OR3VcUUmBM8rVjDG/4qlitMTxRW9km7k1KReERArJc6G3UaKCc4bC5TzNvA0enIbI
+FXL/LmhDLPzGblYOd7bsGSYuCkaQcv+fVSg68ZpIFMB0Q/f+7ydxA2eLThoj2sp11KaTL1gZSPB
f2aiVJPZlPguslyKCCVCAw8RlP5XJqA6NL8azKbNUbs3Qo2okfZ+v0fJ1bmPPUKwcQPzwXSqU+FN
4hn/FaOZBpTor3HfUAjnS1SxwrfyZJFxPsttXmYQlHEBJb3ngMWKkHNqxpAHCHHCklkT6wdU67+o
l301Avkz/3AFCpd4hR3mwg3WtPBaKPWERx1FhbVQWXCNsIJA/ngcNi3XIkq+nLEI9XUlXAmPWGn1
CxCoQQzZtLx2dSABV086n4f4CMS1pOnfDqV9TYh8+iOJ7yGgTwWZ2M/kW3JSyMHQ9bIow/nqRzYN
r4jup+NoQSRoTc5D2l+CcVlipHZI5HBto4+gwAMR7sNGFCL8hlJSFxd5Pwxxzugmnmnx5fxUAh1G
Z8ppjjkDwdG8f81DKp2cCWl9q0OTGq7YZhIXnGVhB1V2zVnThFiKEncvLIdw8ry99xWhCIp3169J
4J3vr1JMiOdOEe00T1ag7tg91FgUrDoqIt0lBZGqIO/1gM8r2IqBNmj6aqQ+ee5Lp4p5e9aR/009
m7H9vv+1hy7i2qLQj3Lg7SURitN0tONu8ElSJVQHFXk9FqZWp4x0VJw6cUV1REL7VAeQhu95nK3R
z5VsqWY3XCiL+/Kn5lXm3NgnNtLxK7A3yftlXWfRsOaosscAhE7gi/Pjg4GtLVvCXjmPk3iIP4ca
Q0XXfKPzAtFlONTMhLS1pNvBVgjg8tzPpJIqaNxGlPCbHrKwzh6ob1kACXcUxZZZvw5uiLNxPRg4
/blb7FrIch7QrHYZ7ZRwG/eYJfwYqDQNvoc/lKOm1uVq+C27YO+i0JZiQARSQ5sBCqFE9g7cH0oX
HitBbsJlw0KnMvYQiTDrlZORZ1gWYZ/xjTzOWEMc8bi+ndZy5i8vwSyIgPaR5eUNHVJnSpbeCRz1
cNlKTiftoaawIchwLt6ethMzfWgf3K3cYJv//C/ObXA4Me5rKbRkChzu7XMBAxAc5vqv/fU03CaE
I0BuD/nuAIiC/syngqRstEaQnkLCETs1hqP9syPspqU9Y8mer7lr8e2j4QySkOqbcqCPI0nv7q0Y
+5CFDq5n6jMj8Im0fESHY45T1RoXMra3P9YwoOh032KWElQfSTNdZ1xGGxHEdWafelSHG8BmOspj
u/KbLu2L2OFNGSakDLRy5vTVu2psMI23WnsfLNXHnwNOHYHwIDVrqFe2DVSoFYn0UGZANqhhtU8I
VYXc9s0huTRA4G3NRgOZxF9a1f1iaY9Wkmpqvp1l8tu5Uq050ZQ/kB+XxBtPn6uHDBrWsOutky09
+IBERy7mKnQCkvYthfZ4md6KOuROa6kvGHENoWNPGcbmNQFtk2Uo2p/Fl0lUnYfqycdlDUpHZHu9
vOCpC7aEIPIESQhGEX7wH+UkEawL/kzz21WsZjXOkLQbT0wHRC8qRWi2CbwkbBMWKgIQ0t1IxCxU
haD1OaZlorPx6i/fr/sd3JPGLxkR8LVAkdNcocXyYP296e/Kfe9n82LU8IqpQ5Q2TKXLbQBYwWcG
PArH36GjIL8r8ZyglxEzd8VdTygCwG6hn0HHPDAu2ora8HPATA724y0unKk/WpMQz6t8ZMaHzcXL
ciqChwjKiR8/wf0ikBDVZ/eMDA4Xj96HTvWHc57zNjOkXpadXiDA4tKS3OZNLdECMSRW02KUQmKU
l+oWUwl9pmO1r3pWJyZH+NKLX/NmS9NemiDl243PF5HKGgGFJVv6ilJCzuxTdMzzEsBblIUJN61e
hGm/+O4yrQlWVzbMwuuHT9PcsFCqC7j3ZMKoMkeH+/xWE9NowleE6msXchb+ycg3NsCH0vVjt67P
pItUV7uifFyQBg2e3PHgnv5ZokAwvjid5ugaOIKXexuTycRCiP+fXv+gpME9cSk97aG1Gum07yf7
x/Z3UApt5aw7sM1WQOWb7/YiGrVBBJxZfPQQdIhcey3yOPEyQK1swGFH7Tdgi1tHtjnkH/fwWEZr
/Pj4gQvaHGhlmC+MsvIFqE582dnRfs+uMP9ql5LwUq4z+dGvG1nXXxS4EfyOHdv6OHR8ZYQ9RdXU
VdSfFSc8dWHC/JInCfrVFGRmKBUV4dG2Taix4xdcV5SpPysA0baMOSbI8AqMC29HMqJUhJItgq5D
qUd07155NFFRDMjLUPdIcCOj1JwcgyTIPFjMCr2ykdy2sXd1Wi8xK7DE7c90EiDVzD0xeyt/nXkT
Dr/pH7NBqjwA+NDe73rJobAf12jfdJR56mBLieN4RcTjd+l2fnFSazCz3F00ROex2D1k3knXbyOi
xTpbxgz8Fgq3um8mS6nciTZNkEY0e8vpMw8dhvAhJPVyxKMA8KCasewpBny8etGAlzdqIXBqciDB
CUIiCgTMPTDbDrLydn+07OaZKFnPX9d1O9PtztVBHMkpPbWdYp6QXRYmGjC6sINRRCZk5oyIAHP9
wPxQNo8KF80mnOzS4W3rVHOW8/xR/YTVybzpF8VsFJYvZA0VZVo1RWS7PKlJjyDwsHjmzKjRmWay
i65RsRbA/JFvDKijnvqR1fx9tlZdYodbcF3cZDq1IrHltk6VaDVA4nePXfmizA6rZjoMurQe70jr
TP/Eun+bJq9YxhuicEIuU6EC5eqFVIsjX4jlB0+H0r00QP2Cc2jAevAICS/FSVZBuy3MOq4p1HcC
E3MaG3cBT5vLnhRZ1T1WN/hTUzdbxs6VfCLQSG3f9ZuitZcTlrA5swdMrYpmWBJ0EfWYznfG8Y6s
BF3P59bvteCi2veXkbdATxUB5uPBOOili/rOFrowfNHqxpZDJiFMC8xDEoN032JI1j7FSna3EZzE
DY9Gw2J6VRC/anUQO9SEYE2BHOEM1IxENFGVLy8mfmyyheqjXG+4Q3JJWFFpD0N7gtJOzfrYk4IS
Ik3u1VJeUVVKIEmoM2+y4Dy1vz5e9C2dX2Sks28/T0OsWhnVXAGoWsRwmbpT9mt1KfaKJOi1sFI5
11/iTzceo3OIEQrkPxDvx184V59SMjdL57CfbWqGQiW7/QJAjD33+7Mn6il31fgyInj414K68Aim
Efp3sUGWaNehQxyRpk7xPfFKy6C9H5vNBKG83Y+W1HV1yEum+jhBQ9VYhvjN981zuUqMEon7X5lD
HwYRlItIglbhmxEMhJagDtqh8hkIMr3GEbTVK2tYx0nwULkIRqaQRAjywWxr0uwYOe+0+Jsaizmg
1GI6dNf38S3CGl4myeq3/AachOxNy9VSeDDx/eEL5g45Uq7hQylO/WTmmSq6yzdw3K5CajTwI0Ua
gSrK7sK1RSexnWBsGjogix2t7tnVbr3G5Nth7hD+NWSCOVCwElRdlfOQh5zQGlmkMrx/r8sYYcqb
PxS+TRd6NSCpq7mUD9ZD1LNiGdfXkPFeWM2i4i2hp/g0vl5NFd2stv33XbbvCmh8NcoDk4T4Fg8H
+Veu0x/IYij+sxGzcDwIvE7tJGRHmP6MtYf5Hz2rbUnGoIOpu3QwevQG0tbUSYaDCdCEi0Mmq5Tp
CpyEz150/dYut82aZ/RKdDZjVHTbQrP6WM0yOBRrb3DSiFop9bzEnn0lb6cpkkRb62vILR6pcTJV
9RTQfly3oi1U4AN0OBBoGhyGuUZGINWUBQZRU3a0X8Ykx8QMIKdwmGeXKoz2K/txIrbVhPPQKLaD
9tK60b2RttdKkraBCqzUMxv+XeA3zRMmGWei55aCbUlGGkjEfKT/yT08hy/ubjGLk7B4PU3N5YEg
i0CPjMPgAD0dNnXC/TJqvtKef+48WVhLiMBBraAsLXckW7D6uxxUVJSxKhuscVmuoShZ2cNPUS8w
SmWJkoHJ4oCkz4bdJxg2MWAEQuq1VtxpyHQtQYg02oanYXTBxXGZITJ/6WntQYyRpE91QpHRTX3s
j1f9Kc2SMV8ecE0Q6m27QBhCh5kyCXYWx//d2omChkAiQQ8lF/PqUFN2L+g09LgKv1TujgftnOw7
TCLZsFlTMCcwunm2hxVtyhZtTGgYhSvUJMsE09qtz9SMUHggDum6bc075XsbVZi9URTK9cTWIN4N
q9AIR9pqCVAO3jR6M11+pIYCv1yFqdc75rPSffK2yfvDIVriHPu1/zVMREEXkIYJqAR/uud1GOdy
hewExdFsDHaXs9w5PNO6bS4gQojAQTAJ7vnJsVVv1huUdurfPOXENTz5idFLt9yzAoueC8WC8dZu
2h3OsyyEo0+g3PP8BkdfitbfEpDVTy0I9SuYGMuA2GlRXX8Pbsy6IDCT9FHrFVXrYRENI5c/RRw0
zf7qLd/8APKG+x+WMdyHSERJO/fiamnyhkyNBswND+jgZFlWlBbKnAr1mXIuySUnCjIYUvEmAVE9
kgaKyn8/GXfi/nyaI/bOhfuuk+ILCwUrdZGTzzXo4tU/RpMjACpRPr6NqQZbshTntGgBt62aRDKT
XZ0KnrA+l6faVn0Kl5YYmLazaEf5Ym4/6uUbFIlAqVIucaLooffM0K2vEmZSiJwNUIqgYgFgJ4DG
cjhwM4qMw3LWiKK2z4I8UJXnvYqKjyzQF2qJXPZ1fbklMOJ9alBerCQINqJLGTKMHmjutrM/BoBn
X6Gnubt71ocS4/AZLP5HfKV89K4RXTz+tutEYf/KLkxq6988dvRMnPQ7B6nx7meiF+p4n7U6l7IC
9sou9Ip9QBwXeA9mI1N5B8F0bj3C3sq70ozPf/WyQFFkbH9CHxKNOixvNCyxMwfO2RDlsdSO3m0l
FXzze7XkUgds9DwF1rqtgrWg96Ex11hMtyfYyeOXDEs84AZpQSBQCvc7CzMLF7RZnk3LSwO0WW8Z
wpdQxIhY6S5q9YzUAHFO4vuwdlfjSYoqalFWr32FzFd1d+2o1n+8d4GNM1EO+N/UgjJjghyKTPwb
6xtdxdIaejMqp/dGHe6+NnhDopOuqk6JoYY+/p9Bp7zu/h7oKm8OcuLVKbKlEoQoJN9NJ7Xm0dbi
yx6S57HAhEYtEacuM2jIc2FGjRPM/q8BNHLsHDF1r5Z174jCk9i/4n7qGW1lJO1itebgvWKoh0il
foTPYK7dHeKeO2qsdkJ4jLy2XEO+sr4AiHS1Y5K+bVdHgJsPn4zurbX/AMpn/5WKVgWEy9P5ZEHe
ApNsF6MFQ3Ump8w38SrMk1qkoYBf5haXowpUMSJzGYyUN2KMhWoFjVci0xyyTQz2nUxKDFiKGqZ8
SFUknABjjRulIbQGr75p2cVmZER9p+KcPWq7VlZRVuU/THoZvjSmXvqmb/NJv1hFXHTwPBjQh/ud
TstJ+i3TvfV+T2QTcIKnrbbt2oB4/dB3EDXfYkyvs/M8N0hdglMTCqfIhkLIkYJPQ62BsrdUERt0
TZdMur5DBe7TXWGCmSYJywL8NrgJJEMQDfej5Eront71HZhchLjn3yonstPuiecV7l6MV6PsMxKI
AzPkZOEq7UJUGgz/JdXExKPr7eFTRGXsuUBeZEYVbWEZU0uiOy13B3qVbIagryU+VlidakVHUevC
xmSjIeANx99qtoMgj69x6XUUHLdW0+V56eT7MUG2nLViU7wot4lsfprUSZKMDEv5rFRLWOfbgjxK
RTsvvTvjaqKOOAiODpHOChFbFBOITagKzqS9vDfIQTl/Aexc/LPKm9j0ZMXZ/AMgrxLx5uYfytzA
QopheK2YOE90BQ0xuTgky0A+zIZ7EiVctEeO3eubx0d4W3AL1ZauKmw5k5iR5/+AvBCaWzzwgJuX
xR0J8jbKzTc0ibKPBwrtC5gz1VW1thn3W8rZ/KBMOBNEKr9QDgO0qz6jD5KmcDWqDp/oniI7P+QN
cA7F48J38pZf5b4bkXERr8sy65B78lZYzZ9Xcl1KoyrCAKkLjqtqqt5MjlXLgEBpCmYD1K/8Abvd
oSuGyPbgmJuK3tCTAtal5Fil1fiyASPJPGFVVqDWuRiLSsBSlpXBDO0hq8qmynqtnefvCVnf44g3
UDIpyAlMEraWYqLKd1o1mha0Ovxx1eyog0ae5DZXNPYkUjT+Z1MxD6qBXLF7LY9g6P8lr2dCLajf
GvR7gydy3O0lbHCMISnuMmrCE7WbnLb7QiNcb1bbJ3+8UNxXb+GJdJ6ve0ggG+2XdIvKbxfJjftQ
J8K8aOxAZ6OtfWYGK+NcncLlHqxGnGS4GQWrcomaah1POBhNg8T4FZn1TDrPBydA1OmVXZANe/9m
qyn4vjBLw0Erk6qyXw5XdPtreb52f9E3JLFNW766qtzzMC7/qnMWWHL/hN1UrF5uoMXJElJSUgRk
5a5OLCfEZnjfUfyVwJp2T4801nP1sX5sZtaRpgX/bjEcGE446nA0YH77dHc5JJhIkKCWxNJWcInV
rwubwpksKTb/U6gu8KIDvby0DaWY3p52gOSAPt5tdL05Fjl9sWOJ9QfR1YZRwM2kpmVTZBv21X/7
qVytJKx4gRShHsN1frvwZ49P4iOxMvSOgJJJsXbh41vBYe9y89FzIMLceEwvE+TotncfWAeFpZBp
7tRSScPBdw6SvjIrAhP72FVzci67HKmdj1w69pImcf8ipPdtMYMiF9c+mhdaUJuBVN0y3uLy3rB+
74Yd84v26KIxfspjcubRaP0wpCSP7shpDqeir5Cl3TgoQavd3Ej8JfjCf7kImK8AXpsr2tSzUW1i
+xhFRQwgFCR9is1cc681gWWU2YfGitp1CidG67utcyL+8i3MMLBdfK2mleTw/pHJ+pJyl1gIeE6e
dP8uBnhT1epjlC5KwJCeSsPaVnR09EPbKiexh8MZchoBp2hsr9y/WcSFIRZp4zf4OrA8Vjujzqcc
pjueiqWnHuhTPpKyn/kUt9CaSbPk4+02umW87qt1kKKzrehsJlxkVMWzWYBZEmLXvkTsvUvaSoVI
ekxNUQYlLSFhOv5KbMLPg5fC9d5K8E57ulLqbqnnEXwhCHtW2JwioDgPE0bK+ofXWCc/TNM5HQSO
TMZe1LXXyBWX0I8fhALavFoo3anvYdoigTCMYsazxyZFbbim/Oa3zcoD9ZISOoRxstIsSDe11BAp
WZLEMxRyormkKHChuX5hqeqFUmJ8kWxjYq+f4CYkn0AF0I3Vko12njDFlsXGvwAyCbWpCpGfkarU
UETZy/jvGz/LBcy7Zdl3bT2yuogOdRr+NjIaDWjQCHnsF6ETwX1ltv4joMuprvvz9YtvNEi5k2g2
+VNprxXudzRV9h4L4xLEOIpp0jpD2dRBMYy7hj/rkaeyZ4ShOVeLCoLTRT8Dbz/asNtf868Is/Ah
u6hI3AaLr2Rb/gRUhhFZ3R1VuPiU7JmaOfdOc59uN4V6WDfbP7ISySETKeANLKj3ku8Xuz360woJ
rP60OLTygmy/hsq2bYsaBaTDuc86HOcOEZUbb5XsfTm2KOVacmo1Mvlg2Igk50DALLnwNOopjoer
pDv6h5c5iQl3pLEmQDa4KvuTphQMQ1XmKlL/2pGtTOGbUsP7b7/3m9XGr8Mvdm05drr1TkVuff/v
DFVbbNw+W2c2CPrFUNIyYzMdFKkTTpjmFgN+t4/+qaAx/LQgVWqujDKSQYZLhBnzUyHPBa9QL7GC
wOS152QdP8Z8o9DEQ1SF0nCRTXJY3pE8VaAhsxLlSsOayZFW6b/De5cYFSTP0PsuD6xmMW3uDBvp
TLE0wFHjrSmNXHVv48U45A6uT1dkbHEkLOxX2e6PMKlYvPLAugzhvOw2DF8Lf9z33ODc1XYyG4wU
H9XKGB5PRG+XBpytTs7ssbZEpPusgNOzX14+8hdVe5HmUOXNrdfX4xLCmxSTfPyEvquKv1d1lMoi
Tn6Xpo6DJ5hWaghTNwM/4CQHBBDL1x4r2OoaqHv4rvyUoBI4P7Y/x3/868B9lDvOAJ8Cb1cYRY2l
AfGg6+ApKcL6mx/RGjqT8gsVMuI7bk932tVY6H0rBUIj6o8i1xEcfyHMtqIZgFoIWOL36BrWuhfQ
Lkwm8EDd95dNpeL9TOmDm1ngFh+pgR8l3nkV7uVrzfNnREoejNZqYCmRDZqye6n9pBqTU7SvIQUq
Nx2nHKZwgDbRR9Ud4ZZBENUIQPMfTH8ViaF45aewtQ00n4Ml2xNeObB6pcExFiLTnhVc0LZ6U1UC
nA4G5QPdGVTq+9ktWLuiUMmFk6XlHEwE4rLNKyFTvRiDGik5KQEun22dN1h20t7FexrWHX3ARmDl
lxDMNDpTwukbpeGO5m5+vJ8cmMxq/mHWpOdUuR55WCXUiq/yjy99Bf/VF/8stYnfa1zNd9VaWn6c
KBJSWA/ErNihtAvFF99+yRNJhr9+FXARSHg+VRvZ1A8/wkHi/eWr4x0DnrUkpB3hrPqZKLxrsPeb
pxUXx1olG/PJsLnZ+TTZp37HhDrQN0z/FLhN5Dh2FsyzmRA3YkJQOcxT4nuhCTQ0CqEgjRz2h94d
tapc1bsCf/2sfqCTl4XFthOOkOeIcpeV113ITZgctjtG+qO0l888Ynse5aP4GQuz072amLHvqcxf
/GqBl6JCh0Ja90uehY4oNuD14XXXL8Ax5Jbx9rldDiHiZLafYh0PJBjbT5FnQfQJbQouKajkRuNg
nx/kDlJ7FheLdOPAAgI5AgkVyCNFZLEEwOZcLUQLjWUsaz4TiJLaPdk7wr0bIDjLxwLykrKN2Vwy
IrueoGbZwdLWU91SGDQ2jICw95zGIoClfdSFbASjIbNZD4OEJ0ItnodhZzGHSvIY+PNBK3Y7ESrI
2b5SufjmVqEKtlKIMv87qqt+sgxRUmRftEqAyZTlYtBOsnixQfNUtGGvIqGgbBMd38jpA3CrdxKQ
C1X5UfArmTorbH02MLsYwQuoqw/rzNwpd7bZ/QE1wfEuOgTfydiPm8sqRtL0blLS3yLWieb9hCk5
V0Ni262ySyEFVap5tir/Jito+UMi0FxSa20GwPhgmewJb8aMfnaR9MqTdBLiU9rUB9GFOHFqrMtR
GIex2js3O785CZtOPMS/el9jcWKBJ352iYLwWpA8Q95cJz9uNSd5bc+IvqFSvLdXRfyBJRuFdoi/
9CRdP/8DFPzc/9I81uPu1pRPftWblrL8zTtw58bWPLiYlZdyO/bV8XtfWPa7/s2oOkwkMU4MkQVx
6tyfEr0LM2jJvuw6a5/m/msvF2jwCkfrjM8ebHf+CfoIlGrxNSC3iqtmFWUsGiCi3eI6IKJz3ilN
TRPFQWYQaWV4C39Dp7cw/Ff0UarWIkGYXtKrraRmH6D+eubpe6sauOutTiKBLRHeIQFTeovX32yf
mhQmPJd5fwZFcXWcJ3v80Z1qYO9Gw+lNYu4O+UBJUnvWUvN5aD4DtaXfp1iGjAcXW1pwyqKTLAco
0ClFWYCvaFASZ2lF2xC2LBkjQ+eDg23zJiXmx64wbyHWDbW0B1ouYaBa3P+YlQDmc+3J3gvDA69m
Cgc6XnfAOW+3kVkH694gEgv4IIdwcjQ7fHaejfe6tRtwyFT0bKewVX0enj7mCSpUBSwKmULKbgeE
JkiMn0QU1iau36FoE/OsXox8vcqahzzChuLNgM61R3mTO2uloGgackjOEpeG3GJanLYBQ7kszYVg
0QzfGDRr90vcJHfyHx93kDocCRYaXRj+vGXH1/hgqXTCjzNHCpK2Gbi+PfZsP5EFyFJClVVpcI0/
nhNoOq8t8qogSolrlfday3qMGZx6yObxPI75TmNWVRO2zXADWK3+BxiGi6b2xE7DCS5irT17L7y+
TqLqg5xxgZrRR8+uZquUdIE2RpRXPoyL/BWM36IBBGs0H0hMm71sFGChOTjcee3ASs1uqYeQctJs
anoNLn3x0tw8gp5+IX/NP4mM/2v61LHLuabsYV8ofkxILjR2VnhEQEoZ+8F9BHtXQe9JlpiOn+Z4
TLrfAyLQgeAYSKBhEQSG2hc99nkFdexpuRgCw2MqxzMDmbOSMImy99V4cE1jGz4CiIk7iWEGh0lx
u8etHMqklYRt9z4Sh1miWDZsOOXk1/FQn1pCjwnEkzSATfsyHKyMN/YI0Nde0Sk/kvngU6HpdUFQ
GEROJ4gLvGOxXZXHEnBnxODYMiYA2MiTqJVw+ggGBcQw6bF+TZibiyxJHu4ZPbt4QHckT7nu07bE
34rEvkKq/Fwgvc6EmElWen/gPkNbaC3ske0PKen378Mefwv4XTAZ+0euqjBB72eSbI+Ma6jV+uh8
CZ3VtvDDQK+bc2jWCp4lTJpU9UpNpqTrTAT+6lKGWwcCMtyop/bWEKmDgYTg3XzDQIq6lhq5/Gl3
2owbxyjH1XydDxjYbYk3AW/2uhKbHYOIeOMycVeOOF1IjZ8Ub8110pbrwvbcbVtKPhixQTtk9Z7U
eO+BO/Be8M6eaxOTWDJd99uMy7umEeIxDEXBbAjJkMclhpsY1xaCrtBpmnhvaawguqhJpq01ayT2
ay9RSY5kvEvc7LFfCN+lvZfqWDTLQl0vA2C/7o6FLhWXvM2NdeF8f30ETJV/mBigpd6UdsH3xtK+
EwJbhAeMq/k93KH7Jz+sapTSaHs8ppAM0w/iepmLkAsvN7+pkHo8n8n1dfcUOXJeF49ZFKLSuXoS
PgCfN3jRGjwllIp/+oYUo135yj6aKZtOzXNisGu2hwj9tbli1pvxa+VIaOLIhEAkYqcU1y0Tgypg
6TlruhwQ4N+D8s+os8CnPVqkhkgsARjmXOFRUQKkXWzNKlLtusLc/HKiJCZpjwkKehgWe2B9Obdr
voZ0/z+G0ioKfiXC7GP5rViNk2wU6luv1kbTBxgqwYfO3BQ+bnsIYDNVMmOwhtI4fNOylxUI8cuD
53UEgm4GPjpVefOkUEOCjJ1ZLf1xBLCPXRgkHfPY08ipkxfXtA3B5ouQlz+GdyHAZPtSXRoGHDWT
U1mgGxkFHQK1GG+G79UA86Yd8xmdn3bKkGm5iyUKOIlZ6Ydvkx5xsnBXo+cpBc9hicDvRKJviWGg
C2opelx59B9nIOPnid4vKiIO1Tu8oS3R5FXH21yul1Urp1vMzfoxaD8AKQEtA3UKe+tN9ZQVBAgy
XAY8/+sGkNWLEyvZXymNgEVjCZqZATH9mupXx+4mtOUG/+Am+H9fwcQZ3H09i6Inmw2hc3RIjvq1
Wjpy+ClyYyEPNS4m6fVkucOGWAuxbgK+wANiYvExnT3qDIKxzOzSNRqT+2DylEPbdalkfmJKnEtC
iCkxJVdcPUag1l9rs9PwxI48tkdQ1z74JZ9SOxJsRK/p5kQziwOWUohKqPkj4b8x0aNodl34Bb29
qBTx/v5NA4XHBGEESG080g3354kzzvCLnEZEai3x1Le6DAb2uNe9iDToSI5MzFxSU3YQph4l27Sd
um75+qxLpJszJAbEUFRy9mX3uWIwDoKmz1jgLbz9M1oSxaN3V0dp59F+mdr8wlGRaAugHndotrEo
5O1NgPVVJ3/ESzBNG647jJlUz9JSnQC+S3YNXvsNueQiL9RbUu9FogOiIJHfAxOLH/Sqkak9o1G4
RIiVmELJe4zAMa6t+vas1KAlUayUV6786V3s2s1leenDBe+LW+Wp8iV8rtz3W5o8Z1MTFKF+4C1h
0mjI63tlIMPS5CLsDCIp9/g5srLj8VyqHViOFrh5r7Xooay/MFRaaqmeN/Fo1U+38wFnFtBfutkL
t7LtJXJs2fojGbA8XKkgGf2UIIlRvRjAJZuaqnuRyBWNaoPGl7DEOYJ/JR8x+3/QyJjeC60a3msl
KK1cZp5yBjPYetURyORp31xTkd+0nY4Laq5O2tvQ0Fd60vWgMMRWUuCVtTpVz5qO1tuoUJDcxhdT
9e4ZeWQQGB4tdX4Lc95cZ/NdHJ4kqhNfXhnmG/AcDCWrGWrE+cVkkugIwyQAoLfeFxToA2j46sPb
23JoV4QLoiRT+seRCcUWnBqm/14L6hSO6hSSf+T1GTo8EyieKM2ILdgj1tngM7bn6IRtH1q+yp4G
7B3icKlFSCCU7gYpayZd8uR57JV5vq4IkJe4QIxwwPrGhfluSEiHU/GnzrwY5d9ebJBGsbbxxCQX
M7SaoWR5wU9YrgF46RzPijLWABlYTgR8GCBR5k+g1FwQXiJTJGL8T8Qa3hQn4pfB6rzDPL3kjJ7D
JaYKMqOtITt2F57FcjolVR2ScqZQ0Dy/O60dCBscKh/4qp41VjiCocyll1sqmsw/x2UcYl9S/c+2
YjowaGseFnUf/te5lx1yKlbcUy2DCRgKix2cBQhtEAQYdvhlAffzSo19N8CekrPfQMG5OMX92crd
H2bKTwNjhIvel0B67KZsdnkqQ+grg+GAJ5ZxUUfzbcIfi1xxt34hA8gcGICDpPHLPz53TqVcQyt3
vQa6x4Vh57QdHpIDVn8pHHGHowPjxEiKix6k3oXjoN5HeXYOLyg/VZfTSbHXbimViBLKoxCWihD1
h6iQW/WDTb9G1i4+UeEs0Bnnnb+baFkiWNz0wINlVjq/eSU4eINwy386OseiOZm9ek0bM3Y3CiiE
4mpKRTxgs43Ed39ExIui4WkNzV5Jjr1kkVDAvTsuafIkf9S3zl1gIwpKkCfeYUcCmszaKr7Y6enJ
jwVyR3chAwTKjsH+MZ54/oMDjUxSItwrQMm/56KeI+7R20JMxmh1X5zybHmh5QNuoj9F3/yKF3Zx
sJP02P171OGxu27lHGq/8/9woeBssMofbOtDaYcOaAPaIdqgsx7zKt1NAxzWDqpV3UNxegD2dR7f
mDHZvKa70li0wBpXEo9vtzgV6L4IvMTwtfp0e85UdzUbmFmPOEf0d6SN9kDfNax4WIxnRBGS/oBH
mwVCdeIF0CDsPvt/CeyBh9/8yKZJnb2trQlQZWlSGc6KbPzLdl+k8v2CnVjXfy0e/ivznoU8n8Kd
8KUDgP2oQAW7YefVPihmm9ONXXAc25Lv9JTV5L6TOkTksqDW/5tUf1AxxCNl7hv42UUp+yhuEgZU
l3suC2oowgkhmyDzRQLBS4yFfVuvAi9pt0I+OaU+jqVeAyHlsI6Ax4cI193bO9f+8MZAfg6ziQ0Y
Q01PWpjN0ld1siaqgA9PrPz7flGDuMWSAzqXA3u0vXvTmvkifq+qyeVXiBE3ZPzPe9bm84Z9v/5o
250SqB24QrJmT+benRI4rcQLBEjY3JLU46YwfRPqfRBk4WA05+uykBcJZ0Ql+neBq8koXzJJoZwW
QXKa9TciSPX/C5ooWq8cbd5zXdyS7Phkyn0YqQilfPuN4xc9LBzvgAF9KARZb+Lp9wgAxmDrzJJh
tCq47i8RN9OOdvv0wamn/+hWsTOTVAZyMTydirWKK+mR5iU6zmDG7MwJsaWg6FhcXd5aPNi49VSX
bO4sQmnjQu7Vk97Pt7AVVrEZ9e7dYrS0T1QN5TAT4DVzjuI0XHjVDlKAKfWVEgHvb4rUCG44X87+
v4t1ebAiL4irxk5MDwoPwACEvzxA8WCve4WSiYj0+XNzYqDbPH2+EYx0yVIIg0K6qwsILdunynLk
RIOg22xOnQrNbYliO9xe8q62z5BTtYGkgyDdxWwSMRjCACSrwMlXv2Ie72YvBsjbZRc3LVdYScch
Of1L4xy0UuBavBNmI9sIvywtXfi/PFmzbg+SVuCRxVb/LuyObfvtdTY1rG8C2TYo3X2QQ5TpzEHR
1nRTU8a1OR6akVSe5uxRUEg/MxCiKt9hREHFm5L/uKSlqfrdEvEvM+y18F+ri+RDqZVJf2kfZcAy
svWLXiFv2jP54gNhlDr7h5wG+ZaneejCTcd4zdAWxGINGqrN3UoWuoKhOcUIqA1zPb9ALy7gpQ73
N9RQOD38Cqtzpwik/dy5pHjbpvEduYzlLwYHqheGjJllG3ttthugNiiiikBIGPNXasD7RfiKA+Gp
wqTbUul4UPBN0/YuoMVjttEB1l04VRP1H2RihfUzDDDVAVs/Y8fTJK5HZARO5P9KhAVkEZfttGi8
Q2G+46ZWtnSpU7Fz+swYz3EDiMwv4bvuwyXq9nAdqZJ763wPH8foJ7alKbGA4i+ZkU3kiX1PqmD/
MWspMeXj0E2Ntt8tPuj9dZ3tCG7vNq12Ao0SwXfaRTXOeGTOSHiMaG12WaiTxyRdnpZp3Sf3JRNR
iyFgsT0ZKf/xkDGbZtKPIVzmNRQd7CFquvoBckAzSp4f0axaiJDhAOQx2u6ibCt7xD6OuGDyjMcQ
ivKJBlbbvuFVP55XsIOMKhK6qbqwSfLL3Qk/58zOAVVqB8g1HlCeJjbkra3RQd1j4zqtw1Ufl7yh
uaW+69/H7RxHPhCv1TCXSl62nY/IB375HSRKDZsgmOVGaJ3yuXZnC/esehKS6m33aOop1hi8MRP4
9UYqb624/pnd/T2j684O6Qn71Qk3uW0Nz/lZCKe0v6Vb5mveNmykh9Hj32GRnoZjcKNzt+FdK6uV
i4ODRVBcKmrogiVE5iX/J5Nr/UPA8UXB9h4j0OVwvOhOuTr7IJ8abcMNqq9OznvEI+TdHIAVyg6Z
pZ+hjJD8ejf9UJoPYeyl62FF9N0jyn4bFuE8/7BOrMVID7bgS6YwAd0od4ok7T06ITZ496zM1Tno
lA47LFi9n4iIR3jHGrqXuKISZ7WcfItmlACZI+LtF02VisIYtq71DxAHgd7wAQt2eZe/3h7x3Eir
O8L3vtP5afn41zsgRwy49ve+26l1/62SUHkFl1ijPBs+rZo3PJuGwSd+BHgv1w5cA0omheBShRkF
P+wnOYlqL0t8xisKy7643y3tB2u24tjo9XrsuotY7hqr6cRC89r1dE9VaLI34cnSDBB8v/LAjvpb
R1dieqApSP55vi6DTuTiFSka3Jr08xlJvGVlz5Y63magh5k4f4cbll/sZN2puzee/sc+Dv99AAJN
nrtYOm9dRoQNBfZHsvafs9of6iehNGvlhRrDLatWQ5Clv+/i8Uc2NfPWG+JSi+nW2rYTQbaagDHZ
JIsGwffMsBFq4TvBTWlyR5FIUtR+pRm1vlXt4ZW15oTHYSZkjqe1Kn2XLDVq5AkZUNsjw7NUdfIs
WOWTc3RkvzzkJhIJ/Lp+YyVhe74af66D3J6yv9AmNvZNNzLl5EAbwdD/E3oVKB4H5J0yIFsK0/xw
mnbPjIyAz1lTLxYQOBWoxNbLFcQSJwNLTZBKwdAJQjRcWkAMp6n7tPmfLMGRRFlAp/9kWXPv+qJQ
n7gG6nN1q6EoVD7CFJW3zdIC5D/y078YmzXcSpSVncjfxm5hmg/rENhJPrjSGrz8tcL+fHvBi9Ml
ymOndqM2p9271OZRK0uX50aMlIZcYh3CQY67W6UuWK3C2y0mZ8XFsVn0LfTWgsVmuY3HFvkjPJcw
tCvQLjnSSJRmeXEsS957pOeDrp2perK7j8UsjI5LdKK7vPHIJHRQNRlmz5Rjrx/1KFHHJsmp2WvX
ClDJtRpywQV36o3iLj0yVLX7WF64YxL4o553YnQJrK9hbKn39Hkf8b9QUfdGUpG1BJWso3ttYJd/
zMyoAV7AsRWpi4UF+BgfTM0ECjdJaFpC1ctt3SkI657i7hoGly8ft8X01IdoDcTDtnCdJeKl6L+v
TM1/8YylDL33PJIILUSsMCdQM4W8LE4lgYPlyCnAcmKGTUD8iddS+GlBuI5OPt+Xw+kDp9mzJoSp
M1OFYAObtv3jxXY/VtnB7hqBJ9clYRE8CqaworK4iuydS0JW7PSK/Vgyf6bOBEHlCtRn6QpDmzhv
MEqHBwTYF8qK04xD18wsPy/JwfaZZLJtYjgnnzQNs4Ek/a787Qx3qVoN+iZ7mKJwiW5hE+IWKe6N
OufYG4nLE95wM57Tu8hkr/3E1ODTPixdq3lpyN1mQ1lTpzE8gVvEW4Gzk0K0nMh1Ni/7u09tIm7U
qQ4B/GPHmO8cMGFVlifuKPPJbzTJ4N5wEYszDKS/8NyD8dVKIufUMWiMkHVcbqmxr3bSN3b2Tceq
4IEygKpPESqEF3vxmCfJY9ml4Uju0+xPwtc7bo3XOIINlhMJs5nPJpL+NihyU1hVhyDgZpiPNwuB
fnQVJHrSPZNu5OoPtwXO655U8s9zBrmY1VnJEDcytsmZkFiUPFPZg8zgwSDmC7PlDK5/C+0UAOil
LtXPXm42MptjDP+0gRerY7dL2hbiug8Bi6d0uQlHoac9x9W07XbQcZ4e3twCo8i1UoNVI0A0keir
GrGMdxMUitpDknWAWI+s6kJj7PNNff8txLok4gOhw7KGdstp+LCEERIVC1Lg1VBFbKEYx8HCtAlg
3BlLP3gEJgS10QNuNrHGMnFhU1uhs44sRCZ3G9Cm2MGu/XHTpk/GIbbkbUb8un+by7Hz3eOkpY/G
lc8U4Rc4CFw2mvIvObaEL4gko2I1byLxKq/j0pwz8HErJHnLinZLEVLJ1f8c+7hxJ8Rc5Ng5/JP8
dguLnPdMuehtZMiZJKVP/QTnbTvBiMVsKrsuGfhe+fGUkK4WCYPdSft1sfnmPQiqXiRG6WcBMyh/
JhEeUdhY0X9nukbC349zX3hiWHE/7IOO2LGs4afsIQYlSlWz8QaHMMgdEPRllhH3faS6e9judfB8
GlOulELUHqgrZpEH5NZw7+a+sZTq0bTb1uC4qpRfF18DKfEHrbhHl+XG4Ngyn4GOveFrVlCb2exO
po0uvUITryqYNOGi2awWgVVqqB/f5200jXRh8MziqKaiTJMOdCicG92cRKKhMFh6lRrRfkFIIVnR
WR7LiKrhrdg4aRtYrO8J2By1UXwXLezwAlJyLmRTnmqA/wbbKlPnibFLWSK8Hz2kaNUEbnUSd7NN
LKxr5psv7/uFnDs+Fwgb7N6TKKWU4NOR5tOn6Qv4z6gRGPL3Ipn/qyJZeN2rMdMP2X2hakjoM+BY
K5VM82hZMTBDJfv6VVQzYiqTfrOt0Fpwqjzq4EWgdeY+0o7dpls5NBn0QEP14xFnIM+dCGEJEG0K
oqMVUEAxO+odQd3DxLZOEMGb22ck8fYqKfoEVoJPwkE8W5C/j/S7M7SBRdHfMxC4f3BB6KlKTPuj
fuxLISau2+yiSOH8ioBqNTDT8zMkB5E6Madyl0JVrYTl1cGM81DUjAk4wsyhE6iDHPKb3mOoIqWZ
SoQEzv37nxlvPaZ8H4UZx9ULay8HpD0fc6bMfxJloIlcJjGebYY4eQSngEkVkojfmHITfM3xxdMn
ZlJPB5EubK8dndUNXHvs+/H6l+HWZ7GnkbTTNaMMRMXOxgRtBkXA9jt28fDgewVrkOwJgg1ceIBW
azKy2JbyL8FuVMyWQMUEL9H0WHptuc0yWHp4t2cEOE/Nnvg/joNSijcyunmT6YpBCpoJBISTxlGS
jReoLHxAFyJnOryU5nhbJ1V66ugGsXFCRyg7xqnC4VvkTkSdJSi/+Ep7ULvjQh0tsEs4PQtFIJYu
hNgTgvb+4vmuClKsbsQf+vfzsNpCkCqsqNvuAREuZym479MCpHEDbKUNluW6yKNGsnbhXtQhW2N9
D8Cn5zAP7KK47gkopm4lebxh7N79Rm0jkhTs7PODN7VlG6JinPHpXC8T4CWBF+6fEcZiCVF/2z59
+j870tSN2NUlJxW2LxsDivuJDXH8WlBM3Xv3vNCArybb/eCK0clmDiQ/HkhjaVSGfflW3POgdqkK
hgXYXwSVdbv98zX1VVxBHXdnSQjEI+MQBhU3AlGlRPTTZLLqllyqs0LhQMPMznvVtTv0Vgh93V+t
3/YjEP8Wy8ZJaRFOGAgiCRUDcUD5u+TbjBJCJipWX7c+7xfvCqQOvyfFQga4puHptpFDKkdYGFO4
tu91Mi0kGa+uxSgF3vvR9rZLE2IgvBTXsJRC5p1CVA22TwYrQ/L1qz6BZmJEsdYIWDs0qDid5jRK
3Fw/x+l0fYNxjledPcxWhJPdwMjfgv/7mhbxfE/kLPGe9WcNt+PXuYSpefx6P3TWdNUYalja7hGa
N36myAuWRzbSORiBYFW490Gt4KpXDC3mtrQUZKIPuOpfMFDc2DXRteyJr1noPjplvDQVqdDGg/9M
83Lh29q7Ugf+kflGy17nRyO7x2/ajd6oWmbbM0PJ2T6ab6OqpaWMKK9CLSqo0F7fcDCbvjp6Z70b
tEhfMgSvJmMcG9zefCtKyJBpDHGu3K7XnAZjDGCvdC3eQIHMPMgPtCzc9R0Vz34W0UMPAQBS/5jl
rucX+vaJLmwjg4a5EEs/RHrBvHjyiMMsZYHf8waXijlJBkTiToAVWcAFVn4vI6mpdF0zdIH8sjK5
WJl8xJ1cV8yKLkQibZ4E9VwnlYyAKk5od6759XfcuiQINkc8Qhvd6bUoABBWIeB8UD1FjhHg9yNZ
RVypQsriksBuCJnGqzD0VrjNzYjrU6w8ftliu7l+WfT7euHqhnlvXccJJvDHG9NMVFtVT0z5Lzc7
wRvpvNkZ+XU1pqgLiY2R/Z45MdeKGW5V4XJwRNT0Q1N0fkhhsD6OQr2Ku027AoVy8/ScX0D8jarz
aCH1d2s6ZZN4qLPEpe9sE0L1LxKpDhUxOp6rIc+ceadgc2WRLl2hA/2oLa/KPDgkHdpI9WxjsY23
Wekm+XKopPOwi/vd+RbZSKVHsQRJkuapQvMz5HKHFOBcTnvWwfgnrCCPo+I0Fu/Xg7n3ZeZBIQPy
hnmoh+oCl6nNNTsWM1lnIidVyQ/JbuRHSISpeh29Yxtcsoj+Y0R48bNAraAYqwa6oDTwlsOpsyDo
jVeYk8aZWOiq2LLYlwetBsSreXvW4pIsVDbrFbMN2U2n02dOezt9zxtQwvWfkKfbODzjPQyRydeu
I7CHUS9bV2cZr5BmXpgtMDJot4of7ttJeshghiR59AIwCAtl/jtO7O8/H6rw0zkbteY5JnFDjZlW
d2dsQZSPX5JLAiU49zevhowZ/uemRASdIZ7eSwVgILQ8GGJX8YJYzCf9GiVT0ntlbVgjrR7zoQ8P
7edSMBQS5cTgXaQrmapfqrwICTBCsLE6D9PMczQWYolCogufju3cVAyl15gl0EUw9Ia3/VePvZRV
UidAffUXvzPIxKfgk1sikW3pOoAren642eBcRMOZzO4YGwetE4s7Pb4VsrMX+dvZ9xWn8w/JxMW3
CpSBTb8ISs1dUHOcTZCny3ptOUAkCwKgciq8pV0f0DetncOaloWM17PpyXOiTZn3wgpZEx0fm7Hn
WtRkx5DI0kFqzNdlz/oT2H0ssfTjCzu1A5CxH6QBEmHfR/Fi30xpF1GX0xRQL7w/v3JF2DLe3aty
BlydyTUWu6F98vJXMzUeC6cuFq8BUQXuVex5Ue5b2gasMiOMhPFr69Uofm1ZJtsqxUPown+CbtE5
pPOfNwy10mtw8/COKBtxUVWmn73ZJjjRbA3YIFVwxGhwW2jd33giCR77xNksG4oYanSV3ijX0DPJ
9MIF0jXqwHIIwpnbQtsW0PwOY3SnXiShAJouhifwZkrkjiEhI21LfsqSNw4UwHE96AXGFnBWl2s6
GE3bENyWwVXrwh3dGdUYf9Gdk3/atd5+vfmVeOQuXNYyTQ7ze407/K1B63UR3rHsxz1edQ2fi//B
G5SjrfURqHVV1on14YKJt1rvOA3o/ZVRx9uu9KEY5WM8O0haRYCLvqG1MPOwKixttphTMRKT7YGP
75HnYHt/umbolmkJjqYJ5aWqBOv1J4HuoL5QOckSLLsGm/ON6y2IYBF8oZ7mxD5FgjEoNZL9Sfgo
V9xRC+DGrtrAHvGLP+oFNfD2+T5zkMcIAyQzcNiDZOyxYJBRTnEViH2mQHfyfPxy+sZhuxwUcl2X
DYXxGfEO9bzI3cS2ppCXq1RpAIeJ8Px7VuAqIKEyFgPiGRSUZDVykCMAKKDx4VSGQK+8GWhcGiJq
DKIEXhqLTI/3uzhIj0aKVMn/ld821hDZ6QvlENZVxVUV2DnNoQCE3EZiVKQYsqLiMeDPCCXy2kan
TcpeOomoAxi/7BHJzp3PIPnqKFEAj5bzVvNoof73tgEXnmOofnPKrxRynOa7QZWVk2BJYI7B2C+r
2phWJiQj+dSAVYbZxqfIcIj0Nic/syrb8rEzehmW7NfMSyy1ZaeBR3oOz/w4LLE2xTCevOvj9h8U
guWAi2drk+rD++0CniI3cI4P7J0d/2jBD5O+IrRpPYaUmWeXKMpVQI2jRlnZW+KXiBlG5Xq5qXby
yyyPYuFAy127W1GuQ4a8iBFcKQjIh+qrMgl736jLTKuVH/jvCBAnYKaXADYIdG9tq1cYtvnT2vj8
YdH5TdQGia1ERtmWyQchcTu1rE4q0Hc9ulhR83gqx8otWhpQkoSV0uOODj/TeRVXWjLt0a7jtuBo
e9wRTcBaC2O+v2prU/TlivgJpR7BPFv3JKSq2uYC9dZE9bnBmNev5cW+ityM+3ka6argHR10i8Bl
//k32PfXZW4dIRCq0IOl5ZzOZJn5OCeKLml5UNntyaFGUEEgtiOwuqKbjIAjC/ncwingXF2T376N
e4atDNrJSqSIQ+G5L7VRDaNaH2IjQ1ahQoa90u3cCaKMf6tdQJDkWtzNT3R2xfWFHi1Rn6E/7KM/
LVC/n8qPReNoqbaG25Qphk92jqTDkZ8GefkVbM5Noch3if8kmtTQPyP9WrdC/w2g6UGEtQMElsr8
4UXEa2QjDkjA3T05rvJ3b6DgobBMrvOiPYmMRIewcR5YvN3ZUJhm3wKU9AjIvssOHhZIKy2uXYqF
L0860gxBLT5Gs18OLvrdw82pMpt98Eh5F3XT+u8xShZlqV64UPGU+/Nb5z7/5WuXfcHIuvgbmm5+
EyLkWD+TnLEC3kM81YABo/tfUjoZS5AZBO+K80BVXo+R9yJ3TYE9OjgwytnhZiFXUd4xDRVGknIL
FMoO4R2aidPa7HSLrKbs8peQIp2XmLpk4+UJTWU93E19Lsr0TD8Wo0Hc6rf0vF8GVCBFlzMPRhfv
m+6K/DuDtzOzRpIpkOxtkz/CGbJJxaDxVXqSFnLkLx/Rf/ct/geggQxkLO83fBrynm3BFl6E5/13
3cIWt8bZd5noHoe6gVBAZTjVveGa0unxp7sF3kPf8JBB5cNIP8nFbBn6HFGyRHrLuoYrNI4aZIxj
49CQNu/HLfgkzYRlMwsXIR6EiKrf8OexrAiJb+sXgUPzjQzedkGBsOZrV7fq0O+tM+QIApzxSeBz
qlSu4WNXq9DTAD4UN9aHSqoUXwMnPQeK4RV7+3USbyL0Hi668NceqQqDj+9aYHnjbOeoQa4IJWDh
8P9WS1iz0QzcyiTzzE+0yTUC9/e9uqN119L/c0q/+yrCuGsaAAnj/n3II3EZ+YdCi9zzTdw2b/B+
IUD7oOeyvRA0KIzEnag1zL5NVe7xaVwrw6LJ8nG8PoBpoo4uBW+1LQpGIK7wXSwELugxwMqgb1Vq
gK+tzQAlfYsRI85U1sDcHAnJIOYC0nSB1HH3zWpE3uRhNU7uW/kqNXfXmk43plCDqIegIDsqV47H
+lM9/marUMOx7Zc+GM/Y1mwbVjtjiKMZvBuy1j8kzp980brVcRB3Z3gDocBwiHJlnoAaOavND1zb
XgeYmjn750b5mV7/aSY4z2wZyW/nFHqoAIOLYWAjCezZjCpkdomIz9DdXGtcMWD8/y0HvUf2SqaM
hMk9cf4mB0tupo+laqfzjlITW7LuXtyMz/h13DOuT4eRpA5hpMbvzUA/riCEsNM2kT6DDVdhYefd
P64uJtRaVZYgnngFexPELwe7yC+vOWhTBaO3xN4itHWFKbrCe0DxqEd6RVKUJc9aC8hCXqNo3EgK
UGDPBkgRKsnMkVp7+ysFEbaDjSgeRYl6c9QX2Cq49c79OtE64wBDwkED7/59zsFIxraPrBa6kXN/
WtIaQzYNK8IFXWdZq52qXzAKkEAAyrMSc+TPQTWM6ou9Cn7sOStDtgWH1hPwDaAWEzNEYmj8FlZ4
zkvGQqWwLHE0/C9H6SnqQhoqm8QVjEoK5VhSDWb/VZPymSB7UDY9CLwTbQnt0yQW3oM0BQvzBPMY
sLhtn+duqR+HHvKXZDfbL0+KQEr/emWwhZOVVqGOoKYsmBWetKsDAhhuRhDopFL2TsLiaOINW+0V
ArvR+DaFcxrBpjVM4jrFtt+iJxaeoM2sAH1/iO6fMZqnL2b+Vv2SLHj7lW5RszPqzlIN+e1wER25
1jx+tG6/H+pzkb48zLR+B1M0ZoZ+0rJuhGPdLJtoifFIJpMKRXCMwU8i0SRzhfhwoT7FBBgn9TPR
xyRI/YgXX+fFC3vAD522rsNoAKoHQwaxe53DHjoBWmMpp4kWaD1PJqg8x32BodVxZm+fThYTo8uQ
akccv9A5MbdlvwwUIw6OroJF27TUeKuFKBBNIbh2IgQWvwAhbg/LS+4C29vn57fpktyK9ghmBt0D
zdevGu0h7jhNFm/8g+cFrwOFIG/2PL5gKswahq/GC3IoVkyapLwDh+CgVJetFtj5ynrIVkrVWM/m
x8VdDZsR2PYTHVtDLq7jUkjQWlrtbwHl412mVDHT+Xh0wQmkhRyssb8WzVL9K5qD0oLJXwHjZ5zr
OcMUFec0iSNY3rWX4bnl/d8VO6EwIjU+fqKcWMkKrvty3Eh1OQ52JLkxNlCC0/vEnyOLllDapoBo
YSw13Ld9Wy9ArX9ItPoS8zcM5gItMF1Oo3L4axQs1YblyCIIILy+OrxSVVXGwIu0obFVmY5sujhH
H+1reZSrLEgc70NPLoWyCqZm0cJdWum8ydvQhcU6R6aivOSEvIV3lru16GcudkwhBsf4ZROIuZRM
72+kBQUAYASKKhxTG46BMGTjJoyR2dzln6MTYkRDhW3V6fKB5INzlqtFAjj94ei9DKbMRNLM9l4X
bjlwGglklFQ1PtJOMKJYczTNwyXnmiu15tCLcy4ylP+wnDO7mIB9y0TJ+CG9620ZvH5yBf/w3BGy
EfN1UgGahMpXIg388hJhbOhFMtrAs7eUbJGoKLd2sQ22A2Jb6B3SeAk5bg29NoyWwK+Q7fPdhG1G
0t8RRbAQTyCgCwUZFKtUmmUI+cifCSKPGhkYCdOPSdkDZJdFgy5zKmTiGvRHlqvsN3YjfyPHhb3m
CuoGNL9G1IxX2ziw2rLn8yXVKEY5GwOUxu0aa6SdAB8vyNDveS+RR22/9vuLjM3VqvMVFd2Zm0CU
2tAPG5fLCGJE6x45+GklyNDuU+xhPrBKcI1kvkPnEZZFmkUTQOhoivkpTstB3e1oviHvtjGZJ4Nr
h2kdhCENBadq5zHjT8gwDwg8rSI0iU0kwF0+UjfpWwCdxjyfRFJW/tiaOI2XFQFPVMCSs1hUNxNB
XlquMwrI1hR8uOGuium52zdM9ySxa4yGnSUqON5Jq1bwtb3FlO9Wb6Kdtbh9rUERmS1JdecAX5CK
e6tdMHi+MbuCvWL9xbtpPUtq26bbHq/3M4IcnKxXX2ejqqGWfBTetOvFdNwnm/iahDQppciUokdx
OHa2eIkxvUxM5E3iMqkC3wlLYht0/xv6DNb1Fn53xLZvX9vylGnxAyQPRtASeyK5eXajhqPemoEH
XthK1ETfwh/3uN7VNAeheBOag8Xg3L86UuHs5JEOPqqdLsKGFb4P3Xw/7hoguq5YU96x+Y1RRhYy
L2Ceg4hXoF2uarNoqKgkBtcC+GAMR+AK4aanJj/uSU9XiqlayaKEo18udGzquVPC3ZZZLor4ePpN
/Cywc5IHXxBkf8B2ZtxoTWGtq9fVbeFVtaOpY7Xz6uIfMM2TeOTf+0I9KP4rQrUw1hMCCRLFWdbQ
Qgpf+1o3TItRjRRvHoXDOFyAPRhZwWxx5R2xroaN8M0KGhKRj6UiDCoDRAlcG6T4mFj9qXnh8391
BBSX8nvlROQiuhCq/NJt/yJAkZKdTvjmcHTXWK/ZZl4T3ABMGii0INZt+QtVb1GzLZ6vpjoymjdi
YgUmZjvXHe4pubeph4aatYyvPPUJsqalqxXVp7z7nJdnZnOTnci8WUf7nWOBUF3etKD2njl4fjrR
R6DLik1Q16H4jV2m8Luc6aT0KLMBf6EUWV0i1+YGKjMtBheSc+t+qcO28mS3oAGBkon+K6vWWUmV
83vYcNn3Xce+68oQ3FUv/nMNauV6IT3sveV/6tpXZXXSOnxQF9AcdQaZmlo7Y6ADcE0lGpnDZBf2
6jDdK2iupIszsXtvTLFYXvz/o3sylZFxG+clXvJULD6lPh8U6RLuF4gJxMZEb//kCxtvj0U2o2Wn
fyptGt9WL+bBFCMZs72CdCW4TngrCJV/nGFExs0GS/kFOLhDQOEoyBVffhWcbLrSaQ8pb3PquTUm
Ze0YRi/uUlbpuauXHtHX/f3T4WfI3gW2sKWDF1HB8HnCb4P7WKoh+pkeKiNEXaXHaOwI1cbroCGU
IC4Rxzd9u9tnMTMtrtBd2bGRmVg0cP58exrQRU17Npo4DtODS7C73thE+Ia0GpNDlmf4nWQqXxb0
ouSnn1n9sDupJhlbOo4gci6Mfzd2yyEdPHB5sxEUTf3nMkPjxSK7Xge0nAhEMYry5F4G3TeQPVte
3SrJYYBcqPgSiQqBI0aiTqZtzrEoTMhVCRq0yY7m2MVLkthlljssGLgEZ0w8CiF1sDdPXnyhXmx8
PoHTFQZmz1Rwk/numrrTaz1MkSKB7ZX8n21ffzpygocSm4/+NVAZTGZsQeJWS4PQlB3vhXI2O/DW
VQ+IaZDrAKVp5v1znm42eXSUt7G6Qcwz83CuBKr5joHZcOXtPuO9hS9jEHKF6e0kq4Begf1hsywj
OKJReD924P5WJVpNx+EUUg1GFePib8v6z6bij3etrjrSfkZlCnVNRz73DAkkNTywGSgzHW4i127s
dekp8j73Ur+ADD+y+HZZ4K87Rbnq+ZCQ7vSGDW7QQvzMWXNNULgPL9anFjb4VPrC5kVaDD8y+EQH
je00nTVARPlI3ahkQD/ZyHx7aGCNgWv00Ghl3riXmcGfVHrCJqOjX26tp+O4ZUQTzQl6Qxz4V0qE
f+vprGB/Judb8Rzi7UInEEfhEC/v8JW1kXnOv+I79wFhZG5ZnUbijK3jps94meFxElVspH54kRYd
ZHTElBIgAylPV48skCBk3p/bAORb9KUsgz0ihBqBL2u3vvGNVvlcCB+fUaOXW9Y0kuiJPwfRJSlN
lk1X1Gv804CapkYK1R8l5tX+DtvAlSjNSmKQo2KOpioL6ryZdumJiVPmb8jAQq4q5qC2lWRDNR+p
7Gq+tb9izYwNJ4dzRl82BygsIgQ4Gk7SeLOue1K9b6t7AHM26zbvkZH6fzgqy7leczOGJDFHGmWe
XGDeqCteJ2zFUGahw0lG7keE3q+jCUM+uRWtUpKPMwb6iM6UkPRN9HkrvuUNVbyWyYxRLLtmCTJL
HftC4T6wTW6pT0G7jUS/ESDqCx4VoqZ7uUk7X1mXEftM0+yGJLlnkIxy0mLe96wy/2XCYwu3GDyG
DNS24SX3MtmvkWMwLnQzmYIs4OWXCHDaf9Tid77oHk+3j+7FrqjzBUBEqY7hwiBoFIMqW0TV82zn
a7A9qE0CI8qeLPgzLxNE+U17bOtW6PPUTZ4PCONNOeN2fF8BR4oRmWv4aRWl2IKoGFjs4Exu7+HB
X2N3/mV5yU9WF7fb6Lk8UKUGXhxuqp39sjKg2cjhdIA6cPoLTrf/1xDp1tAiea+YO2wfjBxbu4i6
LL8dQhNdY/Sostz4xOvFvBc07l1XoYBG95oShXMOBqQSo9q6l9YByN0cewhs7mj2GaSgX0d6SXJ/
y5nheZNUuEdGoXMCfFmb43RjcXej8xQlQgmCXDm6OFg4D3U5QkyncgNT6CT2Y0Fcc5Gur+WZoD3N
8poKMM9Sd8fDMjx/++jZYzrRgwzyQOLfhbUX60FJ8E2aiHs6D4d3SFFZ3IchuyFfyxXR/XAUnakN
5uz3qbIw/ctJVAuja6WuEe6YSNN4mDZhgF1HGgvBHojRYe5s7NRvqH0CwlcsKx1dPIs0JhwdrO4d
U9GLBFf5Ir0aNGC/uEtTH8vaMOijniu1FBmv1MFi7Z1O29B8VMqYe+iGQbsslv4XvVsfcK3d45bb
AHkNXmQTpJHeawZ3yXeHHcdXNN0Rp+6jwIy0RpDdauGyZIBRL4W0/dAcm+83SyxbSHzCmo/Skz0i
QvkXUwq7UeAbz6tIXzR176Nay5pz1IS3f+fsVrePxoyIYl4JmGX3HUDu485oWHmFkGiZ0Zhuro2v
VUI5uliCWqRejXYaB9O3b6nRGfjd7YmlYPnh468MTRksDAWYyopA/XPSQKqujLXbqGif7GMFC3RE
N6mGGGS4YJRtb+G83l14OOQYw2jF27pVdGrHhrc7sRe1faKxhy9HYB17gG2yAdbKxT+vn1X2epUc
eN3gvJAhqqIOlosDUX/G80Qi26R+xSvR8+W4mJCQ9BpruywLmqmnyPkXnx7uRrrJKoGHawN8ae6J
GqD4skd1p1RvdZuCz+GJLHqMp6rc1hoxUXNFNcV5qe4cLFd3j0UP2TwYSgo9uuHr/ZZisGS/oI3i
fm2fs/S/mKZd5IboI+oG28VQohD8bwunHxT4IEXI34eS5MqdJanwQpoyFMKIbLhdMtJlt4UqbY8P
697NejoQKSPbyUF7aQHlqNJaOMYMkO4+yIqqjd6xi/2/HqO2FPnl+GILD38xj4dN0HYSWjGwI1Qm
ZSwL9rvPeyOvkpmmoX027qc+u/zLTO7BjPC38iZV8MkxeJx6hr1nNStSa16Lm6qrIo9ns7P4phz+
91irC7prrQpdG+EY4lFYpbc4MDDcv7Ae+v1tKqWWgsmwCs+oJMZ/aw7TNa1KniYJMJv7vcP2m/Fj
0iVGwABm9Ye9HJTymSvU7yE5qKOBRpbycAwEZqk/c14ops1UlYROxCrQ4XiraS61ggdABICYMfGK
LLD3aBFVeNTdfyFB0tvy/aN/IO8C9GKUEZ0VhgVjj9iV/PCqUZUDfyUM2lIQKsjkF0jDblfIy8iU
JhtozPXfhHIKgJHRJ+HLD5J35GkE1CQ3yYy3hlnavw7RG77MuIl3j9VdisGV5gS0V9UoqDm720ux
xun+CyWK36jfhJ+M8ga/5BXFmfZJ/VPbTgo4Ks/jvGiTusjo7MK1689FO/TpulrKASmXck+5aath
goR+Ut2Enf8H7/V+khJYJ6626pbzxxD8Q007FpDhWXqvOYPBw4zwl/ZATnCMAHdVUAUogqKW3To1
MWx4PHKx3ENp6iYNZODzBsrx0GKt2t/ZpZalItWdT70zURHRnknD9Op38KPI2shNHK3ypOMYMj2e
HWJHrphhayA/Q8d/3pAhUrRzDPQyqj2Nmdi0HWZf1i5zNHkjHX9P98GLPNWB/lGoVk3PCqSnxRbG
17Pxvzj92Jg8Sh8MGSYZQ9xdFc1mIJ7REpMMjSyQX5DsEuzKGOoBih+j6Gd0JA9/b8Tzwjw4hpAG
vb1mzYQ84eGMlFVWxyxuPM/eZiLaNto2Ob9PBGMVDeej/p0aj3H+8GnVmGyBsf0fLqzT2OF7ncoL
TGcsJg5u5bFg/RtJiDkyXgp1f0BVqUJPkN4g+PdDmSOCng9wORDcisqq1fEhu5MYwYVCyqTXt+qg
Db9LDV9XZkX8+y2nDVFU2mriNZ5C2GJc41JA764jA5qF1Fqm2Jen6PKcS05PFUG6MjyymZsWKRKP
4VJ3+Kvv/yviQ7gh5QIX/YrIr8vk2Kh6lsE+hgHgPtZU6wzPUKGPofQQjqxVxH9afWcS0/I46k6J
QXvMoEFtOBvItagKyouxplVXyrS4cxNLntyuCg1Kpz/fQQHO9YXeDBakheq5mE1HGGXb/5Qb7pBC
nfYr7YGhidk8XcInXkAhSih8cHOc+TdzZx7F83iiXTfO+/348Q5+yG1oERQsCmfvLoyyB16eVRYC
f/th0L9L+Ycf+47eHcOAxl3eqPHnM3TJqjWrJkX+pCR2r+LBZsSorWpKZLOg0Bg53G7mpbPuYYU6
LuiFzSgLKfT83UiO1xcjThLoZGSnbSo0eO1YaA1e7kQKqK7/9zXBdoavzVSsxKhDgZj2EhX4yLD+
ika92TNyEnB3Rg+xM83bsHD2L0ClCQSGCVczI9lPgws4UNIkhKaYMub430EQ7k5Rli+4AgQW8p8J
nrm3K04J/l3qOck54L5a2HCV8QwK8MAe1k5gqs5fzUPV30h/ELPF0qW1FEABmMUzJLxqGmfGw/Vu
cM4OWtIFm2GHKfX5tzhb4kRSl3XifdyoJR6J+i00V/3bQG7aeANke5EUCidkRooz8kIHAI36XFEA
/3+r8rBRQORgthkbVFdrGJIGVmUjIjXYLXzk4Y3DsDRIbQcaQVmI8KJIMTwJwwId7kEeGW4bD+ot
wTiFYtwhpPtpaQaCXd9T6LWE/p/uUZq7QV2Lk1xtAko8YRTVJ2TjpeiGwaGR0CXj++gKtmfhefk8
ZqQa7ptJpgAxJes6rlZ1v9ndYadEmd6yuJhcu1JOCY5XE1GVG0lmMcjTkzHwjkt07UjNT3M4trM4
nslzQojOUMT90df+qWRqWFolaWaQLUc94JnshTHJ6P66X/LK/DHlLYI38BtNnCrkvaIS1h8t7/Xv
S/hczmFtn/oGo3kUQJY90GXm38VtYtRj02Auo3ygx4GqtYqSQeYDsl3D8RynF1Y5vey1eD2xRPq6
SaaQTJaV9uQApeXrk0pUSMeWMT5r2A931jdGIHijw9IUgQikSySblXf0q7rTy/g9k/FQ8+A+EZqE
TEMZqXmWwSAw2Vg4X/TjtcBSnbBgcYUHWkwr6pZbULSdMH41tU4yCjKx7OVl244UQwv0ptS2nThW
vlxQ9LmJ1UttOMKrBsvLNL56jyyylVVuLKRT4x5r+E46Aqn5SMG92UPldNNO7WJ665VmRg2IVntx
FOMOIGJlMVldK3ub2rQwV2SRm/gGOeJDiE8gjvjbTcsK5oBJUDl5g0QoYlAPp1f5r3KNXdkq+/Dp
5mF9H7kLVMfQj9EZEOCHg3LyjF2Bvh7iIOYWtY7S1Oqdt/WMoBSebvEcZ7Fqjsi9gCnZqEmXe9g1
DNrTSZWokiJHi/oF7atAeURis436sinLWb1/xiPfZwcXpUQ+cG9NYnilY/xgc3o+Ph1C9jyoxysw
lL4986xBqV3JToLbeLO5OD04zcgjPS8jcWCFrwQrfcNZXjkr4y0MvPhoJTegqdWVuobvseQ4ApRA
MQdPGSNJhdeQ63hGnX8Rv2vKmdjVPGK41t1/nYkjBIdF1pLpCvE5U3kWio91F5Esp8GSjNlOC0cn
m3l9QH4hWZCGNmxasALN4r5ixcy2VxAgqf8zkD7BaHXiN9BZmxTGmP6fItXGPsIS0VccJGyLHmyv
YaaTneF+1RW3yx7BOwz79iNlNpYRjwB8VmTm14Lj5J2Ifh04hY9tN58kywwuBaEFIO39XOQDfhoq
Xy770fmxkK+E3SPKKwCmLXFI1OZ8XIviEvP+pN3pZuGWn2+QTKE4Kycsn5qwBAnPBVuQgAs4ZV+y
e7NchrHucTsrbs5H9MkertZpmDAHu4jbOSrJAdwpt33ESsfT7955HZL0hL0BHzajHwVo49u/jZSJ
zaJNHJSPkr/iEkjHDHynEc3LbDKoHXUKSCsaI208BgKGdUb8Z67r/g/WM617yDi141Ssd8J5EIcb
ylI/JI0ondbwaeL2Ns6cBTY/U4/KypUwAbThzb1OkdgydddG0PiJXRnaQqHByD1c4npcjaya5dVM
nAYak4O9NXRvdPeluSH8tQvE9M8O/dYPvMHnpItnVDDmH9rQbBKRjG87Kk7WpORBRvSycdj/rkOn
J6iLgTpZ/5sI0YKEhxIIVuJ6JyB6ySmj0BSj6WTR1eUNsWfFWUJaFMYH2hxnH+OyBYpUea+HweLV
7yJGSYgc8HjV7wzLo21lR0HC0MeY1ohv4bvdn6MscV/ZAU2o0Ka1wmccdGz5GS0lEjMun/hKl4vd
HEYSuhwPZa39I97R1YYlfdAOA9LgoPxITnBMg7phw7GtnD8yXFchnkCV3Y3hesZSqzKNGGP/zI27
rmNYKYc+4pYhuZjDD/CRV9fvQG6f6RSK3hcdHpDVw8LtxukEnDZFeCLih+5ZvNZS6EGdEeV5iv4S
I9Xc+cTL1rVO6d6ZpAuHIQOeRr0ryX7aJXNI3YyKJGQcqFmC5UbnJKI3j4PFVD9c83416tUfx6KF
Q2a67nwM9CFRINZ6esMrXWN9Axal8CCo2Bjh6hH0aGirSACeYnG/F4+C5GGrfm5tOk2Ijj3bMgEI
J3Q9q4gsdCJnlGbufYOyrheNM1QrSmsFJ88Boekdn2uhurcRaU+eMNqkZyOcgrC3IKyW2a5UM2fb
zbOrafvhi6yXVYMD0weaRUynPL91QfhhFkJmVti337bqVV9Q7+8JF61CfggtyZKyx57/583dC6ix
VsArE6VKH1OYO+OBk4IVu/8Vo7ape/NDrPb7UxvFMo/vfFjgZA/5v6P/4pSsu06qfeCg68sVWhPz
CSw1SNWmzHqNxqF0wih6Bo0hl6FqOBiLkVEIxrG9UG2xpvb8tB0CXHwP+X2d+Ic0Ns4Y2+AQJrcW
ZeSFV0DqZrKP+UiCBZJqgfZWW65onljyBuedUDXql7wdXrksEtXX4unKpI36Ietg+KRGU6cOKyKU
SPdHYG0cewPrNu9XL+4bdc/J5Xm72aIH93QN5uKLpJVQ9wrCMTpZRabNWqc1Wnyvbnos1EVykHI2
CUcz0Lf7rQYiLt+uwfk3R593XsVgjgKjCBX6E5GH2CfGXFoCd/M1JDYefwdh1E4o+XrrGt6tzYOd
UYG+q5Eegw/JlRc5yWw1nSdjv+iZJfBZi7k8d1FlpadCchSN8w/VCxUMjhRMNvUjt/0NUGe9Gd83
C50LeLbqi/GxPRRZ0rmTrrf4mU9cfoYYbkgpicaXfO4zm6ekKo8p4DT2VvOQMPDfAO90QNNQWZXI
D0xvaL6/0uGiDXVdSrQYe90Yci8mf+UijMh/BE+al59qw1H4EW7OMCL/FTAWujDzKVm/6pKgmm6Z
7eChQuKJ2tGutVlugY6ng6mR2Y3e1HfYhl/BkkCgMnYTof7puzR2DKgaTwf8JEjx5tqpJ5Kwjh1i
ukX2d/K61J5ilaMHV4cB4/ggdAwSYPGts+7Ro8q0AJB/AZZclF4tKbS2G7k3TCRQaUpA9isMV05V
DRGHtYFIF/jKwaQ+IGXY0bWkXzB20gbNTqTVo8k0p+3D7aC0DQOhGMieJn4seSQAj3QmIrfnDBqu
ArJ9+aiUXF8GRIxNiG4f/fO7BFTptv0jz7MuwfLks0y4/UT0/sxHRSgvH2CEBgLzwsCT0blw25ft
7k0n8CmobuSk2dgt3HaxymwYH8Ls8rfyMimb03kZmwwZyyW9l6qZEGIubPPB+8sWF0OiXteU2O0/
iYkxhKziyvZY+WL7IDitgYF0/UeInxJhL3Iz+G1xnweBVdBV3RaiwyuWFGr3i7RxBX5LZdJ0MZpp
dtqUtpZgrB39VWklZCdHeKpywE1JJ4PXC8uuK/H5RM0r5tqSdXzBXk9+wyn5pMOu4F0GJ5KxNkTY
qB4nlhJ3F1JPac2BVL4y8b9X6Ed+rO/FSvAVvN27CTNWmI7XKIPVQlUkrBKMQ0bWTCRbScr46JIg
x1CYoPknRriUhzqCO3fTaWR45XpHZDpxbULdqQhr62TmNjbqHlgycJ5FHhEiei+nAImr5Px5sGEq
g6uyC/PX687dY80TLqLbNYKBQ2/fnaE3SI7OcF0H4X7VAGB1FSiHWOKW45ag1YGsrVn8QIjZKWOq
UaV/HE3PJqT0D4o940f/NQ/FfdztjLEKk3gXu0+le4qYNrdPevHQPIoPu5FY215DtRpricA0cGrk
l9PoAskgHI7GPSgJU53UMZ9UrGQZ3IY05QvwvpozNeJszl4hGVphnXFhg5ZzXGZf9qGxgvHEyQB7
0j6TZvRgDNos5FSxvurCZ6MlK2C2h/V+ek5ztplBxWFH0kqMF0pMogmP1uVuvMOImQd23bVwkLkX
bwUXRDuSm1Tf7EsMIiHbAv/nX5bLZqWNng+av7+j69mvZQhYft/Gq1p2eVOzbEqF8yKIW7qUim82
GI0UkD0UUYws84yBosP4LcneHnzAvmEaqa56wCwiUWk6cghZ/aON4u0C9x0RdlN8eRI0CPgkoJT4
dzj1I7hi1vlDXdNNWmsrYp9Ubl7u91KLzVKpfps1RkjndOab/m15y5AaZzM/KGAlY8ARHgMSsC4F
MBEgPCEX+Zp6rIZpeAwRid6GkszIMsn50VG5evn0ya6YOcwZBDlQmNve7lCl03BzAT8WiO2WpoHz
qsR503QdhzLI/qk82E5VMo0vkfQAnOiWlsyi6RaaJ6ByLWDWl8JOclU/asHoLf6SPXMay5HKnEbu
SG6CBnV4r1QiEAfhG+YayjmpYQAjGoW0mxfdmOv3XQhTz5GUAKvNz6e9EChKqbpcmEL5KhQ6v+lJ
vDO0f4nBfSKEqRWkbHIkr19HcXXBYPlTuAaAH+earPdsqkSH7l7jPJAorzNHksaLhBDrIo5uJxi5
0eUfoGgDxOA2NWYi1xGybLddQdCU8ZxceM2AwuipNtJqypcwtR87RQr9cXb/a3719CuM1dEHBfII
HR30Bq6H4s/uLzyecopeSbQKgha+76oyyhxIgM2fmtjV1o5kYvRG500aqVMKdPCRP+BgaF+yaoRk
6vNoo/DyLKWECs5l1qyFMlfZVehzUKedK944KkXDd5Hmph8+A6ryU96YJPzCnv06jM5mlrBTy6EG
FOKD4qNlKvOTck4of36nO4p2RrxWGHxhINcj7JFSMPYC+yAk6dU+Gjz3iNU85vcKgoeiJPny3+aO
xkrWyvhUvtK90ZTIVxLinOidS0roL3a49QpFXlDMZXCdyln6E3QQ0AlwT6Hp4LO7aPkQMToXnWRb
vjJgyPaSQISnKynwhd6XLqLHLiX3xCIFwdUiXOpbPv0NagB1ghLuFDRdh36ivbvTfRTstbCMbc7K
9lkmtXro2yZCnjrxXi6XNlVbuVKCPKgd1DZ1Kg+H2Zjjo8K+gKTlwOvpx60ftjkksWi7sZ9EmaF/
24c2YU/lYUvWOhjIQes+OkCW9EoCntYvlohZjT8Kqjed4yww65krfkRuZMDkzhuaUOUfj821iXUz
ckZiRTiQ3htRrsQMHuw6ix3R4KuqnPkH9917eRaHm14StVTndaWvagNT2+5F96afaM17jkRH5q4h
owHtaJ17Zkg3vY6mlLuw/e3P9hjZQEgh7369t9lludTp9m4CxijqzaD5Z2lpJy/5Kkq9JLYhl02C
FwQ+ERkpB6jslfhpZMII4el2d2ONIT4Nb86r0KOC6h1PPlyYm/spe25t7KUW4tBWbGeYu6xjiTTL
qITht45Q/DSYH33Er+t0u/Y+wYoOAnsxm9txLoUPjKoheVAVBxAyg6ttxu0P3DMrYc36pBbZmEWw
PiKVPoI7ebVY0czLX2Q3064vWmW9LEQjEINIQDxmsltw1AhO1k+Cxp7Ki/uXWaGxYw9YciuBANT4
otHYqF81WrW2a57dJ7w8IUoKCo+SfQOiBI8bB/d3B0Asr8m7pOWVbEkzgVTfZ37tkiIhRXLIBSSl
+vVnBFV45xCI34Ba81eTh7s/fNrgHveASdC4X/gPo7CYp24N31+401i+YIhBYDg1u0SKc84Hmbj0
WM7Gi6M6dc8XrYkHySh5DGJg1MsSqVdaw7V64I66aVnCES/8axzWfbV/YmRVCzXEngi9zXhgnndj
Z2dkGEbUCaP01eTD0pu/+me0pRVw7sKIGVgXDWYNr7HHS0pPhuE9XvLjDCDVwfxNfkMdZmsNxf+h
syzX8dqdmqoOSW3k1qWYAMGafYuJbjaJpEU4smhvveFRJ/4fd25eyzXUh7xVn5btJJnbO9k/9mDn
/YEVauUhXK7x6QatvE45fgTcRqesVYUehnUxvknUjsBW6ozxhD3IfV8am2f6kA36seGpmSaUzNzN
V7GIU6jekOumrouibxQDJ/4lpMcqw/CeY40YE8O3L+ARUDW50Eq4QvfyL//x8DTUSXpZb/6o3B16
YXp2QW9AGGezS9yTYM179p6u7QwD6ewvBC8gQdiKGMyH7HLFwKqGouq10O54v5TT85HPVzW0MymW
SmvNTUx7P947KDmVwissQ//Xzum4O6eUMXkwdoqaJNhmR0PvoRQ6DYC+Mr4t67CgilBT17xBmllH
NRw3o1Vlkq995p6umVDKejutDXCkZypTcy09f16Oct8b7sm9Ar3oViuaz6w6lUQe+8l1yxSQHk0E
9Akd4Jks8PAAkuGo0jSnFPyKs7PLegMDOnHT4/6obgL0gM06icQbLYZdwgJ507B6Saun08sjKKf1
OVnx/p6tyx+zIm1v9p/D2bXpz42YDex8zprD752gshb86GhZCDh/QlDNT/nB/VeAsIyW7SA/8+cq
u56hsPTSCpbZzxhjcQbVf5eUzI8/ENP5o0CgHR1gCNlVdQ7HUg9bybFRModzBgw3xgqGysGroRf/
DqJyu0BF6lvx34xXqMYI4a8n08JJspzQzzeQaUzc3pjjiS4/ST60gL+eFT5YxXlCuSEvfu7/YreJ
K5/+IFQSWXzxyx9udMsYxAeZY91vn3MfZoEXiAGfYMP5NneZl2S35zy/SjExzq+6r2hXRXRhtAqI
k1DWIzOdVHHFHormfysYUdmpBpENgSmKnFRlFipX5bSzkKtbLNOGRQ0pyEjhZlnjUVP0+o65MggX
ahaPQ7tBtONm+BUIZOfnh4Qtxyatrkw19iop4FsRuPiWSyaqEu2a9q+nl+ZubVCq3YhR9Ue7JPpb
cBddjlSzIUNnH0Lc/ymmq4MhwUzN9U/5YZUn+uLdAsZyidaxpLhCZ8zMuRICko/SiaG4aOjHCGPl
ZbQAfxvxhRso7u60xQ3AWIZOCoW2mSWvZHAsBK2FLDkjMC5LN4PFhq6ITvih6DFQ1i/20C4hKJpa
CL/b9KvHh2se3Qk5od7ARg64dzvX/VFl2TX+CcNf7KD0R+XnxlRIO9ETQPeQKKoolRf8m1aPS2WZ
PRP9P2oBvPDcOZbAwUnZbK9FadpQYHifKhBEQtYDf3XtF4yn7cCt2eduibqs+jUJjbDs3lKALaBJ
9MJT6l9agwYnlHx5+HiAhrknvJ7yeVv8IijPTa2ejilq0QMGxFR9+EzIWlblK8P2W+7HF5cv4kLC
U+0OEHphQgGuprHe2d0qrnGf8qtXuKS7c2qlZLzgx0tdYZyN10pjP+A6vz1+GQp3+gsUbTXcHZwZ
gR4A5Wg4trIWiCje+GoZevAjroUkS3b3xzYD9TulWU0ow3fRfdKZgDVemp6rkmjmwoVZisIHm7HO
VNup/GqvdnCLfg3ImG2+YM2jqqM4DuUefhWl87yOoKEJcR4oX/Pff0kK+zQqvkU3pIFlS9KrUiWq
KsKWJlzAhtJlIlBSTu6ghHwohTclmEKOGIHgKDFdqMo2o9gXd99SfAtPYmMEufyixnHrvOFvnNEN
AIpHwedHHKiyPjfcD7XumtRmOLalNxEgFQd6amoIPurz/PYy7nFSZKtVUwqVxK21/U4Ekh/kMPxX
7k6H5a4iwh+dE0l75H5M0MasugnOlxC24OH2sxFQPf5ICR6s/30pMkeohwchPxEcTdIk8khKS0v/
qGTqLo/j5Y2A28dkGkfwzkToj4xkIU/kRX5xvqIH+Ud2jA84vmdhKtKj/+LFlLyoLEteLyBR7LKW
6PK/LheStRU8Y3Trd1S0FRdDdOeTApylfvNnArU8ttPDt+BlM8qwORNZv4LeKhLUqwUeJ2Ehyc5Q
7VaP0UH4t3jcVv2NyfGMdCZFwfOj6ZtQe+CDtC/8HD88id7dkNv73GLEDwHsXrQEaUmSvV5Q47Q6
GcG8UU/3fz3Hj0KfkdjBEhp09dKnovi9grtBALoPLAJ3R0DHsiVjNQQkVIFVKd8rqfgJiuAL+AX8
5tIqbADFq+OgJVeFUaDDtI73zE//WOJ62GdhAhg2pYR/lFvext4y8Rtjyi+R76CD+ALD/+MD7KM5
uBBezXmYvsusl6nXRMmWOggR6WLIISBhTITZomlzYRlgslsso/kx2+xDlNtZAUk7WKJhLCN1PFSV
unCURvCMNqM9wnBi2VddktM768KmpN1/Bl6aYknxb0tKDgyQ0ppzkzfmPoQmzgN3/5kpJTaFRxjF
eXLZaMlhgwDLIj6OVqtkNAtHSBGm9IC6qQLckc3yci8uBQlu2bUBHesO+6reOCtnMgpbN5Yu1Njm
RQBOr1J3BoL3o4Y43TFAfWS9xdjcc2B5OCNq6DBRJdXHquH85ENiMSn7s4JeqqkKxrsbivsdXid1
iHVeMuhWLOth99wTsA4GNT8o3+ivMvJot4CHlHJuXOjC6sUEXT7AaZFvygi6ABjigxtD1iLsvFMh
SvrkUMtHDcUDBTqP0Ix/9t6QvdvPmj5sgeqq1JUhl/jRzu+hQuPSg+QtCa2WOc86UTGkkoEyHSa8
wBb40rJUei/1nZGS0LObkvkWPafT+GYMjONa1dW2IzpPe43QDV4e1vx3dwNZzAImOZZpBAY65dX9
XQkEOISsip/VCgXyqrQkSrNsWhdTb6HE9Cl9rVmwlA5f9lBekTvRu8j+u2eCPhsNDMzSp+SaySfY
TXJym5Q6GqU4t8u3zhPMbR/JLMNLeRVTEAMi9moaWvLhB+TBVTon+lSBHlXdWl9PD6UlxqohKZvd
+pfnmqZr9Gy6cNWg+XqjRux7zKFIzvnKASILoQLFBHqpEtTt+zPHQZnchSPZB2qAOjJQO7ZEGcxb
Ne2D2UsPBJ4vsjHk6xKuzF4oWP/eiM7w27gzNpUlZziV57l+C+Z7p202M7zEWAMGRlRWX5ihRhaO
KEvsMZu32AaFqDwnZSMzHxwY3AUGsAZxvO4f7KwcUJqsdxykaYnhtWeODZuiC/5n7R9+KuVvwCVt
CerREn9451BkHO3fdXVCOJ5bFmdxKqY+ZOaED6gaZkYQsBia9+CaPwxuIUs3lZdehNhzEajJG9Du
xCyIg65PfHZoqkcPZv01CqTfcvdn5auwy7KLfwN+10xK521SGrIbRKWGhs2Hv7ycYbH6MKpi+938
fv6EpqAf8zrAn0G0B9gKxFofz/1IATk/t8o/fxUGkzMsWVFBFYdGUjStDlb4fzHDBjTaDiW4HxXe
BP4l25Zw6hu1ZV9cP2HXDSDKJvnoqS85cJGK6HcV3DQ3NoLAAF3pahYX3XXIeeK8Y5eZEp6189pl
ZQd2tifotjeOD93rfoFin27pwaQSS6Hqgv62p8zzkKw4Ryg5YdyYkDKKymM8S9uIMHw7/fCyLiae
LyCLzX8pBqMKOsO5QF6NI4oGQ3LBBoEvRSjrdLzNGkbv/cHcY2FylqFb62Jhv0qPDWvShRSPN8+v
I7sG+WBBkRXFkWvCj2k8b9Kt8wg/tI+GGRms7nUdkxF2IsnHdYEI7Wjf03ZLrs+blnGyE7hcmC/9
9h5D6t/DLZHiP3QPar/QuSGYiz2RDYqp9fpxXBwZlKJyhlUWZ2T4kka460KnP3JV6WoKe7NfYCNX
Vd1gNpO2QWrrSE+skSKPLh+pc4oGQRs5oW7cObqXlO04qAriEZD4y0jBI5/wXCUoO1qqWIMSAO9r
5Vcxnl2MyHw8sQsTHqiuQRMXfxE/5BD57oJilR1MvKpf5AjVO+Gynw0EtBfyzEAInwLhUZCWTDZ3
FX1WHt9hRneqYtNoeTZ5dVisIRbDS7BgotwcqSj3ydaZMzzBGMC0RHL33ZJtnuq2VoaGIDVm6OZi
NerFUMkggiO1bE+zQr98t+mXo/9RM/dAtzAyU2kdFVmWQObnNLpsZ/71SEyMRCHllrbkP2zJwTxP
U4YwNwKH/Je+SNfPg7RHIbE81mOYulQLJBAdwvET8cKZo4piXA+rm92CNZTbh271u51terYFg1rq
FKlRpzzg3hpLGQC8FxdF63fQhg3HYQta/owttBvTVHDU0XQqyQxKsXLGL+On5Nw5qFYFbnG+pSBk
F2YnKJowQ9Cxygk7NGwJfj1dorkRrEz+9gM3nZAIHid9I9oJVsnkhChzkJynbVH5I1czQfIMNvkA
2yXgZHPe28E857eg6X3zD9cOlnec0DfOlIQwXbtGl5LcbhG4C1+v1ii8w8bZeCf3huk7TK/J73IZ
+qJoGGhKYom1JqxJFRo1Zf7SLai9xyJFbDaFiDMRsMsCaPEWGBoGgAmaOQ8oVwhYCbSM1T2wvjv3
TXR+rZ1HX+jcb5lRphR6V6diQBfjMdUGfMq6ckNF6L5M2CvGoGXNyDsvNiqomeu0W4cnq3TvnIWB
kIrTdqT11STXLfV/zURW4YhBpzZJ4mInT1x06JV+z0wkuAt4QKpd+yDupAm07f7YmLpP6039hctz
UPPymVUvYHulIROlMFVCwhnGDo/OERsUvH7gF0voGyPQZNvaCqBzNhsfbyP0SIMu6jgZzEM5oCZ4
PXcwW59Gm9dzIYxZ7J1p9HXsUB8PhS5Am/RQGEHSSKgNoEqFeiPif85Wfm4DrWjKM/BY8iK+NL7W
B4dmAM0PuitGzYqWjYYpVf4nryS1DmQ0SH4Z0fTWl30cOcq41lpzsbTHaR6dONQJ1ZZ/1BYZojgv
T3ftuxEuarXfZTigzHucYkumiEL2vGj2dnO/WjXXVjJj3WuvNcvNhSDTZpKS1Douj1nEGG+5obsG
bLbEl6Mh6lC5HYhtXAgUqumxNAmmw8DU8onPYinslyi93B4Z/EP0mFxCe0jr8ZCEViS7OBk5Vvfu
qS9eauDZr4ZoNxooQ82qo6j/z8IFwv0xDLutPDHIhQQn5zvduKkg69YZKd7oUsjaQsHOoHdv9WVj
LRuFwYjjXEN16N5BZjMIxWNh15iUDPXZ6p/CkvDuwRB0Ba7fsg1K9PT0lMSoO5A4F/2r313ddVI9
wKLwaePFJpaSLCNk0JspEBXqvZQ04Ua5naHbZ9bB/TIdE1TwU1FI7BJAhi75bo9To8dIULGBRxNT
vSSZswjg/zIe5fYFHIK9xLKY75DgPVYjwuXuZL5moyxIunAEkuYdencHMpKWZq/GKuH4P05c89/w
jLqEEtvZSvIOu/uhIkkubdcR8w2vO7ELX1JUM0LQRMWLfnxQ7/mF9Hs7LjL/P3dvWj67Ggc2rwJz
keR1Csl46MdqxgUqPrM+bMHb1InyO+yxxCFEtOS+t72dlBzUK/j6TNXpCgVor/6GsQL4XtcQrS4T
vyROMoxtvCqbooF2Kn5GDXFjitWH+6PT79qAKGOt2cZgWLXIron1sQ3OFx5gBeeiDeOdeJZuzOwx
mK/cof38hiZ3CVlRyZQzLsI7G4Ygl2doI4JKFIU/BxQiTDJVI1ZGGGpjIXTv1iAgwzUaE/wZPVh+
DSl39Ke99xnR2LhpnHVuL8LBVfOL9fWQBAX17vzu9zQNCQ2CFgfO4advvpz+JcZ9h+6QjoTc+SY0
a8w2FUod3MqvdC+TiPjkgyayPq3Pxmp3YW9qw0gHQfJKrnKgDmtwWbBjVsnRSZD3Pz5MCO3kR5sH
7RZs7qn+42EZR7pB88bzjWtdSayA63TNbHqIqpg1P6wmmBVQrhxp6M2gSVFXbT7QXZx+0tc/gZ6O
lwZNpyaTdO24ORMeUnBR978n0AabzCh3ozDohmJghK1dHNMfYO+hqgUUTdFPEcMVGjtb6tsNLqZS
mLeM8hwgmyqXVjrIqbmwmT5qoPuHI3mrd8Xom8b2DH2WvGJ9ZAH1WWTQTSYqyKbtu+5N5Gn2Urbn
4A8b9cBe/A+ldvvg+wI0bltuNehtI8lTRgo0flf0mriLvbKzVSS/RpPeHG1EwIcywp82CBGf1TLW
ufkjzKgJamcRJs35N6xQ2ixyJh2j/NhqB2kSpS5OcmfEGB0GRCl+CTKlKqi5U2Dvmi+8jhg2nx3K
BuJhRoixGaktgxmAXFDxzSSOqsqOx1W79Ihr+XzDr4yotWHScD9Vlz9jbw3CXaoAQr5DuAQV5mfg
xxJC7olLlBBvp0JYkaUTYwa7dmVmV0vnRw8Uaufhi8sKN7KsJR57yQNsfjRnI7VaJARCCxI8T+S6
NJIVX/yBo19w3E5YP7VSx0BEL9WU4UZc7GWG5lrLnhFPt4BuLPbHcyfxmDuWBqAVPRjwxLG+GYD5
rv+fTdcRxqXASpWXLC8NGpkJS/8qSNtDVTev7KIEN4+qIrdG+AafL9W7BO0fRaPp31mEDz4bKVbl
gFbjl5Mw3F09765vGH55UGTx7T/KC6qEvdBldIfNq7M0qqzSPP49bM3D5eaKHPjKTEKua6n0wEch
zD9ip6mB+u+zHMyua/nWxRKXrTxVl0PGTqXQoAkKoQ7ORK1d3e2JG8BodHPHxyGydcP1LjnnSQ8m
Ze+A0bXBKyysrjhwCe/9ufPPbA/U6tk9Wo6N/JokjUH0TWMqb9x5e2fVjEE66xrySEUQHnuL4v/b
ohVLhSDqIvuzXXuaed1uwbNe/yFvI/R31YoDti6OAVwcoqvWLDzp2TYb3hIpIFXdRIU/fBCeZ5eM
fIsNYYF0L8k1N/JJSX1Kgp1OP5r2fEl0pEtOLm8LtZV7E29Y9XICtiTmQNvJE8ncQj7sUcNdKsQo
TkzmaTBtkzeN3REiKOAZkflsxv1dkHtRXue9DU+FgvULtp2wj+VqMgErK9SK7fRfUZ321pp5a9dA
rgnLQT+ms5+z2fSC+TfN3yPmBqyh/ikKmhodU9Awk/sYMSsn5DO/MxP+QkU7N7bcAb+c/scNkzYY
8vYQwxNAyGOCietS/IwMwsC92pa3hwTgZKYRu6rKjcreEkdhVbH7O/fa7poWuqFe/AixhGdHwxNx
+p6nmemEyzHBFQzlPoDGc0BJot1Y9x452rp70vUeCfAY6AXJkVd9d1bo+SbVtXMPLcscPF3VpDi0
NRpKwubN/quPvAyg2VOLPYX2pk1c9ySKoiVcSQ/hhxG4dOShOlp7RMzW7PXPapBCYd3U4qkInitk
EquRK/F4L2RWlycHLlh/SbcQbKhR6g89L5rPpzld5ij3YxUgxDqB1+LnsZhZ1HLdMGzVoOx/yD04
pvBEMOWwXi1U3AxrmScyw9GPZuJXVd7bTcNi3ncddVApmh/oML74e+HRvsOBtittU2Qq5EbYhg4c
X1BwALJlpkCnrOmiK6nFkoMtM4xh7wccDyZJTWkZT/D2JKVlLswfYS1NLIL0qqrzXZfX4cW3XrtA
sYQznSmUp7VTpYeG000i7Bj4/M9YN1WGvigYbYzdONVvNNVwMaTQRnPP75tWsizBq10rA89aWL8z
h5LNLX8HS7TNMhgFmf8hwKu07XpfKJ+S3HQmjKhDS4475RR/iHSM1mB9KUdvTaI0zHda4GE3axP6
H4H7HI4U6rgE6MeG1Gr8qcS3XTHSo+N5Jg7tah9W5NfrANlwfVjG/JwyZE9yV+JoaoZhSP9v8BKR
gIH09Z8KX2dgEbUUP6TWrDeB0TPSaWEUHxe0aQSDzzLueySsDXexz3RIiglelFcoMkELQ08DlnC5
R0u75QZGb+28cg6BOL44sQF9xAt3u4HCGkfmYFCcj+UQCoO8IAtOaA78BDr9XvD8Y+O5IGaPTBOS
bWnwnGTHqP/SXaTME/bLzdvALdZgNDsyTlxzzbI9Q3PxzxHqt8TA2jEldLrTXLZdDDAUry3jdWOa
gAxp2ktWWazAhonNTrgF/mhHmfvEaGXZ5cpCqwHDhAqLj8iJ7TB8O5nKhX4pKtArzoPRSnOpgAN7
vXiFRP08InoSrmKWbv7an8n7lBVRm2h3LhYGL8SFF+lF/MlusaAwzokX4bYV38KXFPgrbAyOPnZA
sRb0Bx3d3BojXmnPzzMYnOSb96FoKVJ4wOJjaLE9vuQoWo8ioyZJarGGPhx/GAGIyamWIfCMmiCt
DSnM7vRIR/73y0f7SWqaZztZ8oJX8PIjuYwgo+CIEa3IEyEYuHbZkJcZ1WM7cIvWmY73rca85EK2
s8+vkMCDLV3kGGTGu0U3cPlPp1VNR2TPyZXwCP9mpGnhoV2dU9Q/ft0YtmGvMhJyxtCpdtRZ+VEi
xR0Pd1denZ/zSXVVeRQ/1Fn1blcz3barq106MpxecBC34njs5AZCa9I/WCH4gdQ+yDVnPNEVhLMS
uQOEu40loi1rYNkeDk589UO1nWPD4tpU6o3BQPDtfOKsqNwiI2fZV1HXDHK75NKG5vJCDIHN3pAs
w70y48fV0QJmQEmInZ8qAJf1LZ9xu3so7PYDLNaZ6bckZ5LB3TDfBbYK1IDQ3qSz9OnKJ1sVl0RU
kniCkaGnkK5CV22yXq++hkfsweSSa2yt5m4bD3A8I+Ojk5XXOcM2qj8jPEt1jDxVRRyyaTDb0gTf
Pb8jFBRvxKappYV/v3ke1NXcuqJ1h7NpKPVMAw4nLJZUh3awLCtT8OK0Vdac8CyILDHGJT7qOGCJ
T9/3RzU9VGiOqodLzV29eO6zKdYWi3Buc/fojfUWVTDBBj02z+eZ7OEUwn+wmOhlMZXq8r1wVBNl
ZRokK1BDAAyBAb/PDvdL5agCY9ij9dPe9oPQYCddbvTBLu5K8uSV3c83ybgzCJrkcxBgiUkkUkLI
qd6hpoWf5duiKmaPpFwMVKGsTbifF2J4RxsJCLhtyCA6kr9jo0ip6rNB1pYBoveJXmKUUpHQzYVC
GQuooTrDS7P1cztryR9gnAUDpLn2oigqRqMSfdmU0UMjg2B4SuN+3P702BB5QrtujlNpOEvANKdd
4PlyB6+GRM4SYH3l9AOabAWq4AA7MDlsOVy0fP4fsW0u61MTchOoSImqYd9WFRuF8m5nqpM2PJoE
aTOkwF3opKVsTJ7siDDAkGMUnO6EWg2dLQcVm2JIl8JU/nU0INPk2joy6YIJo5375BYgkKlOG82K
kfl+doVYVOli3lrdb8uRco+2NozQlQhQpeGPlLbQoAstLNEUmm3SnRa9YVSodDAHol4zxKs0QViL
o6qapDfmK2pLLvtzLWXZfg/YxFIaXhvhFnEZMwiD6UQx+ZjHak5E0tL6Dt+10NQoomAQGj0zFC7O
NdkOFMIenrqsd9AspC+xkXU5jWvVZteV4RTRppGchTMtbRQZ4lsCXVDVV38z0iOBDTif1y3j/CTx
uPSgDUAuezo2dw/0diBmxjBixYGPJPtx81a1y3XloZlHlkbiVj6kvRCX4d22ocrRdZGPcTHdNceK
dHV54TzGPVuSXw1hFHW5icb1xHXQG7UeTQF/Uhhdpu0wumGJkUys5LYGr4wra4+fEYb8SmN3ju5R
qC50ZmWtl0TVMhMiOHZeD1O3NEo85wY+pbqG0w8K2e1VWMrfdzLm6oNg9rR76wKtk6P6yRi+ZJWt
uRj9uSuVy07MT/Y8TFxPcIvQYQzD/zODhKyvO3/DjTocJBD/JlkjFDfEKURoSpX8Jc4+PvQGMlUJ
/LBUdmsDWaFEBKvzAGprARuhXKZgr9yI+IaGuHau6VW6vYm2eePSy9mHcUIc5jjzdcHNsPK/1eQt
Cu3sju0Z6ry64Wjb+tiQ/KKYlvP16UHAxQADMTygl+KOOdZtHBtTkyFjmVYvO34WUtZuZRnOa4L4
heta7GTgQKm9XtESEQp6yBCJOJMEdRd5LbOGBffQyWxm7fX/pfwbbHWJIWbhbXB4XRj0exKkCkDn
UIFbas7FQbhRonTOD3smNTm0NqOefJv5MNZ0xY79bhNzAgcMqc5Q2xpQtXOVuWIDQBbC1tUim/7L
KN9XCN0Md59ndUFPij9vZ3LIC1Z8qTdbLrUtFlq0vxHH8Ny/nO3j9+VzaJAq57d0iud6V5OppMLr
BTn0ytDehGrR49KIFODUsHo8TTP7kZphAgU4g+49tm4DUC5AoLiSJ25Q6Zq0q67TmGUdEyRHUXzu
lNmauxTPh/j2j8aqLr1LEgDmD1EnxVq5mgUQWCAhyF+i4fBqKkeAzY6WTFW6vpUaRaHeGyrQi/DP
fl4vsnfiNKf4uZ0mG/n1MUy6dXJMleeT8QnWOxnvPIgs9P6x+Vv5uJoGswcZe+rFGj1rNe8uvTC+
YNpC06g7kpudOYFwVTB0HvsHUysTOo9O20a+1Fok1qV3mqTIg3UtH0vc9YsuW46qHOetFNzutL2m
S6MyjGhtJQohJL+rQlI7ZfbuwRqVPqmJWAlAAaUu6SmisYHz5LX+EV6EuqUY42s6BxgN+mpbGIjj
uQyfVGL5JJAqhauKHGZjk7p/M0/DkbwHaqWKWjX4TFB/4xAr/U1892SjFBtF0hvqVAa0TrvkFKlL
TUGFLk/RGn9n7WzuS4danGZ13G/kI9RtwCGZi7ypVISufazXiqkR/zxcGtZDepVCDmCF+C6o4WSz
X6pSCP2x7UWtlM1fCTVeoV7saNyM34G1LPjrgcNE13DUk8AwGtxeo5dJymVDuwVTdQZQfMZFQTyi
LU/LGUDPHnpVFxBX3YqHt19EB+8JWbVoZfYfvyfCie8orsDiYCGNIjJW+ohjnDkf246lVkMApbr6
AvoC0joafREcJmJv2EN41BWIh4FDHU/rvmTgAmpHr0s7PD1hL62i26BlLshj7eMF80g68zt4weMb
Gt1lr8gDqfaLVd1e8Etz5f5lRkKA2T9mEzarpFfLWXnBRQXQ/VKF6szbOKMYlFxdfsYvbd6wdBWD
0V++GK5C3jBAi5bFpDoTrjNcZy7ILQZUMBn3geCmA8i7mFFp2Ddt/rnvGdq5XvGfFxlR/i91q6q5
VdaTx6EFmcft/c0lSNb2zKIC2zFZGteaeU6VbqFR8CE4v4sM1bTbTkVLzLV8K7plNVx6csFMyrKc
m6XwBQkEpk5Ggr6Cs9Isxt9LJXJBQuPywDgAa4Vm6abMP9YcfmCJqsrXJrxNmxW7DONoyEFuHohS
snDo0HfCFuKg3mKBQAQVcVjJMUkI7ki2Gs9mOWK/qgnbsnSXuFVAVrl4U8xBzj4WPBghDwgBDh2h
5xQLu9V05X+8v2djAIempKhSLNTO0aPlPzb8Tj4SaseRy+JVJwDvG00BriGuF1of5MbVzcyd0C9A
bqJJg2wHC9P8gD+b1bE5X52mlihOpPb0iBVH7qkCZ460hLTBPsveeRwmmJIUwAz7/q1bZMPNrAgu
723bCcbXlgcsUpE5SpRrZDBy2cNHYOLQMS94SsefxHTW6SqsvCYGb7GmBC4/NKMeGVcsqWS0f6MM
tpD4EOK5dVndMWO8j3rxIu5mlBTUCdRvR6CtSeUWJfsCqROKN0kSoyoj2tOzKlcKXdKdv5p9MdtM
8CgLg19Cx88TdaEL6Vk4FXey87m/ZDCl2qLgbNTyDjpuFMAchqTlsiPWLOzt/KyVNDwdR0FHdzfZ
fC+Ymdru9vNcztLRyRnzWin7acSgkzrW3CFcE7mYWm7SUnFx+p7WjOKOiV1NIURvG07sH+xmwgvT
Oa2wrCDjQh/p+Cdx0ov8qeAMxlmcKK3GdD+EydeGEbgIcaxZKKdBR/vEUBcayP4GliCAEJrR4lJr
G0RJpe9fxyT1nqanuchomI09gW3ghQlghs1COagsn7N3+KdQZF0zJfnaWBrPmJOlrxzQLHR1Wes0
2A0mJeCup3XXBOLTEq3AG5u7VVMqZMt6I7ddfXCcEfMaMTQF8mksKspQaMqFgQBV1IWo9qtvi5R8
yfZAdbpG6taCq2J3y/TUqzcjNZp0QC/dtuTrEFyee8kHZSdDgLNVZISz5BuiGRR0UDQ4U64vL5w4
FZuJwyN909tyB5EAacH0rKxAy5qqd90oEOIcTMWEVmtrjyHqUD77XN/jJaSC+aoMUmD1KjtNRPcZ
B6muemuiD6dG9odWS4+Mn0dTebrYgyWxCAfJ3GoOyFgoQ8QoeoPW1v3luR0GztVoTbq/vBAjhucu
7nszSa7Utnj8zi0FDaUSca9EBTKInf1rkGg0GMgMvpsdfRPlTBNh23Tqt66IiNg7tNBzSWN5Dj3L
D9NDsHwDqldwKC470aUeFkFZG9hSGOeqPKJylSRFWCyUFbYZ2fpPqGlw4RRwGG71aiEedbEVveqj
vL22sChDYsee+aLHVx0Ok34WoQ2Mihc+jDJToTfgcIVs4OjPImnnrg5qL9vVblbH1gMfanZpmhhW
VxlnNFzaX22umE+N2saZZ+5Czewd/9DnpFsRfa+KAE1j1A/GaEELNMcRqh/65owOV9liQCxX0HV+
UC05IjCRPnPJATHuNmEi40aR85pvAKHq7A0C3/sTH4OfZRqL+KI2sgPDJlNGkeJCNVcOQJCVo+VZ
ZS1RPfhDTDxZkyJLizF/nMSN7fanwWrU0qiO8MiM1G8VJjhDkIWQk9eHKRWx+cSx7JqhWaiNSD2h
rR9i0uIPEZeHa5SfH7rtzBZtD92NvGFJ9VVvYEPQxG7zq88ll6vANYEIgnXCvhzsfv59fTw5cZhI
xgeCDLwZXAcfpfni3PRnBHYUl1GJQ/Xd9Rm+QvvUUIczF5TCziDcP46j/oBiWwptRirxf4b/Ey92
Yx5uHbhamXH96cdoVVUny1CSBIIrcO9+af1xgfXSqiOL3Ht1nthZSmNknTIeG7GDP4QSb6OC3Tf0
E1kAkjjnaeY7NuNXiRU0Nfq/0z62IEdl67kxRWaU8SusIBT94yhobaTw4Fl1OfBSl14KLIPN1BZa
ogicbuP74Nknx76qkBWC8b0FICHcrl5IHpUsj6Qq7ps0K2wK/gxl8JqKETwvALbEAA0ifHZFP06N
p1iboD3fpUtlOmNMQzpILwpM7vvvjfv316S7I/I67Vi7QAHodLEExyLj2hQ2UN7NSjnlPiAbt9C/
EAZQGgRVFnvti0G6WxGv7EdrXZNRdIRnmEHXjEo33mOQwU4irofQ6jeLGd50L88S6cZq8XCeK4fC
vuTXhOr4mRgL7xPrQW8m5FmLVciIN06ikWYUEYTH6ytKJvYtfb1AevSTB6FgcQ8eECxfCrgc8XoQ
wDuRpav6yl33jkMJKBdDuC8fezPumfS2gfnQsuhNFdprhMsPF7R6hDb8a1LYsTk6/o3NhxvsR3V3
NMfBS4xPvrcmhaSjP7eY2YKc5i6twhAC9bZVXygop7CsCsopxggNQFV7vh/PHtXBdViP4ccnO682
ORi7oeu3qa3hDaUW15krAslULtaCgzvSIUFJtNrDUcKVdoLMpXAIE/o4FKnL+gcYByd28s417lfZ
X5RyBsHRULMPZdZ9qdIQAXnPEVTEAgz5GLIumOJmdrx3ELVBhreIoLoA/X38UQ5xVK/td5mF7V0O
b8zLzw73NcqL8znsmX8giiQuBfZ2r9AO5jspylTdlq5AX2szsoU6JSchTjowJtL0NuWkm/f0hPUg
tYQEIntg0JO07k1M9GqEhHFTyvgqVsarUCtihSaZPvY40Qe2Uv8KxhfJveo+QPcyEubCRAAkgXSg
iTrhpob6jW07vcfAmUgxKR+1vMoBgY2adz8qmYR0YENERlLLCGU3wmGXTld2XWMX9x0uHdwniQP5
x/PMGMAJCShWXBLZn9AO9SivwScmmRr2bjcAiB9e21reHmNAAeF97M3hQOYveWHRAqMkxUnqsCgZ
CDLcthQLeNc1n+XpeY90FrpZL3OGs6V+IkF5Ku26btPAgW/PBtM1EW9BDXZFC84Cm+IU7OwSU+1q
SOyeeu3vE+qW3DCyQKfJGq8IJVMBFyS7vjuV+oJePALl4ewLCpH1RcSiUcRrqB1jxxUW2nr7QxP7
MsRFN3MWawwdT1l5Tx6rW61ZP/J9RzvNvmooODluvzIxOYl9oiI/EjSCo8OhQIR9LDyheoebMEEA
25idyxozOUaoDCDZUkSkl4Zr6fKdsXXqipJdvMrYwS3ffeSi/aZV6scmRNNhNOd6JJrGnXBlhr7/
86fz8vn2CQKsmdX7k2MCajFc0yu9zydE9oIwhkiYIB6ZvKjPs/Vxz2IEIayA+nzN2wcj/3lTvf7f
v2ncLfFsQMMm9BhSDkiumbUGlkKokPKDwqTSge7hZ1ULb2GUhq7hXZ8rY/szwmh+v6HgFCXfwvXw
Ug4ZJcZw7c1noK0YQ1pya2rKABJ62mpXT/JaazBQ5m6URokKfdzOJnLbvC60tTf6tTe7DNRwLGkr
pJmqD98cMUHErlRY0U6Gc1kYLWUf//wK5gFGXcOeWl5VAf+r6ZEJdAnJYN04HnSZW8v+x0DePEOd
DZoWQ0DhKGW6xgsSSkOl/uWjHKQlj7Q4GPnAAUJjJyR5XuKlZsReWLWiHg7WNla0D+Lm2FUzloH0
RoN9wBkz+JBYFxDHrO1ZvDMx+eP7M0oNRLF6O9yPePFVTy5hiYIFN3jqdOwaASlKqXJWXXlNAkNt
hPEG+eEjEwy/69OQXW1o+NfM61X+YdgpdhobBWau8ja+MEy9nB23kNiacug8gE/scfM3TgJKfRdO
tv4MXJy7E34QgHlgaxUYxE9UO1PwjGJGGiiT1h0+/Fctb88ksehdP9NuTO6SkMD+cXqSL0bYOc1G
nYVWQYb9ibx+EuJnmXQ2roHBTEoQ0sJbMEWfC8IiY4DZT7vYhuuYn82S+FIKgpfAV3zYI0VfFdye
Rgy+6EA+TUr25nxtCMwvFQGUZOSTzBUtzl8i5kT72NeJQD5ljOJYcOKpP56YHARFLhE3TVkOb2Rd
jcOCTUnV7jao7WI1xf7Y+zAYgkc/L89Gk6/IPYUi5/jYCS20nBk6qwC0Fh/I1V8dNay4yqPjC8Jg
sC5bireR3943gonrn18Ne2wERlG3LxwU8aznIVzEDbKt1w1FfSipXcB7WyVzkFq9jlBx42XgHdq7
mVLSYAB+rpp+MX9WS/yIAYP8oJZ7doBgqnuMR2Kki5NMFMsXPylAHPGqPSoKf677IbeZ5OYh1UdE
yNqfIx9/lNaLCci9WQE5ZxfzlK01JwfKPChxoIukuD9pLHp0+N9SYd/nuQANKQ+D02RWyUiZ6OEv
rLadQ8oXOMLXYPEvX2pkAsSN7485GJGL9iuiYai8EQrNOf0XiNylO/SnDdkkf7MF0lhIAwmyHSY4
yaMYPWC7RK4pFcFWiKUJdraOAQl0Rhng+1RuxlBKeSYNnjY2+4VrtRqxmMhL4BGQpRFaWhqAnmlc
907I4l0WXgQcEPHKH2J/9OvwLhhkSpBvMWQ2xH82A9BIFUqLQpCmHf/w+TeoTxcnHuLfaLc8Hbag
+iJhVCErFamP4Ik+buUvJqm1whN8wcqFexbL5CBk1+gCbaCfhaWhnH0CPiGGGh9Ytnq5wCmxmOoG
/USsBihSWWquhOmns/dFFmHhKPUbfU97hBQ9Es+klEqTfdoM6RtGWUy0QEfqsLQFjvstp37flqhl
EEGN0AOd/hvHdpQWvO/ZHStFHPvlDlQlsq883C2pBLe1uN1YskFREJkjVUudzOwZpMEGTuRPx0dO
X5yB5UyO0WXGv7tCkIsyJ9HmU+039VsUxDcFXYvAFdnFm6YaoDfVcOCzHFcBw3vRQGMPQ262oGr/
4f7rXxdRO36hN2yamE/x0IJ8FUGc+rQFzPdoC/QufobkwPdHcGtdtzVjtzTcXQhH8RJ2qjiYmXek
Ar6JwJ+Sk2TPcIFFOMZxt0Pqhkly4qs1BH0LV8q9fNmU+CsCQSBrlnjYy+GhAbet0MHIy9vWO9kf
bbKihswEzO7q4jCaZFhs4A1ULB2A0sUVTTJIKQnShhkwCDfjSOcLYS+ynh1BRJWAqgsNo+MPWUqw
LV6cHUV0w0oCbBFBmrAmcQJ1KBzp3U7DkuinvGG5OCDgBmS6rRLmDg4vp26W9/2jlM1ltDVwa/b8
4PuEtLwQA3YB6EMuRK6szP+/PD1NqMLqkC3C8c49U4arYXlQ0fgyHyQYomDLNPfz8NEWXOBsPNLf
IVEV/4ktgdgORmqcAouaxbDjGKIcEk8uVBwENQk7zUUsuY1I6RtWuKLpRnq8/Nd6ce9AWous5n1f
gHZwsx7cfXxtC4IvGXMkXxI0uuEoy+Pumt3n3T8ldXMvGpH3LYV0mLgQOcoGyKhFeDz0c/lTUdjV
GQLp4MMCm6/pJyinslgop3/wXQwJ0pHNO2qX/Rif8kBiyzT/RWZFNpWFG/9D3PY6nU63EkJeV1Sm
3sSPJVbg8O6Ty0+3GB/5KB8BsN/4IF8U/lvq273UIbAHzvhIPz7QKdo+4UYNSD96LrhS4EPIFblF
fLUfMiJoTeqsnYf8ebtToTDOwiK7ySOcvhl6kTc7sVdEllQQzwDMT26TWMTbiTUqEBGe7HE33wvJ
Q21irRmSxIrNBln9o7VRO1Va7FaModeyVX3+Ipv5QrUBROkz7/+DLd1Q9INjew614Pt3suPpS3OK
OrYS91FlTdUfpZUg6E1wUrEZHRcXkV4Wc4EKqgzOnzmCrmYnC/zou7H8n67IiWbSGYTrTF6WQa9Z
O1gnpuSbsekttVKAN5wdOiG7IAYXz0VA2TwXBYJimYrMBQ128qsY6B6YYA35KmbruGy0/ysyckBa
h9MplHpYZ0oKgJo8nwLWDW7JjrnLzbwmATB6tumXP+qOvuTZy8B816vz4WepcLS0HMgr63Co6ZFQ
CH4fD2gTOX9lQPxa2ocUybKeR2p6asPGsR+cB67+2H4AJhw8Cl5R8PytjtLCW2L4mzC22wXiHQLT
BzCOf+kckvZAKZ5yr+Vnp0z/IbujGFmWANN3qBrNIVEfLHSnxvSQShMUNUIUCH1Kym5ek1KSbo0z
Ldze0hg4F7FHtIQmcKtguNTsZBxrdzs6id2djWrRfcRggAMZUs93P3wz7HxBuI53a/7fO+8mw0BR
j5qWScZGtO1yzdb61+Qd9n+fOyMf54jNuncy1+EstNi6pmlRzyregwM6smnqswBOra66WLVDMTlZ
ghxZ88br2dvRnQQf99kDvjBJPjfj4zCi0WvNDGAu781Q5vcjydq37fjP+N/ouXl0n+E1/tl12QI4
YzLYMOmY0OMqK083iWkmbpeWgyQ4T7lNRjI7xmD3xfvibwDHrHujhEmSnmW5x4JIX8EXox2a6N3t
kRre5iVF0de+y6RjHj9vLkR/t2h2M7kMO/mm/dLv73fEamjGZeJlxYBgExdApz+fyHYXQa2BQAi6
E0yn+1ux86wSMRXGaFRkuVSqACsZDrzefOt4nvXZy+ZzAszIzPaXpHt6kybnoFy+Vm51pz8C595Z
5RCdoqo+6cRj13rjl2aPhbhvJEhaoCiXrBxDeAykjeGFimVsTboQ4y118Rsh9mN5i/oWTeJNhcpQ
kGLHGlOLf+m+qWDm1KZ/yTtBvL8JgGU7hkh7dQir0AiTYs8J6C7rZSYtAZHj/2KwUdS0/6gifxCV
Cg4b/m+hwTUPRZ66WO8c01HBPJt5FYRAYHVZasQxDM7NPQLJ84yuEQoP+lUIzUEmuSV8Wv3oyESu
LO05W2qcxoxicC25GfH+G7rvrTN2JZnvLaQ0McLYNu2jGh7RCwIu7vSx0IF/4wEGkgwFME/7A8/h
ytTPKgcliAxohWgT/Gy7cch3Eh6w+RxCAUsRc8KtQUr9Klw+BPxaAFCqs9EsMYj0OK5RGi5+0caK
ZDVW72NL5FJimauZXUwiyr0TUzMXb0gUMx8rLAFs0zVT37N7f5l427PU8okpZeWMKnPq2fX7V8w2
p+i0w/MWLffqE7lege5semjcsR6NJ9mXs2THtzpSiK8JnT+2xmWqhyNIjbLel5ZhSK9ZvILx+Gl6
KUuusqk8VX3JPNbmBhuaB7DCGupAx2doe08+uRiUBaTphKXqNKXrOLAa87NprRZhZ2hyteDQIeta
wM1V4mUfuG7Sq+uvJJuwtOM4epwOKKtfPXCyQKI2guMKFpp7sS8xKmmJA+th7AJbSRZcZdZaHiJM
Tq9vsFPH24ipjsRiMC8gMBFFCL/Bs7MAwlM7qfXSpXdpF1gihJ5hA455UBcUlw6pom2x3oE7b+5a
bGZIUhlwZqEtQpiN1/EaGjfCA2VcTaxCr283+BamtfD59MXuBggP+mYh/NIuVrtcl4HzyKQ8m27l
oj6hn0lzDB1IBvpQrr6kUAPz+7F9W0SiZq1khCek9KUhWX3jK+beBQbr2Mtx6WjaU33vUBynYCOR
0aDn9YHHLxhqPeviMpkO3gg7usW4623GBemGpBkD5GwvaIRS1d9XvxnKDVxdC3iBfjX2LYmF4LUm
3cvJS53bNO29Sjtfy+qng1XXgXVtGKBf5VWt9Rflk/5+gP66aid1sZYYKUfsj5mwVDxQzK3F1mh+
PxJwJ8wWXCfKueEk0VXA+z4omz4bqboKmfF3LoK5Pt+9ldmdxnObq9fzeG+L0aDbXwqwZVpEYoC+
EMsFYVUO43YKJdsiENZBMHfuyp+XX3ppnYzmInuisP9AceIKRIQ2Smu0U7xKk/8hWqjeMJPpxzox
prgqG1pVnNy6putdfXbKCi3XzDl7zLfm9pHa2q081+05mKW37YBP3AVRQVV95L4Ku6LusvCf3v/s
vkYaz9ZVaACYbKHM8vYxh8mDkuuq37BQXtP3VfM/Ms8pMLPm6+58MoefCRL8iKJoXz5OfPKNMIfY
mQN2VLPb/7MyaDcRFCekhQuCQrZ5uoFXwz81kBCvLsntbRjpUWXBM3OQ7AoJX+uW8l/8rNqhziA9
/fMowhg4ZJKxDCYfEALGugYMqWQWRuHMo9oilr5psSaZUpTAzQ4VhDNEeR8GwGoxG8oQR5I2z79r
4uV8ohYIQaOclAWZ/I2A51/qJGjaXoZb9ITDs9rBsX4P1xV3atsXMiwt4IAo75iEka8h5krdmOqq
rj/TBvsLnCUvuVcYGLIbe9p2OKp7ZtJoub8XvYTAB4MSjOClgEoORlKZNUJ154C/SJGWSGWAlpiH
cXxX16EU7k5WNTw4fsQUNwbWJbpMtxVCLS1xjz6iDhMEBwszwjsjjf95lUf5b8+5prlTREbXcf94
Zmgeltrqy7h0v6x/vhMrtri9cP3oD2tqM9igt8AOnUHq+7JOJ8x6YTyJl4ihWfYh6NYdoS+EqS+W
A931uS1qkq6IP4z0PisNoJZGShCOqPudPfklbN5gwiduk4BbirqUJT8c0l+UMqU+xK8bb9mWFpSY
pvivDryJgz88DwZVRKKq04HY0Euycag1jSR87n6rwRUod4+3SXDNANr+jFBhGqpbdB4+hSPkOr1q
RwI649p/iS54Z+0MyIkmydppQfiI3sQkUn8JrrP/kf7XyZsMEMCxAde/MnUMozd6rwh/3HKVxGIt
su+KyWC3gnORv1rSGawFyuT8yZ81aZKGtv05i7VfasXwIMoRl6AT80pwn2L35PEMAi3faINHBP+v
NV7UfDiGneLwt97lQKOPcCeerF1rLzA09dyWeuOgY+7MovpRDfuu4j6oJsD4YHUNJWNrluJ5G3SK
53+oeI0pwKf+tkfxKGXJ2A8DUBMnzsZ0m9yuK+ePej3EQ4iTeeAAxxWDoQRWIfXtyMoGi1hhfdjk
UsewrVMtII1fmlQjQp7+GDPVT7XJGRyNTeucLeDx/O6XfJ+fAO7MVolJ8//p/ixdnuaDs3g7Cktm
Bmll0TlRaal8vUX0OKeplKH0CZ8gDCtaHBSsIGGrcdgyv/U3sRmIHXQFdboP5nP2osDcQNL14KQQ
gw5l+mBdSbTUx5MXnQ5PFXbTu3AabbIJladlEKfVsGZcSpBT7slsiet8lguzbkOGGOrteLcqmIVh
HUXeSaYxYdW2U+sALCeB3vNVbg82d+i/jZVB1pj3igRVTHjWko8GnIRl6sRs536tXCu/UyVRB3tm
rf3UWVsoPfXgKQeqUWr/Gr1Uh1wDWIFsvTiFa2XG83ZRE8BR//c+Nb5/Y6Hts9nsRYjt9HyJj14N
NSYXBVSFMRJDY03wQJlEAMctB62MsMv09V84QV5oZg/rrPcji/Obs2+82Wi+kUBrjtm+UEQ109hC
M4bAyhlcMhYA+PnwAR9DWN3N5sK1ND5Hk+e224dlHfJjgd5mD88sV3NKpFT86CObxVjwHWsyj1+m
Cl7yYzTOdubx4Lo2IA6Lyf+gzHSesoYUlvLSEzAgfkRDyYlKkvId6ciSeGEi6oSoTrfxiBTDVJOO
5fdenBvTll55Eyf5YAbbbtru1IKdchsaLdrrkTPIx8qaKxwSs0IMvB7bfuzswhWsOYejU9dtqa8d
MKuqs3bSV6S5pYyqlyOujgXfqoWPlpJbmH/pUQ3GIfKco2lQSJFRzzY7mw0ro9MAoFHvkp0I0oyM
bQ/ZtEW2fIbtix/HneEUPNodX4VzPELQaV0Mv0i5WeRnEYKjwVxR0kgmMVVvH+zIdDywKHFoc0nn
JGN+AZY1RGDzI2uwyE01Am4HOSmu0i+8Y9w2XqsuTR5pMLf22YbBnUv7pCd3ygzR6AbOtOiMpq68
v7m3vID0opuObJNqjAsU6ml3MF5MxoQIV5msRKf+I8C8hDpB7oV/sAYOVrJTrVw8sYAMg647fWg+
A6o0j5GpB1RPHnNoo+f6OHpIeykIpIprT4Z3rk+L00fmXYIlB6aw5b49KE3/8laNFZxvNzz9LEI6
eTamh5FLZynV75ugFia1ERlzNBvufp6EI+iQMGfFBVO1j5LS0LnHCZuYe9e4MTGOAvShFdazm2Rd
2slACnB+FcMBeOiG9BpNuToZiizcjsq3EFKFqEqNCQNcE36glz3ZiY1HveaycfjOTTXJdORqPPuA
XP7KzDo5pVj8pFSIAZrqCk9sPlZIvwoJhzhMJP/H71t247wnNp15ZIAtr+Vc/rIwVFn6FvF3C7/R
flGMlmhuqRZINEz7bTOHvhuSTquMQehPd+m0wl2H7CNWtyB7A18xYqVUQLaZpUDF1PM5nzlML4EJ
GgUS59G3dZukPKcODXGC6B50l07Jxh6kYaiRwtfo5L6fiwnmPagFmeu4i5WCcQmdABi5nnFtlYI4
ffwmyv8NfcK2QIvrS19iqmmAoJHcho0MpZgzTA9KV+5ngwle3oGzIQSbxGCLttovWUKstmGI0spF
holiRQCyrA+N902sIpJh9/J4il0Op++IXOsSTc4gwqyVG4lU3wHhV9vKqOi/V7e/FaKjUPxOObkL
YGn9EXmqPZMf0Rj5gSApxqS53SLLf4wdYRCxCn491AeI+rudApKjHYXF0o0XSionIAnv5BnJVbe0
xAhn7ycYvxjLS3CiCW86A0m624FmzpXfoZ/G1osiw6pTLml+ZO9sVWG3ASamkfJ91lSWCjh+zIDS
LEdTyOi8PcszfkDoV8u5r2GjOqyRFEHHCEoFikJEkaUjoTdhvHbzcHrIn9fBV4ZTfz1FFaOO4nfT
fsTp29SrFSk+5oV0JJ1bobvUQPPhjxJGvOHY2uqMDCWiXmeH7otuhC2TBzUz1ywesq11tqPe9PsL
8eftBbCrivTdOvh/lQz+8FwjTr8U9d1+bp3OD/PldOyjKst56Nudwq952YE3PRDC5D0FO3b+sO6A
5tVKQL4E52Q4/XBTC9kRnSs8ntzTVwYyQAfbYwJ6Dms/Q5WMYPNKcrTNJkVYzmto8GgLsc0wH6A1
X1ObopoEYiUpXdulhX02oNMJPf2gddBboRm4IaGSckCM4laE+hdv0574xJWhxeLGy/s3VJn2sFaS
TeypWWhoBvJPtIHnb8ex3hSX5Vlod6Fe+XcP5FP+l72YQSingYJgDqhK8kLYcKLicUGEpRQt3uI4
tePP6pf65pt4hXRUzbNyWfkHYWK3rehqVV4PzmqH0Pe45SNGz6thgK1hUCfNear85EJZKX/B2QhH
Xs4jpT3ymdmfk+/OUTvn1lkf7TJxBrb9molhyYTCmvfDP16iyY6xhuTrva+T3p9cJAz6W0pSb2qT
q+3OuTXkTaKxcVrzxSu+ZIiFvI/uSvLLf2mFj2bJzTCQ36JcDtXVm6SjHYanic1M5H55EPg0191n
Cy0P3hf6E1cpnbYn4YIju4V0gqoKHpLm0zQH8hHgczoC7pXT1j7c7Zckz/rbNAb2f2jwPp6LRTWF
J7Tr446kudIbfJMLtuBsGxYuLoNbkf4HW804zK6kbPZKQcT9lSO20jzMMnsD+6TLtgZvwX8i67dv
aaQT4VljD5JTIjbH9da0P5YokAQ+togJjXGFYCu/715sOGDjCKLWXMCo4XdnlULhtri32nYzwxos
JfZFGyOV3iZFpiAGNc4skq2m/0+MjtQOeZBzAHYZL01MF+pgFrOQGIj3kUv+8IG5ms9UnWJg5lJ8
KszptdQmdUOYnUqSnmgD9HgMnFyGdqxMjlmFKvxhjJbu8K93wag48iHasEIBJtb6iNmag8xiaNs1
UgC6cy1eXhZr3EkO/tjDO1rHRJleJ2vRcfTFq4kyuqbJzg91v6jJ1c2Z5UgbqBq68xg9mTTD0qNw
jg2tUpoRxG5qX+S75JmiY47XtfOiGiYVP74FRFwa6IYaAqjI36Xte8qGQ1jRzgIzY9l7kzG2wBiT
4TlyjoT2fapsTLKqJGzPvAgO2GC0O50THzGGJKSm2EYamOy2+qI65/2bBfRTCI165uhVLTvSRmda
MAyh4iuaRMOyqDnnocDwluUd/T8r/UgNbxlT80LIlHHrlmcK+2cLtDXToq40Z/DNRjgFk49FA3CL
tT0kRToaZhtbTK0Rja41Ewp6DZ5rYx9T2eNGXOGdU8DsYg8AOt4QwsNz65CYN+W6J5eIt92ihB7o
RT9si0e+9sUBCDCIqhN09qTtCDqHJ5obM6ppdaUD72qylW4W22fYj4v3Ei/MuKAnBb+9ntYAYe68
ozldEL9Ns6OdOtGrV0fGbSEIBMFWzJF4K6RZZ0/LVCOl7f8uXME/XL2lFkHVcyYIp95BiTtcCaOm
H/ceUUP20kj861dSVDKRNGPf34D5dXPdZKhKkq8yZJLSw53wOoMU7LtDCxokgtm8C98mirSXn9gd
wzfXq/Z4vvSfDl5lahI6qy5phX0iuCB0pQ3JbjziHlDD8h8ZRna2rLaRnyZ2DYWKeOjQZsvUm78y
MuAcqZKsVtgMJiVnH0dHQMEcXvbLdmxO4m/wzMRa492e3F7earFcQFaXdTpbPFhXAnNJVxaCuhzs
+MFUNVlg77KwyrS1cjg36c5vYUkss+YADWh4m3R1/RgUzHvFp/2sMyVmzNutRaiu3jTv9nNUW/2F
Qic1Xxxc0/cWl+YoYpEL7SZXa4pGcZTLX1kPxmKK0VThF069xkyzHcKMFscu2YUgzz+fXQa9rPNA
KpTIWoJVV9RS0eKJzFn/Z9gFKeyAjGYmADl4mFHEET4RAm7D+BbS2vxpKz0+gYiGZd4bI1ecPDTW
L3/vUI/oh1OjWlySEqOTgn/bgdYwpnIrTM/cTE/iws6BNFJ4uULlKaBbEvM0B+kTHbZsojLZWLC1
HTyCmaNbLOYU5ofZ8+p4SYg390Xaz/G7sKP06lR245RNp3vv8WdnoYt3xOt/Sj0wKSj1cdlK7fGH
+2K0xauBLC61j+AjoL34GehvBzBu6lNbbb+Hc8MFTbBj3Z/ms8swcVN1wwFNw58FUL5YtBIoEyKI
H6FUNHaOUIxZiejlyvvYQE5LhyZUQbSLiRpSYVFB+xLCtBswoqOEVK27l8i2qchj2bptpvZJb9VC
2qiwU+l0D7ocXY+KQbrdk9dKNtyhx04DqzzeBIxRyHV5amUdmDzu9d+5WhQQKPUWLZbOcDMneqqA
ht7wVQWtrJ6S7jOKMvlCjrB3k+C9hl2oUNDKuVeWo04IqN2AjB/cCLRMw/fU2Cmgsl52ddw1dgNN
wtK6bANC1CZ1nonkEQIlyKvGt0KVrPry8wLjQlTTiHHNm7FXZGqkslcaKl6L6Ejk43o0NAwqUAXs
lahihc3ud+4ZZTY3YkEnYbNIQFMeeMKTfF1iPiVSWv3tQfsvyG/fE2CYVBYETknCj355Kf9n6MSN
+QuCTQKGuUEZGbmIK508WMKnm8IXPYRjD9vk/mFc2PLmL5bHtORrm9cm+48IwnafYt2VdNPRzgvl
Rzx/0e94N836CwyMbAwfTSoWWDKF5NOFpOvQo7NU0JKWXv/7fv1WygZPJssg1IXmFKJuziKk3TNk
VHvA8+gv35oUZmLmhOPGUY2Sw/ceYBSVlmrI+C3w6sixeU5OTExIuePnjtisQR5TQbnnJADFdcOK
cL92Ic7kvvl9vtNELPms70xvscz6bW9XD/m1GhUx7r/vds4AcEF0uz8gdpj4kJc2AeNet9iOuwks
n8Nur3yLdlDVvdp6GxmQ9adw96iMud1cS7JITMT4HlIo1jidTUC0cyPJbxpd4LLHTdQ8Qzp0P6Di
vLvfPUyqg/3Wpl0QCDwW1LM0wozqDSwobKU7e7+e0mohZkPvfnUk2mTenWvJIL8Ta7oGZVs9UUsT
+zeJRHcHfVG7J6fO6xWT/AH1EPUcLEBfEJTswtmTd9Q9sDTf4IWJbz75oxI5tbPdwJyU05OsOg+5
qItceeBiL+dnQUhr2nxn6cQTpObnd1pzwR8hP3wLaUaH2w/CB0u92JbCfulLvdlomVeVUkzZ5nIX
TquLL3PhUzrVNkIhZDWKyxmap5o6vxkm6B50ARUOoRC0nDB4U3mIQycF7pB9VDLDfmRk4isl6ON4
ECh0ZO9bwkl/N19TtJlSa6GE0BrIJaI/B75sLCgC5aVm/5TrniPKrBiNrDSnjghw1HIHygD3O0TP
JGdi6/x6Czlyuhk4ouelvLiMlInU1/m5aW1s6m/St/QhtGz4I6ZZLGnzH1Yd+F4yQmI9nRUFV2hY
f+cznmt84KBlRZoCCMq07yhcVGuSE6Fm0phEeCORJ6gh8UAKEwIho/nNgKx5EBm5lNAa/sua7PPd
8/Q+PjNbkKySvBSfIAriC9SWXT+yEYCbOdmVLGEANHS2LQtqyNbvDFPh5VxBt4xtpB4f2Q4Os+xT
FBL2KNtTbTS3ECdWI9FHnlD6HBg1rsfOVty2hIWfYtMjgH7P8oG3BXPUaezRekk+VCpjQK5r0QG/
s1RVdFGs7tCRViMr23VnGctgJUBvhhSuYM+guQVAa053/HzhuzeihsG9/QMbVNLWvGTb5YuwnNVQ
UeBy8Js/EPaoM67HAUCokCwraDcVnMrq3ddhHZYoysfKEBzh8qZmJ8gEyAeubNc8uYM7vRB2esUE
5Ls4s1Uw388O+xYb+3lDxydao51a6lJfy0TH8FkxHUUTc7TJWDVIjAcWzaQscsOr3vlSLLkApIOX
CVmFrj4Quuq1DHMb+W+TGPOjXelASS+lP8ujqbAqSFnDV1CKrP6VSiVvNObOAvdpMtX9YobntzIz
tHfYdoTpAGKw5xBLU+0hUC/Ny3usQEnF72tudK0cpmrEdJFxXQK71jk1j5iUnzvWyYre5JfaBBWt
zV/pkHsdUFugZpDLAaw5zoOmem1gMR+vu2uXY025TmVYmIw3tKDbs+N3OYgBcoQcjYaP1FUpFcMd
khKhVLlPyAjsj4nSTk9FQ2UMw5nX0/iSORH+SJIBdrT/a3tqMRqPQ624CRzCGlO+2E0zlGAoNYcj
wmYJiB7bhcZmNjt2tL85DBayWxmfaviEd/1uYDdZA84SaaOdPBYFertU3KaeOauDF2ycCqSBSmsq
3l64R11dJp6wyHYGFgGdfjeNBZwTaMnBPUFMCVxHGSLPyDE9TenIE0UpLGlXpHEWYGK3k+ITXbdg
04J5JpL6/MDcHIJiaFXC7eJenZDFyHgr/23fTIYV4zonx+7c69piJhN79WAAlaWpTlOVZdsaxy/L
4VYAcJbqjBoFrT+OZIFYXJ9nBY5maKS9FL7NyYFhgtwj4JwSXjQtLZFsfaGdiRMaicPStoBDjLIC
VuAVuYRqtX36gmc/vwNz1Q5IMTrFIUTnFuWSXp+MBnu2tooZzlk8fwMXpsglj5SGz5ZiX5xzhUta
f6d0CRQkh3yAm1vuBPPJIeDwV2wSkiC+lzbLFg1t0PyeZMVsBvtsA/EDGDSBbI9S8j/9ZbsZBmt8
z1V7iduZc38jeuFk+M+v9levDIjKyHbTOM1gR3fV4Sk0XS39+hqIVgQyHXlGy6a/LRFmTHBxV/Iw
vOjWcG27L0hT3TTq7uWCRt+Hrc0VzQ1ANS4CvUXD7NwLfF9iztUau73wKuKBWH6ZmgMPe5XEtGuP
YANNmDSA34VxV7W85a9T3WwYv8uvDYGRbPCJByVrlPXxdvAVgqUibDnrJYFOF1zMkeJ55eEBUAdm
fmtRr0pIXsHXBppJdifI1ysCyX2s78oTr3kce8PHzZPjr5WZoIvFDvHiQS7aBrY+OdXzadnr6NkG
1to6bQib/Gc1vL84b6RkbZahedbCiXjRxRm8Gb0ufvK9UHO18qrrzsx0R1u9QM+24F4iEtw2z+Rp
JttBD2HSB1cBdOSALhKme8v+DkjjvwsLsSV6coz78/+/0y1AbYTiT8WkoSaAfk1jN3p0NVF2nnAE
eMgOhZDctddG8VfyBtLXI2cRxW6rxnQst7HbrkNlgKUAyKnoeVE17yR373FXKh1hvW/qy/O2dfXH
CyQEtZ/+8BfLXtCqxdi3zrPwmUXm1Vh+s3RBmEHb9WqvBi5ED3i+e4A+vxc1HDNTO/xGZIOKXalb
11mjZLuXdmR5SK4Gms1dq1xj0wPaJXX3ubYM22xFNjnC/zffwHIgiW9pUau9i9Z1ORs+B/iYF4yX
SKeGUC6E6RcyyGqIGDBE3HuGcZPZNkUEAeYa6kyE02OyI924Dg5MeNSuOzIvH1VVIOmtCxkG9QIU
3RQSiQNkiovVks/21qzwgl5/aXOkPPA+XfHP3GrumXI1octrEDDqyvtz91y7ScC/9OE12luwmGRF
AGRix84XLEw+wL5QQzo57ipYNx0oH+BPrhoyJs+op26aKgTfevNMpq/G6inSYLY6UFeZlcWkqoDl
qLEaN58AeEOcBbHkpy2leeeQsKMwqUFCvPtuL9eusmwZU5PONtaE+lSWtzh8Yl/Z17HeZG75wBQe
oeiw69SwUnG/zUn53rqaAhRm3WDYtoAN9dksA5j8Oc6cZPrgsMLQi2s5JFF+xFtxxhEc5Vadstwv
BR5mORwxT3wpvbaRk5oR5tPxl+CDoYodZZQaywTyLehELDGXFH0pCOr/aWtcE7RCz6gbuow3JgOG
TlL3gE3GAW0CUoLzHM/n0aM5xnphOpkquB6/EjKKZiwKeRx2kuZQqOnrRjVhZGxt7DHpyYfb6BiC
Ny+MWKMaHL27RfACOVStienMBNPEoTwUWTdt+2wY+msSxDMMzKbPLN0vFN2QZdlBTrfDIG+nurHZ
iWGVmq9U7AZKIhMwfO36A/cPq/pLNCyDWlKlheV1YFN3ijv9n9DBSYqHXHrmJb5gkoIYv5Xgx5rY
NtdF6H6GN5Rw2V9tgsezoa/7ROILbxaocYJPdsZTaxQunFr6VWDTH1ftU8OdwL+e7IoAIpL1dmBN
sikZwZze91S2Xdcp+EKx+U7BexeBbVjTq6R3Wj4w4/Ts0pKyLn/8vYV9Oso4eWLCN0M5D154ArpB
70naSxhTKEb1gDEN2EHnkFt5bKQQ2fqc/ZY+ZZL42HPf19YdRSpOiLStkmD7Ju7u5F3ciHChpJjp
hH+BpjXXwD2xfOJgQ1HBk8XYoRGlNWH3DfymIvlBC+xBDFPWb1AXtlMPDjeph6uke39O+3VrQzh2
Y1vLU61Q7mhYB4RL3EpOfVUsMsniXdotMapRupezib/7cqyCS13yOZTPauKQfDcEQOWK5JstVKmY
ONwo6PQhqzxu4+j7Tj+rB/v6PWmFgogoN4qdP1gN2+KvcktxKJa065o/I15mQYDaPeL55x3AcrBV
vhZN33ckn17aGVsKH9ho8DjcKpmYnEqpttgAP+gm9cRg3ZTDUt1z3ntX0diJTne3wBX8qjHf97kF
so+5ynrwG5k9Dctb6EjV3AlOE08Av7j6BW5wKH3c6Ob73z9SqIzkU2heXKQyE84/xwt2VLDfaMy9
RDFdAUvrofU0x8gfXGztJQGAebP8v94Plvr28NnCE3qnPcKDWAYKsNaECEHT5xdlphRo54CpO2hs
ha0rit1ndoZEqOX+1GL2rE72aYGfMVHrlpOE6OjEwsb4K9TICt7fGfP1nYFYVz9LnzSqmVEknWOd
xSjGusfw4wPnUk8Sy6+xK09nAttSZZQGlvj4/SmPdWxCKUo4Hhs9RgLj2xLAgXRv9z8fxyDB2xnW
0HLCNok+6gjx7ieX/OsHysbI6d2ftERBxI2tns8HuB40YkTFLf9ILpkk5ch3Hsc8nECNknKTvqwM
0oefZ/11cguCV7H6tuc7GpQvh8gVgO+v5T4kCtbEBlWevIlKOSWSDH48S8Ra+u1gZIHIrgotIsSz
Y/OtCQ4Hg51AqIJ7QEShbGXoKafuo7jkv2FLmfYhlQYLyrBukyhug6ZPG2cipLp8bcsmY2/dd92k
G6p9WImlRh+5Vg8H5L5zoVSK58tnBkfewTUKLX/8yTRIVcf1G25PqNCTOXnFSrjMajgQNRWPY4vP
sMjnZmgfUBV/Ryp6D+LQI0TOpPOmrpOOnS+6BD4cmoozlp6jDVfebvDWgUd9m2xFAD0ISsPAAhvP
QLYOcaRQsrnq1UXuDEgzvOvZIQ54MepcSeuw3JpmFDHT9GkSLJ+ozi6chpfZB9MBgWQT5SIk/Fk6
sDrwlNsaVFi4wdx2WkdQ4LU1qV0fJfR7a/OCXaq5r5QqB+d3gJJ/33x47rkYtSh3g55Y52i2pbuI
rtehXpSdnIfBbSLgWTq8D9RdVSKlE+NiX9pwWj95+fhwJD7+azemnBlViT59/HkKhWldygz3XxVG
LCvSMfVqw9rtCQU1IiRAeHceWvMzCrM8HJaEk1tif6t33LVQ7A1u7W4kg4PvZt30zANuIHR46pH5
G1lQmKtuq/2VDyGuQAU2YjP9E6xFv4ggjLz/bE1JGR2ZAktyRw5y+t5BR0MpOA5H84XF1CPP9fvA
lUARyIOGTf95SqCY2UE3cNnTnc12UctticRsZ+6Ps42BoCywyY8fnMpNyT5JB4esoLzAc5fWObFs
5zpE/bJeI66dQFKrwri+gIiDsd9l6FoqILnK1bxH68DIMYsF5gTkm+ghWnRZ8FC1ZG66wkPfDJi+
SdGYCsmcyldlfC7DUPyABSRCJ8aBdvJHPVhiyo3OrP+7rd9vi3xfHMiKmv5zgSfBzvCQKqgTI+US
Hoa6UW/+qKRtbxYO8OYIT6y8t/MmfwMGMduGObVRQ07e2ZoPud4zPm1vokU9BZNhaZ6qGqqy838y
9NtfuTSmmtUKSNMvusQo9aLkQ3eP8ZTFkAfEoGa8Q0KQkSmYMu7uavds8sH3zLZer9nIotpISUat
RPy8HgN+FEdUcf36HOM6YdBDRf8mpDoKTvEjnLxKZCRn9JiAi+OC7wMoqJ7GyxlNimY98JJ8XVSa
rYY3OowyrLLLrUrmAMV1A22bJZfOes3JD/oGK4BYRlaSF1hzPRAFR79CAXBhIZCkLM5EhkhEA33a
FzCcwVrrmkx4gWaiCu+9jdvJ5JZ9R5a32jn4omAy5X1WFETEXjRbLu3Qn3fzvo6ruz7mL7ToACgm
6QigWEgM74xNAqkzHw9BwsS8kl/HdIkA9UkGogrbTMnZYEuULwNcLgMpTjwymhQtOIgVyIueMUob
dQxaXcvAF4mClmQ8jXd9vt1Kg6sfWSQEXTHrhkkMIyye934tqQYvaWGbOjcIt9IBoWNRRNeXG+9e
SqaXWEQGg6aV5JT5XQAvsNESDJ/hzEZF40hxgCpccuJpJm4O4XeBPmdpr6bY0TEnzr/6ftW+yidp
/CJlx7SahyTFXNaW6AC4PwTyGUX2JErPdFBA0VAUXXMtZhrkp04lwFFpocTC5/EtUw0jY/6M42fX
5JgcsavtjBQUdyB8Yzrsy1+Gdy7YAanAy/z1vBPkKgzJpaoMjIPrN12uJ1t4nTBMIrs/drBFjFvN
9s4qlyvhBPeGaAmVimEYPrYC0IGz5OkvKBR8JPsyQ47KLWGv945aMlmpU4IOtP06n4U8cF++FosS
4GquyJT+dOPx60orxxh7DpAzXBMRjmqLWc2nPbNOpeiqZXdHqUUa1ztm9rmAU384uc1bI+NNGymE
ZwH+RYD6k6H8NsX/9f3zf6kJzfjllT7rwHtCq8mHtV0oPoFQmUD/EriJryLHUtMynjBNxKU0A6tr
ZAysfxBtL0CH7Qu9qLzqkAC25O27okVkztBLCTuRl7uwL6pN4dX3C9/umV1HmXJy3eEbb5uOH6SZ
GQlKzulQxZ/Lq4mUlTNiHiDkZlZKo2NYHcoXSR/5LijusxySbtn0zJv/tdAe2ALxJ4x41Jhcbw2u
YkbK//1MQP7KcbKi9wSVutaxq8ny8Oqj4tZ4BGgNTV3lpkNQw76FoPac0RasHh5Zvg+xvV4hGZN/
0qTRkIDIdAgmKATbZ4UZAmE7dTgpXy4NzBbU9Z497l0dRjz0hG3bUOPTh2Q8Y+iX9wkzM5O5sz1P
V9sAnOXc1TxNIB/EAuL4i5aAI6KDitkTzcDQK2b8oNLqH59kG8YzKRdZ2yagXlfLmKuRcza6ky7w
Z3Hpbw/XMTzM27IScMN4Q5yY91yhWrCLmu4wTajHZZcQshEglfO61gAWDZftjZleFZMfU4lFjMbc
3blngqZ5IVYCCs2gDiTd7owcrvyyIcGuc71X1J6bUj6ZCHRCSke8F+3YuqNXkU4FP4wt5nKymtze
JE3Gx/vBx9wse+s1qerWfPD+EhMYwHGPVlHBQedIZwlbdbZtRqZ62G4ssDif3Cgy0r+JxQPH1pL+
ePcVg8aMJaPuJpTHgX3RHpV2tHlHtXqST434r2vdHU2RLt+Lewr+GUACyPAshs1LXl7hENMRANko
r4fdPFoFPVstCQOtPuhXiZGfplkKVfpNAtixlFrRtuuqAOwdpLM6LcOftegdeYjiFPJ1BWpolw25
HzWmNe7nFIezlHn8lSXJbzak7dlk1USJBefCIYAI5e9t8LBD7+0mYh2fT6dRS0l8gDQ+pNWdwicw
ZPMFJNpgxTEe9DStuyZ+nTEFg+gMzxKGOgqTp5OZ5BxFFhR34sQj4IkpiX+8wbNb36c5YgrSWiRi
ulCk2qzhDF5pTZ15kiuucQLsnnfD9U6Wv9xTyPNTBbppeM60QB5ajoMlqbqUSJatTcpg7b9HOxd7
zMU/RfbYMFXN9Tss4O3q1Z1y5G2SLHH5VAHAK9bQZlGAhZxtKV8g0hALuxrFtFgK6SCVgpuuTaLK
yjHqaitW1PZbZCY20DG7TbDXoQYKRGtFaCeRyX1SU8GwZ5nSj/eVO7APvwfIXRbz/SuzFCAYs+wN
un6KbURu7IGu0amO5LFJ42v/SVUNACnpWqdDsMa5cyAgQLkL37+FXgbH/s3z6P4AMbqzf0UE3ONF
6iwrfKmpsQGX9ApEvDaxvdS6KoJ1xUCtMefeX/4TKt7xLPWVO7D28wb9xe3OytFG9sxX1kU4BYP7
X1CbaFBOaJTy1rH8VkmbteXyktRoeI17UjF1g5ShUDcvh87k1xvww7pQJuixuYhujkI9Pl1GmQyY
GbmJYfBa5g9a811tlNMuYE0LuIIEUyQRGXzBfCDce9GzHW+iUz8TDT19DYmMDC8nNpPSKkDtle7v
AukeFeOV4wAJsdjnNdsMjtIIUOEMuotEC9In3xTN/1nlQW4JUAldLgjLCDbrksgkMdjVF3Fp13Bx
dfjwobPc4TTyF58sCOjgcu30plkXkdPZn4Vg0F+7WhfI+JzuKi4p+XH9VCGg7WX9wNCnnAwR1dKu
TxlMG2R4O6UJQXArq95bPm6HYmRE6Mc6/780qY1i/Vv+CSEjM6EzjZdBIKgtKi0wBoBoY/N5mtsg
MnoDjWkz+5IsAtYWWerfEMuE99q6ipLlNg6XKs68F0DjqEX2OXnzNsREiHFZZJmNCc/qLNeaD8m5
p3b3nBJAhPVILSKKzFqBNOrYyLT1gzQv33JgoVW+vmvrOrU/k3zE+23ak0lWbBvoig1jvHa4yHBi
fXA2OoV+EGHvvBdc2Ge5XSxKDFza/y3KZk2vZ4I3QLwe+HD49drtuULg+at8pd9HdV6K5buZX7Ed
ap9wajqKgwNhae3eHcUko7NMPrHZEgD5us+0C3Cnde50qVQMOeJH2TT7KQ3gM9FBLblQzrOTJOdD
wca4yHdsalqDQ1rEPc0PMoyGZ5RfTpbQEEZWVqyow0dL5mC2mXrXo4s5w5Lg+9rC8Yahw4l8Rbmq
VCwY4mU1tlWXYxarfTPPghglnC+T6V22AXXAmX451ueAvuENuUEjTkM6f3gccOseBHB/gd8jlTqS
UQztwCgIDbHRX+2PnVU+NOBl262dQplTn/PxK1xGXrcCYTXFaP0FKOuJ5BjBFglTZmLIM/zaloVV
LpL7Yic8z0QwiYNQlnFucWwt1kRtMG+aWdkIVf/SzHSTde7DchCLo/jbOPPdIGn00iFlzXfksu/r
OiiDwGfOmmbHgqWR44vFLPCEuzG0z3g9BxoXjk1XZnwI3+PlUQ/B6SqHH1TRQttXnhXvY5VKaX8G
LcxrpuszY6wVkSJz8c8mx+R5LK29kMfLkzuDKzObld2WdjVAJyAJy1N8rxf/08Cc6oD6YAfnD+wo
//YjkyzGaFXkUBzj/ogoR1QXcON+662r8L6AILSKtohFfgjtTKcVIhVce9gJS7Vs6l368gvW3gCR
r5Ha5KibTfBxptGLYY4F30nYO49s73fOo3nlCtMpgv9kcn1X6vXA1bnsVgyTZw6Pnh9PAFS8G29j
UKD2WYjjhOViUNSj+fHeTQ5u6SV1EOg58QPD2IOirS+GxVMkgED01RC4T7Uqwx0YisbJqf425pi+
bbVbf/aQUJuQuNaMqdegtDOjAFskDeAz+G6JXcym9UOoY15sFfDB/51aX4eZUcWQbrZuG3CEcsRE
SygwuFEzpiChCh41oLI/sNi/l0fhDzUAT/MxbWSgJ3FEz44xDn0F1qU3lEl3Fac++Nv1Om/H8pPc
RBzWd7cSEui+vm/MMOQ9ZhnND9DgrpBz1iBJF+eHfEEcqK/d1KENdjF+tGxCuRBCZDq1CY0OWQVq
3sJsP1IWqE4/EGaG0/eX1fhcE4Rc0P0mOT6lD0vN9KSUsePwqEr6LgEju99PxBPt63prgjTYqiuD
t6ksngs8lXTxLGXU1Bd2ABBNmCcW+rhFgRhmlfmQVpnTA6QrQXszK30Qn0WI7BI8UIuamGMHX4QZ
5VE3qgupEz9Zucsej1OeUaSRltn/BJRQP+E+VHCVDgBLYnW55jqbv5v7BMplk0DFzbDutD66OCnc
jaSJ6nC8Dcx5uoxFIBznvsLtcGzbj/JURoBZj7kOhIIQCFrsXqdbTw/ZYu3N5CLxjhD2mE3Lx7nk
6NG+OJDRbne3H6qyFKTSiybN/i+XGY9zUtv5gJZzDQ5wJPmly/7dMD3OELQzcfkIKOB9IcZ345v3
Xvv36s390FhMJ4GzPjIb1arVuZbUTWM46HynJAIpUkmXLtpWC2uW581zGiNsBL0v7CIRkFTzOT+Q
VANhigfSC5zYI/5cYzDIUFCc7HMc3W4yZf7X43q5bA6HcoriI44lKtYlVTq4f4oK+ZHPj2V6+vbd
kqXKvyUPL2MkEnhD3IzWrUJqDhtQXg+OvH+2Z0paw//T10mSl6+Jqd3jl/Mku5mZXAMWUWIDM8A+
/7sq1935OT3/Szg0G4Y12+ga5BhC9r054ijjudxpU8ro0a+mmp8VoNq+4xDdIJlO7JxCmzOus7Ki
RY5jDmQ8KcFiXXuOyN1eAR9G8J4Peuubj8mm+/RyKQ0JPbdcdH+77u2pj6TGQfFIbKfGmzJudlfj
TdHXK96bwMO3/HbbUVN2BqSOVlXR86KEGOqC0FrO4buXc0g2aLW12CmmuHwwNnjLLwxFzOWeWSl+
JkqKCdB0dxycZB6Kk/y+woysymgSJ8g2PG3CaSOWXw70QqpSmS5xqtfQeQ4oGNF4FCGKZbDzzTbU
jIWxv9RJqPU5/HZMBSCfTwoVxtH/rdR5CJ62cWNRdgFERq7/HZMws0Fq4t8ACs5GZp3Rr0We26/e
9/Vqz2pfbZs6QmSQgOJFdNw0FlRyd9+lVIj4/ROltLWxrQUp8NhygcB7L5wBOKKTpKgd+umowdSP
U8+msPMhpTvau06VqV1oRjkrDPQy086KYuKMmy/WjUwrhQLEHuzUJ4oQOUDBuSLHpGzYHK1lC0Gd
BmrolaO0aAbtx43nxt5M3SS20m0evkdhAxj6PrQIo9/S+dqP0ADvKW1uapEfs7CT/Bi4ZrACOgJu
F4wCw3sL2XfRegzeryu/VT1PbwIOZP7ZEgy9nBP7mSGi+7b6nRtO0RRycw72jNrk9kaRNYkXJaSH
DniSyljlhRvFaJVeh9QWfIKz9OpZIgRam+H9HDk5xdxUYGQE3k2LwfU3z2RwZws8Kq0M5CpDFoka
f4OESjvK7GYZYlN0LgcJ4WvTIvU8UQPD3nvwyCVQgK/MLjsi8hKRi45T00RB+4hc87XC2/XROrtW
9UHweoHQeALnota+Qh+u5eZ/qjxa19Lp+ctL4YistrY1PwfOmzPRjvU3KFoYfOncgCw9iegOW15Z
M4nmoPxkpZyb0+Z8WchlTvrAlODQQ+mxDggrBqUrjtMw5RBAPkq0zZ0e/8nDzSLjT4hmDCFnRuhi
IYyKbVjYXQDIr4/EDhcAxlovXwj+yRC+ezuMV5vvYTK6MbFpCMxin9M1Csa+j+EoQQ3FqJ+w6cVI
07jZ8jIoJ/sSXywagCryz63vdyBTu+VXTpTu3M6i2zkGia3gH05+jv6Zryjz0We2hKmaZZCM0eK6
pPG0jOhgDEWgfJl/7uOYFYEm817LDcwf23ajq6ajqvYGhKAWLjkNBq9low8DT/cyKcuYKnPBv//g
Oju8zlXODMxAxf4DI0tO8RGo8exSXimgx3VLZ/v1H9Gtj5+1J6yehb5XRcsEW6ZL1O6pe5HVv8g5
kePUte0Izvn23wDmALJlMIXdRR/iqwHQZxP7Kn+TacIkvLOAqReSnZvm8ZGRGNO0CC0N8z8E3X2t
C0qZ3VQ/iOVF7HMIo8W3yCzD8uHgU36w1SL2hLv8hD7l+qv1NWPoUPSPNGxlf1G1PYk+MSCA87dq
NbjMVHJhne1BPKtoVZ2GZ2ikwm08eCNw2YgtWhCIVzH7IWYNZ5IOalK7ZMllaLuelvb8btYJTeGn
TigzGvkzwHHOQhc4uS5bQz2ovQYWQWOEmUjETUkiYFD9v49BZfx/piVEvG+1vNrfwlNmM+VU/LXn
bXdAUe151SfT/OeyUfZ1ZwgtmIiypoLmmVobONPe/cTp+1aTH3GnWGuRqwH/K1yn1+9yE4ONexfn
5vdoyoF2S8/0dAf0njbJDpNesmQsxkmn2HTqujfdvdZtM0gBG168oD2GyZVGDczq+qWNeHDeNltp
BrbTxvAJ5dBl90vfjZIunQPkTkzIhrvdI3JbGylbV+f1TjXwRYLEjk+oEnqSDkbz2nrFjwreL25o
GbxxkZyk+28Qj2q9ykNv826tArwcI+e86ZryWV5V28D4WLdg2qgciRbA6gcga1NCsU1+EVGiNu9e
5XDgfLTf/NKNVoKARVokkeWnP0DBFH6GqaFXaro8CmbZLvPKVwDBMg1KsQLvue2efyDtOvvOKXdO
XIgsyi0GDJhfz+eAsVP8d/AhuOPpu//6IZJBlAFTTHnJqKJHkKFrH6hEmVJNfZjIrMv95E8AB3bK
oWNUMZZ0WA7Ftg5B8jwfQxmgWQuOBA5O92mL2rp0Ld298LumDKYGFmCg3mIO24AGcoezXUMU5L+K
7g3ZBXx6QLuscRvOPaJKxKKECdIV14Dr1vYCc9AwDfYCen9O+3HleboCrjftmgAWyyegJd50HGKU
swNQDObRg2UpxgSzsuBditTMNUmCjfUHdHt/71SJJH2VWNAVPOMY+cTqGyx7Pw31npEo2XnF7pxP
Zetqgp1CzsZqUZ5jHU/LgUMRYPtniZrbSmg7u2yTyu/hDXV9o6QVKFLeQoHBvgy/qtYn0o04knbQ
hnOlt3tLvBh513Z3WO4RhBqEqzp5LjbVFiaL7ttVMzCte3Xd++vQKgMS6CG7YG0UIxyO7dPTVcHP
INYMu55Qpa/BgplAo9PiBLo9EPaJBNexQ6XUbMRuQv0ufifiGzsaxtGZJ0swj1Ba10+wEnaQc/z1
Io+LGgUgz36bQeQ2zGyg8ncY1+Mn+BMwvKC6YyW5z9vHVZd6HmfvEi6vOOpljHG9smvOE4Bex2DJ
qaIPI65ffmMAFtWMKuw2q7QwKqP7QQ9rIdDhXPk+i00LEHmPvxkIcTCC3CczbjDLDHylEWO9TMVL
SQf4EdB6AsDhiRuZVvft+yKK0g9mINMCme0Z/29cs9pyXrQuzItDd2GsU3/oNk4mbhcJOvcsuC52
6cGv868SJ3/VNHtOt6mqOyEV3g8AGqvsrK4wBnwOMwW4JEutVBj6iKX8qtRrfw9niJujUcOQa39m
i4RVBMbJASD3S132grF0rp4vMivL8VGSMO9LbB3P9oyYqHEp/w45zDB0zNAiIk6QkQEiJgCRC7GU
ZZ2/YwMZzX3w1zGWIybNYWG9apQIrAeEv0An88V+n7m4KE0QvAZAEXUBgXmZ1igfyoLcuMi/QjqI
871NQlDcnsWNVwF3daBz48P+3sEm0npvOWxbEC8SrZSOHzyL5UlUZtJFzGumEdKW2AMpTs8jokmj
BwHvLZufReAKwUXFEM144JyufF+xxbTwD96bdXVNXNDkDk17VgDJssHBZAfhb/N110rteSvJEUyR
FdZVQVJHuG9yUiCB4TqyhDahgXuDwy0PIXDp+eWuKEc4B1ob++DcQB2YbvQyptVj308/BBcwl9e1
8lK2FTt6aAYkITcNtitkHVc2xguXHqJVFz5nf4wk75n7p9JtaWKpcYcD7QFUcRFX0g6bYB9U8Gj/
UIBcd8BPWca+WESyFpPy4gLe1wF2M7QuP9qUK1UBllTM/WqeyWAZJEJHFVFISYXNRN4gQG0aIeTM
QmEnp7hcmr94TmzjcdW/ZY5K02DsrKbJEd0dAJKF/qzxAXxsCXzFSKEsSlNnQ21sDEapUSUpS1AQ
dz4CJDa/dmC5cABSFii3mDzjjxmRl9OUKUzKbjDCwpygtUsFQhQDfV3BA0ZRp2p9vE5KjbyQckNT
NUKOeh7ygR5recFqF23ZZoXmOfrgHq40wwk26Ta/5I9KKXRdL2KMBORA4vX86bki/M4Ib4ueIIh2
tOD9cNC0jEDB3bMtAQQgpcPoRtG3DfnYhpB4syZwUgi/N+jN4VbBtJa2zLnzMbU+pgAiuxq7Wz3W
Ozkemn5IdadKcP0JEjEwVekPKITJpDQSvfcEoMjKLaVr+6se/0aha+1SxQszLXpgvbsxkukUfRGd
ZuBNNimBxtj3sw8baZv4dJQqJpM5pFAfkWtG1LPGaIptxPBjaWdVunxrzWOVpIoYn6SIUgE8Tabr
cGLu+PsUFO8djlIZDdFR65qzvKyoNl/MY6nSA5ZY0Cy6OXxZf5gUZb5+s7DtOfA+Q32cea3LcEAV
7kR17uEYoyFYE505oqNtwQ+bA+yBudCFASE4WU1PDuxtbbMS4TGfbniNC1EBNWcc151kWRj5MPSS
PBmJe6SwagDJmfTgHbe6QcKD7r5Z0gFsW1Mv9YHid+v9bP+wcheoTdNeiVkD5lg1mFOu/YeSqbtk
z0ycd/ekhGXP4fncj7Q3Q5QNBnBTBMNhbxDLlL6nFpUJ1k87KX9w26EhDjcUEnfksvpK8AuXOs4L
2Cd8EaxHqhF3od+V2QdXvdAeLB9B4W5cR1vaEleVhe7wUuhYsTuuSYfkEbaY/OVdQVTWcu52Skhm
axXqYkPKk0D/OAbm8oQL7JEGXV91f0tgYqjGWKcS5M7gQkiFXzwvOu+pPjydZKTFu/hjpOLLrlKH
rpeuQZfLJzwA/cenEV3vN/zu8KWizZkdntu2dJDomIERLDSThPFLUyrdzkCmdMZYTl/0RBvWDgIz
Iw8/cK4r3hZsjcKg6k4s4XzdTn6z8KgY+JF+Rmd0Dj0jLxycgVXjXEXwKgxQf6/c/ipNlTIzdCAC
4bwl7Fpb6lMFoCi3FZ+FPeFJOI2m9LHbyXiwIi5jI+a48QI/PjdQjpvzJy+RK0GAYtTXfPUKMJKI
mXKM9X+oe33ntwP2ujvNagme6Xm26HPTbfozVRTaSEiB45f8pmE4kuNYxtgy+aAyVucEWfqRgZWV
ol//UWmvOTX+r75KPK9n1JgWydP4Ma+eR0Xi5Ga4wqBOEU6f+HYoN+z9UZQT/aueL0T1/6EhwuXA
b7jMrXS9UQXwQFtzYpwufv5qUu1iqxKyQ0WM2sgs5NrldFHj+FpKldncY4G8zaC653+nfux8iBWM
QO4xdzksC8u0bDwWfAWwJTueBogeoSaw7NkT2L5m32TyFNQ962isfIH9wVl5txYc7htOI+mEr502
ODer2SoAICkGA7YiPuTSC+emDFGr4uCUH1Y5m0U1unH4D1l7slV+EkhAWpdzIkKuxrBvJEDL5Lcu
M45D/xVaGX4EyenLf5dvPuE0OoxnEI5OtWclEYcoiybhk/eRIhzVs60c8T7c0K3x7f9YhqiK7f3F
zfJyqQA8YB/wcC+/IJkyofz97r40HWWW37HnDOWW2DT1G+9rFSocg/F44ENv1OM1z7wyNCVl2jrq
1FGot1MGLT0OCnJw4iDqNzBESCdBHo44/AwdW6khdk5L5/qF1FiD5rzes1y1axBJ1N2HfHUOtiiS
0DUiK+a38HxPFrQLeTO4aG2/Jbbj1mxNjvwqTeE4Ot9QVkBSbntwd/cd5tNdr6oABdYgCTKF9nnD
t38PRzD9gm6nrOngVm5ZwVxtR+oyBoGaMDbAEHmu+KI7PAw3TvazODK+1r2HpxUCeKVJtPSDpgbb
4kQ2msvsiy/XYV95tBYmCgrKv+kYkqc8Sq62voO2Fd05YnTg4IN/vfSNmWGKfLkpwKpRt7v6Am3l
e76oZSYlDXu6tzbh7QZt6wmUtYP+JfEI6NH43t4UCqAJU4q9rQDIPmUXfLWVYff2XobYhAfeXR36
lxSgZ59l5y7dUoIRTi1n+dBKgvODPtKn2QZKR1en+PA8u7xFBqc3mpIaK4q8uFzscjhi/7nUWIbS
VcepZB09/eg4OXiQjkE2rqnxYlKC9OfIGJ/LSy0EkxuE+bddlLhn9NCAC+o+llGc+ksSXTXbavOD
O0CW7ko4yRkjeUdaxsWjFemNzBEnyJM+qa2mrZ2L7lbiS3uhUnwAChPVukrSuCrKitfdf23vTBiS
2iKm8vnLdEsGyedUDOFJX95az/2OlU8UUPbvj4cBD67IiefHdQgRALMnVsNGUD02VagXKvVkKThQ
RnrvlTwPOTn20ChKT5JVndDEUiWnAklcUT2uDc8kVNdxwNcVb4Zofmlhh9WwCvB+7cJ6gDOudl3C
PBytaI0wUBMq7f3Oza6QLqiccQEWKDEIHCD/5ywNSx9TISkXlcENXsWfEN1zQ3nAp7pkJwE+FSmN
pFOjkVkCZSE493UfZHulijZ+7TraWgkvg325rso3ocOrZ50KXoHKaf9J/Xa9jr4AtbphhBPIYNPV
Wq/x3UeIKuIsP1hrypX/wf+431dg8SdNcAl21ebByvucOuyLahQ73yldbrItlyMnv3ntGY8By9mx
zhlzZHVDcREIJKrKL8H6S5MJr3FlCqd5BFK9KTa1dgRx9FEzadRtxrcfK2AiKXF953tGj4QylP0y
7EDSn1F3XU8rUtD+2+5k29aVfCx1pB0lLXcRvRLGjeNEaFXv1WPXnmTN/w7ejxZa+z26cIETK6x/
UqOrDyrDQkdYWV+J5KxbCtcezRnLBPa+L5wWuVz26k8lTeF2SySYJkzGukDD4LaaYhCXxACtKKvn
C/3KUr9wHsyfl2SRVMfXz/bJEqfzf3uZ83PEOKzz3d0rS31gLz51JaguZz9SlmgR6f41+dCAeKCV
HQsu2Vt+Texpk+gBsaIJV9qsNKRzdgqieBUS4L/Fw3AI9mC01/Avi3+NTrpun/WE+a8/hD9+fOfb
A38zlMJ9+mpFpc5PfMHyp24V5SeWq3P1qmmMNpWlioTtboO0+P+KfkN3bfF6Vyw39ZNvnsCjqq6O
C73wqcK8QVwsIYA1c0S6uWfxnV80kuHV0slFCw3zGkMeulRHK+6fxC6A5Cqk05QDtLLJxlVYTx2O
KXuqJ5mL7z+ZwCUj7EGoOZmpe3K15AezMWk8CPQP3lPyhurWif0Zqdp5LXVLdA0x5pe8/K557T8U
fCk9CflF5rGjlF9YHKlJdFYhBtwI6gpJt1+g05AkBCmDd0IKwBxLa5JGrOsjyJpJ6qv5oagHUyEw
CnEoZKpEOh7QLGL5oS3X5lnHKTCy2tR2Jc8EFvGY9+tycSJ8aWMuGCQDDSF1VsujVFcB6e04e+ak
lwJ7A388bnZn6Y5iFZRJy9xxP3PPCzpyrduCEZzonnxfpKk6W00j8WQ7FTVLapbEk7g/6ob8gNld
TuFgpZhVv5g5DJxotyw3bo84l+Z8ZTW2VoxE+SCyIhSVPp+3DivX4W3u3F4oJuLhUE3teqEvg/hW
4SAYBiER5XJX9hEi4lEfAOqnn1PRpKEYRw6q2zi4gVycUn/7VKvkUwhL37207wrLWjs7TcjLEWA8
iQ1w2pj/QVo5qL41KgCK7eBtsxwNQex29V1skzrKoY55aX5qFFd4JjWWaIYcqW/Nh23p4RHGQJWg
V2G9o9cGUDH6YTXASQst6vdHMPmHc2Q5T0IVryvnTvLhCcBv9wsEaECoVRzNMr/vaP+uCbvEFP0R
nphKHefCkGabgnhpRn0lPQvkVnHtiTlPeQQbDzibGnOuLJsbCxftJqnCY4A2wpn31oA4K6SO03dA
u/quypjr8MRZIraXEN8sG7+A/IN3H29bBANdUSaKO2HacwpapvJNaLE90iZlcqgwCJV5DRFioPCg
yHCeU7hnIQIKCakJ4BkKP7a1ZQg8IhAGfpu1suL5k+4hl32d2x0Ndz5p35yvANqHIJ/RnCt9BkoT
zOYiRiBcHIy371iCirBY2Tho23xptj0JidM8ZhpNeqyEAWeOt25pAMDNmXgJpJ8phA2fklHzbuAW
yBegayo6kw+ku6Zuf9k5YuCJ4emVOo7f5a9fkLnw4Ek09v9TpapKYf19KWW+erJpGcYcdJRyEdx6
i4gPQ3OsDZXJzW9hw78AewVkcfBCWViok/0PAoIVgBiHXo7Las0+aJfSUcdau91yYxOSeTHSlMQt
0Mt2ym/jYzQan0J3zzSJBgCR9LEqbuM9ESBq88KNFCTD2GTM3IibFFP1oOUHMhbWFOavcDxkObXv
GMcLTKOyYmaqhEBbbOU2SWDBV9r5C05PmUARro3ywBdeMZZZeAZyXIIT9EWG8wcXulsjA1WH00if
Qv9Q0bwgL5oHO/rA78GpzDb51bGG9jbIQh1SfoCEQfVIpzRIs0q8znlRR6Y3bOr05uoNBKgXiJyi
ypuwh++KXYQfwiKPf56Pr47jtujbquoUm2NtidJjGh6HCKSOh7fwQi8Ahec55RJ4IXhgqTlGfyJN
vGO7ykqsxNClwbo+kpmKwsPK34J6hBtfG/d8LReI7ZHuKnS3OXjOCuSrr3Vm5eHD+HN8N8VH9q0l
eAYqKn65a6Om4voKI8tCMxDJM4GDwZ8WzW1F+gAhN9pZfKkLhximfhgTp2ggob2gJ5ZPkAnzRF60
3drPQhP7tUwe450DunrtAUdQBqRulGqd7sGpxwZXtxmcfWU8OR0EpyDxFRq1YEYc2U9KwMedaZUg
EtSoYIFdkOfTH57GdHaE5/S6Ws7YcaCWStb6hrA0lMwmpWVrThaEU+NNbDV+TH3mBN6nl0tKkNX9
ArQj4kveslB8P3Tsky+kG2TihaSCybAW2je1I/LknYqHWBNCJHRLA1EjYjv9z90o4dxVCjqt9VCq
OhhbU3Fb5BFEZF5Wxgb0+qWu3f3FCEla/2jW4EDGTgksnCA3APOH4Zm0hhJ+T8B3TFH+22nEnr5t
FxQLUhucA1WKWpTuVKsmtkqWtolGO/HDuDp0DkFY2fqpqrOVqKeNlHg127bc7AznvdtVxaLFXQI9
kiDiZx4K+tnJjYRzRxz8i7cWtFHCAV0Ppwpy9Ie3c/TzQCikLtPp3IpioLAltftxTnEdzbW7OLdr
tTGlXNZhmGjmbkSbTUa5G4X37cG3XD77qoDjyNpJs30Amxg2vplXLclsOebJyJFlsnPRG3j3xaQp
S463+5VOncQwy7t0IJSExQPp2YPQSW84D7UeZmcsHdw8EZvnOkCXsmTITLqJmtaXRuemgnPpBCLs
Kv9fxuCpG8oSPkvFOQqlNXuZ+Ltv932xdcdX4/a237tHdlnhCwfizxhNSVgW6LT92No2qVwxMFki
mvCJdkNHWCMGlQKK7xoeXacr/tegmJxNaTAxP/onorL7vuxGhcJJX66HD+9ymmp69UeoAlwwIOvZ
e8BsK2E7ExmlSiautR6UVOnsBk8LuHzVJr7pnHGGbiCdvpgHVMxpDjgcN6/id8bdZx7xhSi2uGsD
+IMK/fwq55JUoSuu0ZA/t2SRvQbKlzGNgry8XhMoMaTyNltD33/+hcP8XCVlk1Qa3ir/8nNik/uk
nzfPt7fARKAdFI/MHuUKxRGT3TMieBEJIYbEv/reUb+d0y7+ZybWXuJ+IqeokAhdaZV58nRnilXj
2H0fNVlfTv3a4QMNiP9ivic7GuC6GgHb3r82t2LDgEI+khWddZMCbWfES2OgFKwQAtEKX1g700oL
81uCbBbBI4KzEqns2NYjFqwzy17Xrn4+PvHqaTBI0ctf/oMHZ/jEfVw+QIO09tiRT6c5bwOYZx2I
VVxlx2OS0JnAcfjV6XALJF97nes4PtxSGDj+A/D81PxXT21fcKP9BE4loTKOptP7So7NlmhTRGvB
1FpZtVdop3X36C86/Pro7u/3irumwzuX4LdADHxgZmJUv3YdWf1MxF2NUQdUvrlijZz3ohOHZh8K
g7DQpyzmHTSiCshQPXRSumVQL3E99LWMNVkthn6/Eslullsil+qG4t5PUCMJmVbersCc76uXU/cN
iuehK/fkQyWC6Q6Ob+jFJVARZAGLjtvVO+vYAskbpMm+WSZb51+1sWxngav6iezCSI8HW3owqhfK
ApPd+7Bpiaz3tSrSSlxac5XkMLgsOQ0iFX+xBTXi915k/E1A2ulDvVaOYqqnOftCPvPrG2VmkXDM
c8p7SyYOi1x7Jg7xU4Qirh1RKM0rZo5Nh8sbO6KfjkpFiL96LK/BGDSkP/fi8JRLTNf50ohZ85nB
0NUHlyYtQC40FkbgXhsQfW7h2caPoYS3A2keB5TlbkHuVk/wWLPDrqCl4piVg+yGpJVmrA8maoKH
K8XD6qE/iRU7EDIcG+eFuvDu1uITi1jhPfWFRbCIsXtxwV/bqi7x6wjFHpG/lXGaeZ3eCgn74KgV
7p1YuZE+IvfAphEMZLXsyMhsm0GzeOOIPsdjAzgPbOAFgO0XN7qcKUNIEhRUTpVppfcvpziKeQVu
EvihehWY4MrLIgdqZqp6qRKW0obR87OcjYXyWHhXUxaFa3TKkEPBFPHK6kHdDQfNMdbuJP6OgNYW
UZDJiAVrdZnP4ogQRXSl2BRD/k8R+eWFpgqZkuCcsGmo+Y6uRmGKpITfy4WgKZYtel3GVVhjHA6l
GVsVA2Lo/i6SjXDEkdclSiwo8BafI7KUCV4JUHCrA4yMiB9mnpjwnQaHtfG2owTi1McZ2yG254V8
EsWerzr18ePH24GTGIABDZdphtWt8p1s8V/SNaf/JCYpKeRC7aFP/z0lc+zsIpjYYFsGRiUxeRA9
93a1mt1RkSzrFDbRir2SRlREb91lr2B6DWLrHP9hdh+8hw+Y4XZmpd4n+tK0wJc/Em2p2Hd+7+WZ
ZwM/2y69gWZ0NDTJYtoFHnFx/HLR/PMQl4ofWZ8lhgVU9u3jU6acAYyr4GUi5V0tacwSfiAG9bzo
YC/+zqraRg9ju7MrOpO0j7ljSLCO5Jw8hDVFw9pbEXAerUT9HJY2sC/Y0aTFPp5I+gatrENK7gSY
d0TwQJTeMqjt+bMkp+k2QcRqNHHGepqa/fsNIijnzrgcGkrMbI/CvyPAjrjfvfjAzsAqOMkcLlfx
XjUvMrIMVhp5TA1Gwb9Toi/Z29KT0VZqAKDre3h9mkPZekpH+MAAQ8fTNCd4Q0i997Dch8n9/jt1
2l0ykdVyF7cgVd15RxFr0ZVHsHoCE3MM25SUPaynCpcBDbZmRkrQ/S7x36t55O/CojUljOpUMLzT
325tXAbO79aEiyYRZAk8sJiMrfwxrz2O7DodQu/WIgBtcupO/bsArBXJo7oQqcUiQTeacwWomU7u
X5P0+73xgkJZzGy8EDB+9hrcNiI2FSMcjxcGxaKfmFxqwg2bvr51XFG5Y5f36SG3EkZMhazMY840
FXiUYMAHfJo0kSTI+MkxfKS+k78ajYQRjPP8wOi5YoskR1ghYYPSAE2/CvuzpaptEdjxyHl9tZ04
SBolFdIPQKqs4D3wpZZGLAOT0miN0f/xLA2dAOCzmNGaGt2Yx2fB1Q3QcYp7ioKyNx+RpBtdjiw8
XbAsN6SaKVglwAW+/2HmyUToOnuxy5aaPrD+l37sjQdhBAss7yfzDdNt+tsJcX6YGhQIuvJqMw2f
JnRQrFEnF0LrbYO86LDkRoVS38SrJv2xXElbDWgn9FRyf3JLeJlDA3K2p93Xt1lpvw9A+qNXzd59
88Z50Upg+vphopQRVUI/5aASEUviwVWYwa8Y4rHZ+TiKrD/gPAmt0Bybd2PTPlOtrfCafGi5LXqH
vH8rs5Rwe/5Vikze+usXl3k7GBM1fBT8ZLO9h7PFMkVXIVy6lSEIJYJv8oNm/zqUxNfu5XYapg7B
cwt3WbBq/lZelT1RT2N6o+KIgCUiP/TrPJLIWc0Xs0Vz3Uk32pCTYJc7mVjO9beyfPwfnAXwZDBU
C+IoE5DLvmehtMPKU4G7Z5oK0Q3YHGKZwkvniHj4fDEsSVE9ZYIukx49sixXQVQUymrFnSbmVT6N
3pPiMlcN64TrqCGcNG0RLNfiGqOQorjaCwqcZj1YEO0vSTgbQL4sFwlEBFxCHX+9piMaSf3w/Bvx
UpEsA8PP9DXN4P5lfEFL11gUiwmZloj51/yJWd7H0lM8HC5mCfTl7ofc6YtnrqR5q3nqMmo/afjb
553P20rmJQBKCv6EWQ461Fss3hgT6+Cl6rj9lnSY+EZVCUiA12SKU9yxTPQQNFB6KqX+RxGjXX8Y
wBLDjU2MMjVw36oiq5a+pwSUCvc/xcDDjGYifLhWW0siDhK6sOrQLMNUcbjRLY/BpXvadQee2K/M
MCvSLDdRSdmphLAUYkIYusTUzopp94Iypqo42asfB6mSraGaaavBntZYj95SCpB9mhMTuC/1dal5
XGS/SGc2tboKmR0ZJW9Zo0sz98GZI9CeBHMcMqFJYqegxg5aQ/B8EIroHF014BymNy72WHl8iRYw
zdpSBejLoiS2X7WjzdB+49c2N6QnjrVn/P5C8Nm4cR5PrfSlGivACBaLUGWWLtyL4W+eSHFsDSsD
jk5O7vA786qnxf7eyiubarmYAT3tpionCmXJ5/ZE3yQ0/sE1lSCDru+8m5yJSxZg2FHvueTKNyBu
S3Pc3q7l5v/GkuK5dV4MkTVle+lPusR4svqgZngrpUbPXuDIFe0Gc+kKTr8x1buJHPIrTD92e6PG
DxxFsQfcOa4hqXQ/hKvsTI/om0QiaQElEFHB3rCtKh4p+deSx3XBtFvizHg8waq9P0+1W3WAfHMN
kKa0MvnyoVl14Cti1PJ+0IQ11WkLIHwupvFziy+tYGITZXXT2GcYzv6+sWKRmchvJ+mOv44XSTGo
ZQv24f8zO9NOGzwHQoa4MfJsRa4v1W/SDcJNWxRo7LEH0SXnjTS0Tt5m+AkMtxrMTTqZLDpWAMT+
DVTk4jq02Ann7GS0Ba78mh4qvGZQElyi6wPC8XBVzLcj1UfRRXyvkSXPSXNnE2J+ST6WHIkqAS01
iIBurmdEwLPxVkRWTYtGs7/MFnAyfAsIPRUg4Qq5Wjlarvhw6LmR8z23vQ42fjJpVYfLOtkvx7AV
cBN9iAn3/8uiT0xeX+daGfCd2IKmEQVXXhQh2k8TMv1jqmbhZ2PnN0QBrnUqoKIZaczra/efMoG/
9hUOzKzF+6L3g5izZQ2ENRQbb8OJ8jZp86djkPxjFWpjc1RHuAZAn4se4gHbZpBixlMuCGrzgNby
MOxFcwAr9NnASPNIdiRcnNJSjbgXsXSxJQkvGAoDLA9TZW/wuLco6xkyp24Hb8YxceCK7fNuDXto
sjD0mmxxZ6s5OC6A4uWoONkDhGwkt8Bqwt9MKjDX+tRfCkoLQNe0RgxhTzd/is3PNdPQ/PVXBhYz
IaDLD0Ga3csbSQRM5IpbInX+jn4MXVKvUaPJul49AlRoi/t2di3OK54GCyCbUMxGVPJzAFKYdfRM
6XjCJyqVTKSQYtoH9IwfwlqrdBkuWDyDVP/+hF/3qJYCWrcUKkik8tUHpyW4STGjS8vM0M2C9g7X
cLlmJ9s1agSdW6s1fyphiFJ7lLJa+rZhV8fuoFa92uKgS9PuGWkhrDGa5T0Lof+sENYGc09ZMpjm
k7h1Xmm/nhyyJzrm0rHLLOdJzrX9NFgPhokxhKFRgfsEIAYhuYssL0SSKkZOVD/BIElmJP8iUpp/
H3SCI3MYJ59M4dBQ9bVcpi/U3TeZegxIqbGV2w7ihJmJrDQnYMcZUuSngfebjyWy4NEozaMcYcvC
sp65cJuOn2sPCoBlxecMQ/XkCuu+1l6jBi6uabqLjF3DAIf03sQJ+b8z6ZbEKCzp1QobKHvP+8yA
2t0fe8j2WLkf4D6zTDJYXWZ/0A/yW8YDLduPGh/ueEjYxxnz6/5+o/HJq565q9flmmDVt0kPvePP
257ALtzCZF3XCVeNyrnCEet8Zbp9y/2DvQ9O4U8Cq0khqURkZCr29nHhb0WBE3YAVtL8xnHAY6Pk
kHcQX7OGB/gQm1xBtfUgX7spL9cJV0VEgw6WxMX5/vsevZilanLli4RdukYtSzVsS4ocrQA+fanj
z8BJO6c/Qh0csnexO0rP9lRy0pcQ0wQU+438iwybHaZDxI+pHOG/FkHddhWzn6LECCSKKSIi1cLE
oAgDXo4X8jnjLJ50RQtF9NLUtq2k48VLjZkeF5825wIGPGfmEGHvSkdd601pPYpG75BZgws+UE0H
Imsfyzf0rIeQKcg7H8yrs7lzeOgr1XJCy+cjUQV2Ujbeu1FsdT6CPJaYaczGcfGZH6tTIoaE3waU
p8pjdTbiAWu/rBRCRto1x4wID5iDtPMCEVu07dPbiTdC52IdOrhw2GYK/URllGGCgd76Ym+F+TDP
kzr0NOY0yrp1rMDUMQKCCWjr5m1ixw+mGUCAzepYWiSoYh0MHDf5BKm2m53B8iwLxuViC86icv4z
P7dDQQnehLnycLu1XE1sFN+QARadcPDJqsXxq/FUXR3F/du4oRFQ8zsR1MMz4cPDajwDXNVB2AjJ
2NVYWEo+S3kfPqRrSTN9dyx0SV+zu1bPrLtKwW1oSoi+w+O+lnoL4MPxbIRDScnLtHYedHORZJtL
HxZdSNMcE2sda3FJGVkWr9XNGoJOIsBJWY4HhxbumTAH1a9Y9QiS3IPIng7Hv5p4XJpHRRtMK0BY
uApMq7wtnAm5uRJAZvUCvkL7jitSvMXQIxZr3b1dBG7OqhmTP8RwpRlg90Co6He11fn960KpF9ZL
yc4UZiMajvfGJLPJ1sKpTR7TtnyftkuhG97pmSVeGvUuvs4/koKkmJDPhG7IXFxobxpQipodMFPz
hrWjusTLslN5v4D4lO56ugeCG/WE7QMzxZKz9RTA01DZkMaAnAqMP5NCQX8639y+xBxNq5SNliM4
bqN1XOUmb9EknctqU0VcI2E2osNyfeEL9AqWevQ1KxflUv6mBlg/kOQ9GLDA29fBwcHyt/C9wSJr
Ln1OG5+dAb4I57z9ZEw/J0lRTGJXIKOTbymRlyvlSSGbBnLWg2MOnAerSxqnUZXQhSJDnDOCl9t7
dO0nchAS5UiJdPUmVsqy21+1u4o8TPKCV4NHQqzFj0qwKyTOCKVtjemENjgC1N4Z81uIS+oLGGNk
FXQahWUo7fSs9Lmu+mCVqv8DD/jq2V5B3PqwCMw/zZv+n3yQ00+hOTQeGBTH+6XxXEXAQ1vtC+0h
g8+Q2K72Zxf6+k/zlAeC7qm0kWdadmdtwlsHq48dYdLNAetFnpE8ILfSAPTHq1TxLiCfNX8Xmf2l
wH3eQbXdBPSRUupg8DiA3T/JNydhcoygzRwlFPX4aoFUpn1ug58MAb1Ugk8XTdPW3XnDYJX77kf/
CJQjWiEi21YMPjX1FT8VeaOhojhxI3Nxat6CMYUPM6wdK6JyQgcZ9Kx/7BsKd4WrjhqpEyhvZEB8
vAMSKPFZ8pcWpu+Y9Kvew2KYG5ckFEQM6+43dU7zVVHKIn7uQRFl4joJYRrZhe4t0LpLiyhJGCJ9
WasxMBqco80WZ9aEKQZN41sq4ara+3BloBqgK8E7aqNlM/HKpdSS6Qw2ITCXU678BN58fCrpGZet
EuERrrNkckWBf9UCqZ8bzJRvYdC63uwK9qH3fOKdKzp+7jV+sJ6J/qpq8ZlPUhakr18e6vMDbBfX
doatV2J1SzScg8zIvua1D0k3TMqaswvNSIUS2iz60Y8Dj7Dl0pkobMGSG4kmBcrmIl/m+hyBk8XD
DywDVqntzdvWDoLmfeqQuLbQD9vGRP9/BZcctkatirO+O6fHI/qcsY5jSK20Zu4PloZYFi6tnO/8
K1HiVdOur4hvFNIYpn1+IuPGT7ERuoy+CMyGsJYVg6mrL0SWe25xJhoK+O8PJS6nIAGOWtqsPZpk
5hvHacFQzFU0IJcqgI8kHivUoIh2+2tzYnheUkSQTCT9Njlc8IfQUjUbUNJAwQTjIH0fVOYqe8Ve
AUt6Vy94SAKG1nT4+eRlkuIYCBLUlwXwycp8YufNUrnbi1xVvjkDFCpEnSAXygeX89cWXX+WEq0u
f+R3Q/s1xqvDtES6aPo2UQJhecXSy3mxVuCGilhPKT+UQ/Q/obMni/GbPAiaaeTnICe9j0/ucq9p
VJK5mjnbCyWy0wM6pEu1jYi3WuoHapNrXdC1WDmi8oZFvz0PdOQyaIiTKONNrHWdhHGzJkFVBFLK
m28h2stmML8ePpxh4WA9ALRNpBG9YN6Njpnsai11rKan1ln6+zqWTSPXdKPQvum9uR+19Qxe87pu
xI6O2V4xtdjQBmxGOoOi+Qh3xF3mAuMn/S+BAIBSW91AThoIVW+8O06+7e6jWMuFLGpnSskARBsD
I4MRUtPxmayRqSEwHeBJl5hCPmhwbPexhzrDUOPS6Ow/ZIcm7q3bIogUCqdgi0GTKI1YHH9hUPLm
8ObHkxl0cdhyN1wMXsIMm4MiYuLU69z1+QAdycf/mXFOhB53POHFBezBqnoZ9Z16HdUyU9tN2iIR
oNayqAE+XBjAzau0pUjGFduopjPCNeaQiACdWBJ8gn92PdJRrNeHdcESgrsoOhEUaxLZvI2dJFOy
CAIaVWgCGaksWMfrVPbwx8TT7JU45U0ONuMJhQlw+t2cBRZ3yj/Xe6W8fByCNImrXPh+Z9SCwsXK
i31T+yXYCZ4nShYbq5P8sFdqLLY8d8fFRnqjD/E8dBcmYg6r1NkrVR/rpva5RzhrRmCSVurKVVSz
JP9kMJOLes9n7l32hlcYktbwjNvO4eYUGqiSYz5ipKvUJimw4eyzPjTqcWAmhmpzwhwtk8kMzgrF
nVMEoJvbuaKf9/EOAHsz8+cwe3/JMQZ2IReVVNxIsNoCayQahc5vEtIZGPJv2UCQrHyrbfBEBDUL
E8POk+jHrrsdu7WvyEER5wrkXYqlk+9/AY5e7aZcsLKVdLYb4enGEK8vBbjbi9RuozZME+SsGXbB
hhl4ozFnTuQR0voBgrlBEoE61CV9KlNKegE19UnCkPCb3CyEoemGfPBjBdC0EsKMw7x1qCFmeCj6
6u+9+BFObEj3irKytIbNU1Q9k8Dv1g3s066m+W470i8IQR+PLeo4anSazNn6pf7h4qsbo4X3uuHJ
E6S2nxdAAF9GsniQcwfTjow22ZDWp0FwFQprTabYxowunOV1YhbM3khnHB96j3flERKogyUcYPla
hnUjtXCHWZukD/T9424lknWRW6kUbFdQ4FbZDTbj1R4/6ukgJR8icR1c2uy1QfCapU5Mp4i/ppXe
kgzTBSAq04LONrxuWLIHpwlj6uoKlSA1LCsn0dhm2qMk2tlBPLeeRNFWwfZfInvfZnE+4x4TIeGY
NpRt0GwXAXqLjgxTlw5wRbdNrS/BFo56HAtsKGI96eoohUI89NT7rBTD1+nS2yqdrZ612SUl0WP5
ozrMGNs1ELMxdQfbehZsRlKgx+AiqYUb31paWVUcyPImrB9BltVaiYUXpC+/4ReQXO/1UBVMInQz
f/JjNCkvDjufvK9mdEd6ar6Ot7h1CCeH5zDXOIixbpj+aNZT+pKFF9tfAKdZtEHNsKOxXwaB67FQ
HTUCmIVxpdAv+QFDX635aoPrztR51bd8cE09PDav8wjODqxBM6zB25nvhaO+ekC5JGPixKXNPeoo
DyTpEKqDVb/1S+wj9nyBDOH6Rwpxro1jnMS2LumSV8T0NolccgQXHfMvNDl8AFlvAq+yv4HzI//R
BeSD2wkXTUEmtaJtaw09Qn5lRK+dEznpEPuvtL/9iEMyfu5PSqQ+/kXINAQacreE9b0jJjYtRuG1
1htn8JkuTPDt5M0C+L+ZAEnubFfT6O2Vopa81GIB5KG5sQxE3OogX4mBql1s7sXa68xr5q66KftN
wdgQ6wwokv7i4oS9/Ly0FLweWl5cevn4krjjTYgIWDdEpvJmysOoC6XB9lS9jfXuKcKwFz69xrle
OvI3vHFVcgsEMMJ0mHzIy+FBx/iG3lwpO8dlYfZL9yLnFeeIR91Cs+dzuWB/b0nBSrVDjCbT3wM5
XfCyzqAC3u/PZtyn8+tdndOYaC5EPGsudAEbQcXQ+VsEiYqbmVZpqVp4gcQZgYvY+2rRp7gOXMsS
xgJzaz3CsWGbNnBhNVZzZTgn7rxTqX8M1RrY6pGrItCtZlxFthTjbQAf4sdA8KW26ZzFYcfRMkaY
rJzROQbmsspUSLMDXMev8Epng684IRj3CsvjfVM/0ZjFPsf4lDd52XxrhOB9jZpEvr2Z7PwTQYVg
ELn7u3XwP3qcH97FkPlClhFdROsqjmXkYxW2XVeZeLhctlR5VS8ZEfd16a/k/7lPbv8theic0W0+
dA1M5ybhN4Wg3Y2y829G4y4hU6tJ0uVNi5P5rDA9uHGeuGtQMIUXHdjtjBMRNevFwRWjpo6IkpH5
r7quBCR8RFWmjD/+DEawdi6VrqWKpSOCMY80B8XC+/lpIuK7i/Jct1cV7Fwto8Sh6faJgX9QB2CV
ZWydojnxNpTmj2Go+AgpQxF3oVq1/SlxkjC53IdQBAnVWYeyAFsiTMyKXk0kyVqBjSSC7Z4N1qKA
eUeNypSiFzB7IRDH7IrTQGdzHaUMh52Qb81FAqQEQ+kzLCnOlFuX/2XZN7cMfSFIlM/AdzD99xK2
biU4I2N5Txm3DLIRwF+ASQwdDl+ub2BCtGHvrBCYbhWFAJWBAgkxZJPjH3qDnD2TPmDwh6oEhyr2
ncyEgg7XOTD+jrZ+nqcfGap4guvYXwFR2Z8bDRz4dP/jmbIHochMy/w4TUviog1E8HWZ3CJku5Xi
vb+oCeSRKVvmhe1aeJshH8CaT3FBKY8GfMbTcazgqhbxYvPK6oZmMAX/+RuBDe8Zny8TJ1ioooea
6maCZgWI5TCyOECn5Xr4pZGdEI+bkDJxvLNe02NkI2eBNV2/b1GrW/iXQqApnDwz9UxHD2N9CKyQ
/JioYRcDR3AQo+X7T2UOVWbJkbyqxZx5GR4DHYo7x4ba1YYEgrCtYZrXhkcXGA3fo06kWeld9jjh
EsBbrFua5eMr0tKFb4BR4YmqmI04o9rg4YAM9niMIWiLPyoOqcBEn7MqAjnnYFfrjCESvBEJQYyx
WO6q7YDDemZq0qqih6ydXLxKFCGCIuXU2hcznxcPEoju0eNyn9VTKIj+PVTZSWFCq2J50EO51aiD
3fJgPBIx3TiK54/PPOsJFdin1EJkMbLL/4xyt8ISBdtLCvxTbya4uMvu+cOs9WZsVx1vXh5LMjNB
xsPq2AsRRmZqeFPrYF7oTTMzlAIULjBjz/hHMOZS1O+RWzlDSeeWrfyGHtP5EojumEJFsRY4EcLu
5LNEuoS+UWeIxMAjMHseJOZcYGg5W5R+L3B4I4MLDQjL1D02RNU9cmsNuDqzi9iTtk0wKeQ+AGrm
kfpXd9iwWb1dNgnH1Hec2PA6FHInZd+x+BTC0f5KQthpymvfZz+YY+AcOH5c64F5eCzy9eXWDzdu
CCW2qC9L91F8fN+l/IzwhVRXtSNqfOQ2nttq4MzM8JxJ5R/vLk+VQ+G2FGI4OGsTFqBKpwCGKKN5
VCgx8eQoU5Qk/rY3iGIHAH24FQAffjUAy1L179b4HASIbWMteZKFPncVrC/IjEAwMXjGQ5TAZWmE
gwxEHVNVxZSCXMk6Y8rQkaHYdx9Yo8sqDrTbtNcZIPWLzw4OHmSS2//h8gD4e/QiBXhepc6C3pjm
R0MVQXHJGIBCMx/CeZffVWYEKu9GR0lMGe+TMfl4mE2qvcfCl+LMnnq8z3kP78QSKcjKPxGsYlY6
1YqISS8iKuRO/6yDbFeHS3Gsn3Ys0kuFkWPMGJ2qPhqmgWdN0BvANTDjVuZD+Ufj0qWdD1YNJO3i
K+V1iDPiaV+L9lgwtGeOATppN1eiOKHWgoHSbM13J/w9HP9r0SvM4CO4X/JjJnf0iUCvypt6vjr2
N2vEhmgeq9Q+T82yVMtafZsQZUJlW5/BOnn68VOAAOhSYEAzFsRWgxJHLC18QNL4dBelCUYtQAhQ
G4Dk9bFjKjz8uihQeN8IyWnUFS2CKfYXAJk2jrC51EUV0R4Y9qEitcCCF6Q/27pz/pD4Qp8COB6E
62HOLksjEEtPI5xYzYRWAVeKaCTb2KT5tMBykxFW/eIgshRpGnlL4vwaKm/WU8dGU31YNs4h0jZW
WF62W16HXkjqg1C84kG7B2CfMPGfoH/NP8gxnRJRlI+zZIW6/YpE1NQOeZ54+7hjkc+lcpauYTD7
fO0ezYLMFZhBl1vlJ5Tb3xEIMGgqbR25ll08VlS5ME7EQlBmnS1Dnl3BwHjWSzocx8L9A87RK33b
IN9Tr6OYw2RVKSiPmtavTljQpXZHmEY0A+ydMuPPt9E+3e0keGycpfeLSj98F4NMuxbL4JvqYB2n
b3o2f735HIsh7NFZOYBuZBjo0XFkxvUdbpXN8B/uEeJB6cLYRwXhQTfZ8kMMma8wbrEAI6S+Trxy
iBApGMpnkWEzzqsDCp7ABSyFB/7ErfcjDS43CJRdhGD7/jrGAN09j5PQrTdqd8LuYaqmFgBeQ0xa
9VlLgr+2mxe8bwZJQ0howMEqqUsAhmkZ8DJWgqe08w9urF3YUF2nO0sWt5bg/8g/XInM6EGkZiPd
r1ZQImFLfltkJnQwCDHAVwBxbfSxHl4QwVjVSe2XEFTA1egPJJ55YEG6YNqLhwXeQ8zJ7e2E1/aG
OD23INJInwpymihz1Ni/M6FRK+A9vF9m8zJv0PoLjsqNcTHCWqWMjSETEtsCRT2eexOHIZxMpDZH
e25rTjU6pKUg0NzbX2w1635LuTabFk5FtgnUzoNZvDqRHEDfp4aMBegU8VHuANK+X7Kdi60xmzQC
j+w/MdO+iot17NQHRnxByrIL02Lc5NP7mdtvdrDNmY0Dfn6/kTO6eaYEy//05uo/91ot3cwI3sfh
x1NZH1jIqAkf3drYcIoptjcdFSm9IZORvMIqt390rRfeTQVoFI0mYBDy+sk9iZMnHHB9FspnozEb
8I/LgzOdUxS3o+EOM0p/FJkbGDvl8fETz2HDATfY4aiCraBLEZrGdg9uqF6kg6dVJr4FgrT/kQUa
8zqX992b5fVpfhEi0BF90FUt6gsa2yqbfD6ENqoQbJrtPZ2aQcvi5pruWdouq5pJCNk/Y+OrYE7w
S6I8NgvEmXtKtlazTLWOdt6ZmHyWRFhRrSMqdq0viaKFn5inwCniwcT3fkyiAYNaMEmyePP/T3VJ
8hEPATfi5D7swApGAmBrEDHl+4Wmw5NEl8vQ3glpPgHIk30xwl8dNAoXSqgTQk5TUWmKeNQwX2TH
EfvWmma7+32IoLajzoPUiFW8+2QrxeAfSszzIGrP6mcNue9ZOVuJ/zpgZirUjrKomCJS+ym0z6yd
cBOGth6h7moSncs2nUVxq2874F1XHjiQ+szvv7eYV2NKb9CuSxQ2OK5xlFCqHB9SMDykactcdzna
RaQvufgw9oldZhYyxax0tZ2Ra5DcPsN05RABywildHXuGnRPeBZ1QaI+kycyo1CGX/fZgBoIOKNc
NwEU2ElAs762+2Fy1d66JiXQEk0Fco9Kj2p1UvseZ32pDIlG4TwFbx60oFBU2LsOYFaTXhH7QIjV
EPVkLq7O7B2DdlfAUktyRAB3sskrIuEGKNGoVK/389Ot+w6vDayEixSvWqFkFYun9SAjwUgHvgk/
jArofINoGf9j/AZRCbzQhn1wuB0fK58Dj5EjtqdPTozjpVCYEWcw+2+uAwJeMyglxeer3lrTWVgI
Zh9tg78k1eey37dQ+6mSm3Bw6Sou6F4JEQiseyjY8BGp3Ek4+wJz3HSbuSlgSXdEDe8+iG33JpOb
EaF6Q0qRsyEne52YPRzujaGEzK9fWhqjOETRC+LqDV52t3tw+g4AE3MeqdP9xa2T3M8FqVJCMdVL
6Bc93O+dRy3Q2XWL/4DFN4Ypql12Yp7XaT7WlhGbyemjPx4xNKkcGPLoE4aLQFztfUo9pxMA4G/s
hnEtozxtR42OQCAAj2sk7woTwSq9uEIsWA7iLM4LjWmL5UOqoBjQuR36Q08N2MMHwCgYbkZ2FDSd
sMRhdrq142w1gPN60OsGSFFD6jE3F38wvl8FDfnz+k3RetjIdjHkeFobD447/vzT/Gv1PckNv+cm
GJrGTkmu1fHqB8LigD/oOldiR+YCUWXpSPK9hNHriYT20H/0rXk1BwHJjXF5yqT9JWGWEHC/Qt37
eefqutFKkUk8BrKh2CFr0NNXCWMSq3P8LEV3QbbGjKHIxOLGCW5QdN6QKuukAR33OCT6K1sYbUJT
KIrckISDTvXOhQGdZBPM4yDWHwp9d4zEZGnwZXGSDNJMsl9l3RrRRPKpw3b5XnVe/UOwBmyKwRy3
gIcOoNIw16d7tvrI1rugHbsl7Hzcj/3x8WtTW2s4Hf2sEC1B3WFQoHnYqsXOWs1WreyjnJPeggvG
s2ki98A6EmQOGUGS6UV1+9y23KjIY/EWTl6Mm8/HgtfO4f1ZZREgZbY8Qe5rF7MaPCEV3MePePO5
7KwQXuIKdL/0JV6TbUK4qn5r/Ihjevp/YRrL4VX931gfAQJBprlz1ptxqh9CxKVtN/LExn1wtKml
pO1IQVr/qr6Mzn4TD5Mw3XhJh9yYCKHcEIoKoblYGtreejNrT37ka/q1vtkLEY+PU8dTeKG+DQ/p
vBsZ8HSCY3WBSm7/IgOVKw3peI3Xlfp2WXpXZFV6xL2cbYXi4O2V+y3NguYGJvy9Me/cUUdQAnAC
iT/V9yqQSwc+tkZvPxhRoJVq6gW2yhxynryQszUG4qtalJw8V229XmUY3FIaA+/fbukU2LlFEw3A
iptiKdoopK0Z/vOt+mCzDfrFQpT4pX+bUCmR0y5AC6H0VJC6KtgKlBWkPFAKjzKUSGfn5XFvMAix
m7+kgdlsS7ptCYNM6DFAb1XHolSkYN3ofR5Fha1TP9UiEcmrl9g4qP7DNN4QRdYtqTJSZ2fO2QDu
LweJXT+zrp6urmbtYLc9LwRmw18RieOXBSRbWbrcraFH6vKkluHrp5OZl76c8sA/fYww+TtZ1Z+I
u1Ju8vc9nu8V5y+I3y7yAgEI5/LNKsl1El45r/3KtGvVg1+Ozf52EeV8FHJvoQFE5px/+Qu+WaUf
D8QvlKU8U9FGnOCR6I91VFiFz4V+5c9mfQs1lXQilHz6Lm8r/XDpt/cOVFWtKCnTYxfhtNxGSYNC
QpATh83qFlbIqTD5jUx6pcfhuEBv9ApuT/sTblbjF2g2ETjfqRFMrLN90y1ZJSkIi5FsSBwP9vdT
hmcr7MQP6YF7d+H9TbS4muPGcb9M7qR6Y2Lst1qx5RedGCjjZz+7JiO9lmsr1Ll6wiOElCHv+/Wj
jGB8ttVh13937Nbor5IMJlIsGpMZ/Gg7rdcL/uw0ICvLNSaQa6G+VRtpvPMUR+NCpHNLV6R2WQ2R
V2C/IQSvrMOWv3znw9ei6EB0+XJXhCrFRUtJ4G/HSk0/2UAltE/ksU0nh97TIbtKBci1E7ub7Ygd
qc1p6/RQMK/e0mdVhoZCX0ZXLZpvSfCq/YGIoL0vSeN6/n+8gJo4QUT7eo+6DAwendWOh1B8cdmW
NSp7w1aaBHdSSlzhZHaLgiR+IHDKOOqo9LIt+fbe4p2MJKd3nR7lQMAgxpyzUZZ5EmHPhEijjxWl
TbavwGgWXNvJiJ0fLF2FjLGVMJ5oLGgy3T1iGhmtWvdmwaNN/1L7KaSOboyFNOKQ4clJzqxz1vY6
sDVUUP9FIiuZkilJ2+/feJlrBzyTRIhvK9ZTNFYyRNj/qyXmHgBT+feUltYwWMI35nXJfyvibaO5
ni33Gn6jdHFSh5XMiUh+Yiiz/x7AfYAeRZQSTydDLUihMmdx93jEsv7HGkZTnlWCzYqIAoor/TBq
SvXuRlBflkh2ufHV7yxinVZ05evQcQIb26+owVs4fTlX9jc3cQMFbuH4cL449imqu1dgPVeSREn/
BA6ANtqSaoOHmzXO1h8rSXEQ+fnRmWI1CoX4sl/s4+Sy8INPL49884BCTSw572rqFWP1iPkiW9hi
pgmi9LJUKTsD3b/OzRbVX7DC+nIEzWSrOHGA6oKbEkNoMWDZRbgaEZy5LXbNBuy4lmbO/YMxhYnV
lkt1zAKdoJ0bgjgWFKV0Z3K05MvVHfQLRN+vwN7Xhc7wTgCRazdevFpaB4UHAVAJaWxmZaYlxvkf
9A3DZaOkFar5PfuMz0wYcO3iIoitbvIR+kiLvFfg8IQijGO45PmIJQIezWkFIJ0XXKIhe/MkT11M
PES2Q7CYoNBLiTHzRKkJ00jwoCNPTaCqW0aOTndHq+vJZkEALa29QBBht6TRDEuHFlq/WxMFwLt8
DwklgYZiie+vAx+9n+2IgIaMkRck1wfZgkuHLkS4khK5AjX2376ZKFyYxPZD2EjRyuKSFJh1kVlq
f5t/1huLkl4dIXQT8bwRL1U9UuXdmUpiGrWqEI89+DUJleYqFEnkx1mPbFQNeczewuCuJuIY6t16
/LzqD+roDk/U+FlgPNeb1LK03froOPg5zxnq1gS5+n0ra61TT7OeCv21zF3QL6XDVwfmQ7EEIYeQ
PXAf+y6pJqr4KvSVt8KA19JbgdGjH/LG/6b6doFoVTPM+okq2c6kuA3z12vkEg5rVjdIeHe7cX7M
ux4NjDHFTXERrg//mDpk/eYcB5FPgb9OEbPztgqNkdT7YFZ1xIpNSbnrhJMOp8/J/U23vOlUfxSO
V4LIah/C6n6+nNNCRYoh5TOl7JrjmMc2KvOxss6lAkAkNZsx9WCrZ0C/PdKScm3IzrPEywB34Gz+
LKd3WqN1k36HOOeflFizjWgCCWKAlY9tIU9YTKDYwwLJFiO1sjqralT0JwZUgd2+wEt1jgS08bV0
xvsXRr/mgCrLgT7Z9gaP1NIqiX/W/xgBgKbcD3SWg6Z2XMkVzEKFgysDefygC39nrwC79npZBH+B
QQ+1lIjOgD0NU5WVMYIv9oCPaGLBbBpnLoRku+LnGIIpDv0AGpZHezn+rEtJP6KJWJLwt3u/0vRF
KwtnkWmOOKV5mSR5geqoIaUETUfiBgRKheZR9LjF4CaK6GsREM5HWEoqZfMDHPMdTb8qYsH/FbW7
9mL/SHdz8G9EfU11KMJ/OLfBLT4HXaN0Y/s/gbQiVVLHPW9TnNK7MKAeUJgui3j4tJQz1S95y2kB
ih/I7YGhMumnNsQd5oKZhnYfykqASU12VHFyuQailko8fgqKkLsBbC8usfg8f1ekUxhV9+vro30L
nsjVePLbHpEMU9dbCDqiF2RqC15YsfTDWiX+6ciW5KyhRmKEqWwi5Uw72H8PXdL+K68qpzutIUpC
tWzjERRU0EMM8B5uMm73cyHGIfE58JoiVcGJn0ZI+tR2K0LryDUrOE+hGFDqQ8DxpSvSZHPlq+ws
dzZl0igMtTm+OGD13Z6BPQM32fvOa6g1HWWgHcYo7/QLHJOwHwlxNBeCHZOZe3V0sFwS3Do5Kg/1
1H1arA/O/LqZgbZE79cYY8SiBzait2SCx2HzPx+Cf4aGWKzXD2MZlEtgpCUGjV52IAKr4xVEp79f
fVQMpFGi60AUYesUa+Ox3+x56BD1eM74tuCARpCRxusM02DBBg0+/wVl5mqN0fJWWUBHLNmo9SHF
8ltmkWQjF0GY3KqyeBqdvdTba7ID+8wHktT8iIDVsB2gFll0HfuQ7Y7JSJusl1epaYjfelFijK+7
VVLJiaLb1dW3JuKka+euud7yF81aMhfCyuTM7hN5yOpe4f7vkIx/NVyoj/sg0SbqGyXyUjwZQXhc
maNGiWXi/NdF9m5AF3SISZyBkuhQ/ynzPtUwBN5FXQU64YxWb3CkXURyNSoh9eD5S7OaZmav+wdj
1vHzpH8a/l1ZTR8YQAEe4DZ4nlD3RH8t42PUvcSOAHbmp6Js6mq/Fbg9H4/zKMxTIAaNfpaGYUtf
CDXQoWn7POkvG0AUTL8kLd5zbWSJQNEmEN814ukXI1l5uYk1uCRKK00aPlN1K3IRno56aGDGib2u
rF9B+sAialQkCTRc4iCMBL8+51X0QIoJ+MVou4Rllnj2McdA8N9+zvFHlb1UZIvAgmzYGeIsHngD
c79IQp/s3pj+jkILJa6hJvV7ksab++XIQxZkqTibOjrSPzXX3oUF0uk5Z+mHkKB278ugdsu4J6eu
N6gCsnsOhWXeyKCPAL2f9GPwgConVlqSPjgDVcG/VT0CIAWg0QC5ZZr5qgiIs4WiJIIupBvSV9uK
/l7eGXsI3Y3lNAEsQzoS9vtEJjMshtaLxgo4w5L2eFYdxtQM/uNuZRhbcRx0wao9cJTmHFva+OPY
fjj00+9yCqfoNedrOvSFayJjoZ0arEoeNye8ofN41LYGyM6SoNIbJeFnwvsaqIriat/ZLMnml+R7
e+Ikd1kS8T82qnV1Uhf+6s1TcTw8UNX351vY7l+SH7PFFSjhP4RY04ic8tWAb6YMiP3RaMETCHHv
wsgk2EqIVTyHZyWCzJAAOklzXc7Ii42HH7e1yUl90I9bxme4ZtI7dx7CfDAUuM+HKit0qU9YoKWB
v5ofvcMeJb+WQdwugaRdHHC32gFOxAoNqHdK3Rbwx1B+VS5Ak/E0eC5a1aXJy45AwGwiBxw3nSu7
yksZkfaKKT/a3OmEfb3jLaCcFHUOotblPjykufS2Frdx3b5J01Rh+MrBlO92Gj74Ke9cYz3R+675
tlMk3QfeyC2iRzc2rFlMqxu93RGnRD9PqsYhbZYJ8kva1IeLaYJBwmO9sUHxzRvG1rZBbsC23w3q
Aq+1IKIs3tWvKJdPHIQyKF41U/KYul7HiQ+CixZVg9hkgL4gb1C/lHEJ+Wfk3wtbzv3w7SL9TDfC
CYU6bwLI3tkI35ZMoqfNcMUS4prZ6D2ww/+1EorOshwJODGEtjhMGU346vvmwx/BdmxdGqblxjtR
D6INPqV1nDGsvFy0GARLQpbZEdNb6/5xvGrs1xLQwoVrgvjXniDcorR4D/mFJghGP2wg7ksFtbBm
CyquT1mvX4i2yfavLXpw7KKKvo64dyyBbwlMCjX2cvKcR/h0sPMLW/Vtj+G7hMIyy5LrzupqP1a+
EOApH6T4/3MmqDpasz1zNTVsXjkKDiG5Su0wTOhmX1XbTwGSzUio8kmtcNaXKOuwsGjoDAAP2CNT
zeLMnnnldT+WCUOj3kp3NOgjfKPdK+kLb0fBUYdyKcQSGr5IKYHTg8V+hAc38JzzDEs2DlbaA+wY
GMFzz7/Vq46ZUPk6hpxLKOmYowihniPluZkeR6xlSrr/qr5Hpf6XWl/ZdaQvCy56ypJlfIaH1HUM
ecr19+HpP7YDTLLOll+0dKP5pCBau7sV6kVdf0KlAYZkcQZprV6Tg42+oqTRnK6t7ug/1rEfftE8
R1HVYSlRGB2RXfwaWcqodAkpOnbX9dDPxHTETJaIiQjz+dGMSQhtAYQgJbG5dmO8GCRwVVRreSyr
gqSyweImAmIry+6xW9lSHiPJnOR+m84VtS4bQV8qyIQeifgKzsr3TygnowqDaSfY7T+DwKn1qYEs
Pd8Wc6e6jxlbmF6LdOO9bvW9zyxvauJP3gzvfMoBLtfpOoU79GmSjfKRVoG1G+zEx2Wx0oQ+nufZ
fu7qOF17fwHDNBiNkuVMTXVary+HT+kbRyicRRr/kPsF3WIpNxz2Kf/8B4iTzDaicRwCbKSOgF2B
gIo8LEiPyqVivGVkLTFX+qBIn3vrCU8F/nvzdpIXBX6U/r5Rnj48WOFinMxfJRzmMK3ndnnY+3XV
oTLfqEGKgLRXInY5EH0H36yt2AzpYWtNdCLzSmqtLcVs7/NxnT5M5kagfoLZkc5UDu7OPOSF205Q
qoedZdMY5ztMBbhDg/uX0VEs3LRmUcC+guDNkAcLW/YF2vJ4sfUgSS42SZkJcFBNHxtnHA+14Y9T
tSjoBrRYlX9DhY09rchT3ncXAIYXybgl7aH+SrKK8vzRVwxwbSVEFjw1DiOHn1M1hTOptCy0Bgji
sImF6fK+o8efPLqGAXK2nDZ1C4XSMJFZdpQsqV7It3ZH+3seFnKY5sRHr8R32nhFR6yzPP4KS4Vu
x2VbvUembhRA3521Gn+qv0Q6JlcW3V+WuaCIsYRd4ZSaVfIEjP5zw1omWa/gklq0ltCzUzRJtvMd
icN3k48kael42ANrxdXKKKmt2TUcQwydy1V6ivkeTXbhw2ECOun65SjZyRNZrz2eEo/UOwOzMndB
k0BUrGEYErAE3KYB4PqwBXzHLdpOQ/kbrD5jYiiU04rEe3LCf2SClvjK5ZOr+ludA1aSFfExt0KX
6MnZRqz8Ez9buIeHXTvZjEXwibj7EJPhIr0ZGBcMXSmSIMEDYui/K1dIuLCGPldLIlq9FTump8Jv
Hs7JIjbjwpTM5O8l/IBS7LRS8Qbdw0djRJaaWsqZqhb9HWZI9duI9yZMu9hC+NpQCaa+uE5vpT0w
VsMApWmU2Y4gjGNrfdDTvnEy5DEsf7umTB5pNwvBtKCz7Ya/XHi5EhdICYJp0BPeElr2Z4tHcsWj
h3sdYv5lvz24sxhMYQGqj/6+Ck0WRVz7/XBIt0mmXCl+Z/EqCVbhcc9KuFYAVYZFGHxPxCM48FD+
7OJ0nze3wQs5ynLh3HuPXgU82B4arcbenrpDjowDnq03cq6mc9quVh/4wxxm/VHcid8G3m9bZp3+
9xT2LrlzeNUJgo7EzG4KV6IhG1CVjs1UlozZsnW+HgTp1VoLdxfi7/RK9XSYv1txM45yiJ0mO0Zx
74q5dOzat/snMajGUct/YV3gIdWT14XC4U1+wQe7mqz01kdd1lVytgTBPxxekqaYrj0CQ1ed+rMo
nyF54nBNi0VTcU8WNeKFS3FfeHXdmnu57T0noG5JwOJuInLL+zRiAq5GWE3UNv2oGCX6t9FgNLFb
77NiDIzozkrfYgkvzPCOQxj80uZpzPh3IuCV/nXTgU9RkYD/wsSnUomNoXejs5z/1rNVkKpXCDAO
nONIIHaEErHVEH00watW+/6ZV+zEXaTuk/7s75PRJvbjRQ+kFtmk2QJBh7qvg+6GfSTgSZXtvQmZ
VaYfbpyAYIv8Qby6behaw8Dgu/FPIhYZvde+tqECyFjDqxJjyqlWZ/VKeNn0JFuVVWVHSLiZwpnu
A8OkdhZ8nNR4OQhIlJt44z/WoGWB+JutLmbnW50tyiulFhgL8ExjPrEQMKGQ5JRbzPQBPWnKFJfG
hJcAD284EuSC3EEbb6sCUQBkB/REGMgbLJtuOA4LCp9xldiBq4RUKUKOBzNGQEadZEDQRStFj5lw
dc4gKmDZQvZ5zbFJVhhoUYlsh6nWJW+swj8o4K7gHq4NJbIyMRoqKxM4+6QVLC4MzeQZZpW/yU0D
1DZx5EKcpeaobi1riQXlvpkD38gFv9KSFBmHeGiM41AOyGcyPOOewfL1FI/JpHg2xXM6W6nmppov
4vAI/JhK05JGsVdgahHspuWRVUvmDWgd75hQD7dE/HgQ2+sLAc/viMyL1FdBNYtUIXd3POEp97br
/PnM4JTcIhtCY63ujPJGgoxvxJNVCmoCxAsLab8QsN4OcltY9vTX7wol7/B8KlnH/y7gcGryqLvl
1vEumP3C6SR6DsAo8p1TlMwvXdNN7dZxZ3FzDjKgda7ooHvlNkVLNnjfPtSVRHFxV32hMbTZF82f
ZS+WqIGAOQ0dhterwWyyqvwtYLfSb75AXM7KVvttkU3HRZhqblMSLxb+RsMqQjxr3coWuAMJsV5X
BsLhAUXzxI9ya4AHpmfR36ig2u8bSqASKV3fVKUT5ea65X1rpXNxG7ac+4IKspQR+GYpvzvBj5th
s4YOS3W9YR7Nsoi1ASglq8r0HvUxtkckatY2jwXFMtqjFQ68newwT9M+EILQGXMGj8w6jUjpKBrl
ugXZUOph8VMI7nVtiBDFp+wWlSCx5FgWNmbnh9lPu6P7mGUsNqssKQ5YNrAPvzZVcESJ2mvA2gn4
GCh4gW+qJ7WdjWDRyAmB6VZ5rI52YCsV7yTWO1OtC9Q1g0WFE98d8n1U2mIMtgwn9RzDKUg2HWwS
ZPspNHMI7mjObEMGG2iPOfLADd5FkwPMlQKOWBQjqim3bCOD6EKJSLS65hKo9i/D2F2v1i05ocsb
3dfFty0eGJIv8qhvdHQxTEfFre4Q7tiyUXtUefPZSqfUst2p1aDYWJYazmZO1/IPphVeyNepyICW
bNgeYudSdli1v+eUA8je9pzM/0GJm6cW3JTZdsoKUP7fEj4DjB44DZatGrdxmmvRVYtB+iodyMjU
fKCMqcSgmtrf3tK3ZKIksBldExRz40VnXckoSKgM46IihxdyLCDTwPTOC7rjzmKByUwaKKAmSu8g
mU5OpdCI58YvhImUz2cDlQyeULeY7OJe8r8Kg8xGw22z7sUon2LIOuD13HgrFRfiGoMjZ35xwO4d
zCsZd/fSeGRS7YW9q+cox/StiKbHt12lvLfy/xM4Vb5aRZqDoLCfGB8VEqUZBFqDW+uyvIdrzQc1
lmATuw/aEBvBmeRU5favurgEGF1my+RwTMTD2lw3Wypvjc6boOUO4YhaTmo/YeowZJ9vTwJSxOz0
L226vg+Q7IiXSNGhNmsIIlFPBeAfZlbakaB7zE0+Ino/Bq96x3Hqzz7UosVmpgAxO3//qykNfF74
7bXZM2B0jda+MFqmaP1qheG1h8FyYWxYFI3klwwbMZFt8dtEZR+yiYdv3WQdcb96IvvNdaxNikfC
/fXyP40kSHJjy5hCQBkRyNr4FYN78xpGnS7bmhYPo3pQBuxnAmgFlnbo5kr+53CrYJmNXXdVshhg
FTSV4OOUVj6+cQeGM0KPCrRdKzPRIx9nxr4BijT6TwjK1WwBD1RUEuI6ilt6ejyfJFXOpGXeOgIj
IjlzwTIWpbTfZ738KqphBCPKc++CKlOjMKVKLF6ZZa5rEre3PheKjPILEudp6yk8DBTNhKYE48UY
/NBV8fsM/nc0UfxQYXHwSOrxkHBk0PBEHL6mfhEaXCcTFaVX/XbCcIxf2WPbsxWb8IizXkj1j3gv
8lo2mKELZqMqKGQNweLN6MFwzzPjyRS3ZNhipaImrD+w5aRtndMHNDp8gy4EBK/q3cnFThCUEZXJ
JfjWmJaK92Xvzsv8LBHFWr0XR22ty38JXaXIUV7slnaqkHoROTpRFhkSKnsrN1N3FQHtSekLSdcn
Jc8uXqfhrxdEXs5uY41h0koVkWlwEbbMc0NGOM15bBB3FGFNrwkdQfF4oOAt6oI1MuOY/QJqsr61
PS3y5r3l/4bxWzN/hJENm/p2z88fdu3wXwlD/lQx8jazXkg0wM4kAjIRvMbDEeviK9dqvajGg9Az
D7/nGETPJZPAH/G3qUUOTmyNidO+QHKa6UgYtQsickjXc5pQQzzwJ03RT5ysfPcO7qakxGku+XDu
xW8PtFrUznf+S5ongvuMmU7S8wQnubURzBlmB8QteAP2PICsoRchyP+fMXNuN8DtNbqwzlVuDxop
/HgjDuMLjGWzALm0sXpMFf554Parz24sod/2uHpchmsQmcIT6MlU/jHh7Sr+Kf6ab4P26ShjmcRg
komuQUeF0jfzaIlPbceMS1XXaWR6gE6wLaxW6ZyyBsyA0Le3cfxNzfkjTZaFx8rzJFxThHlvld2A
AGOsnWpLZAWSMk49wvu+Y3jlY75h66YzrwGlLneOz55FxV9sig9mc83/zE6gmKoDRsM+61qQ2sZM
Uz2TtZevLmbztVpWH5DEOXThvDqG3naDOhIefYzOWYFGZXUGveZwv35mHTSuAeFY+wd1dphU1jn2
t1lWNTq+VmLN30Pq/8S4ylmcLKtHH5GUF6WkCemof0NOzLTnOI1Mewlm4a3skyYOMfGtg9dcx+lD
DIf2SQBZVU1DFAVgqDxlDdGsVvSrdgDjwyrFCms1KmfZEtX8+0O4Re45lnAgNoH1E20Pu3xGUe+Y
gw0J7hgBQklA4nWLuq+dKGxMz4vaKzUmH6sOP3USAJ9E4xY8iEISnHWh10IgftICkGeNmgMx/3fX
bvnfRSMnycJDZeMvn4IfoAMAxoc167pudth8fGgJBvLdt1NISdWybxCee4zOr27Et+KTBWHH/5Jl
RkxNwMeoy0ldrD7PXGlcBs5LeqSRQ4fOypxD4vRODJ1ef5z6d3fPKwiIHDbBSUDjrj6cRp0njQ5j
LviYl416H5olZppP8pHSRpZcYEQoMa7H0z0dL7HYD9TZ4ykcNMHM07D+93dBM6IIA0f5mWyFk/xQ
dKwkyvTr9s+rZcDFbPhDtON+h1EF9CfLN1t7VImOf11rXcgKOHfHtUf+9xSRil4lkyVvpI9W+Em6
HjolMOPLxZNRHrZvWcRV1MQRajSuy3IOAa/Gm21JBUQkxz7BpBmWfivWxCe1BzBtGxZn+H+Hzr25
Os6K6QIJxU5t05KRV/BNQLE1kW+YNbpD4AeecON+MeFFi+7pST1hmhyp6hT9pNPLBJ7cVMXlT0l/
wVWZJYxHf5ZjTbIEP8qCsi1VyG7KtgPzyCpo2HzOJaNS6V4a603mE4wzVh8CFUFc055rJjmnN+a4
W6vs6YSBpBggsa6rIvVChgfaBwh9DG1ch8sr/e41GMQy2biJAHpXQa0wsvdy7pp3Ci2R7iaZcxML
sdRQ/cMOEDpBR2gaLVbSJNiEn+l5yvXSMeIIxHVROn55lzbSj9QZRgzhF0W4MMXlZ1nqW5MLviLk
BR/5DDFx5oK4i18r7pZuosUQ+I/Z/2+RERq20j9o7b65S/jlEUCSz/DpbEl3m0e7RYIfj0FTyG7I
qKo971SBtaMKJqPloAqVdDb4XS4zMcfK4sDPMy5qreLbDkzMOq6rRly7ObyGw82+uBMa+U/zotEb
sW8ySDJzJu0ulBHJgtJSS+AN7+PqyKDcx9eQLg35k6FZAWXCtrOxLAvXeSSQ/AlMjL3xZnVkggvd
nQQvuFyLSVd5hfotPPhk8OklnAjzI0ND5Fe77FLdgC3lmfr2ddPfCiBkVXS4M1rgXqwSPnKwQl8i
Nq/0BYzgHLtokViOgKwnzyKIz/pKOot3Pjy3HFJJep0cMIrLNFuY3Ot02O1Un2IxaKs+MaS3WZ2V
3kKpJP0WwG6PIuGvtaqxFmbCZ+PHBeNU/kC687808fTt8VelAP01DONpcFIDze22BnclcbFhBHu+
96lozDD7/GGjFm8lDs7nrQ2cxgqdc0E8WDk/uwH8ODWaKTf7F/V/Ow8b8JysMp22xIUb07JMcS4R
Yie3k8eT6OQ9KZ7zu7xgJqPBE0LwtQP88KjKabmqEeqv5BAoyWbyRVFVwkNYonfoF1+ebiEk3EhZ
jCxxC4PkuJfkk9qjpvGEHPA0mHlwHH3SNV+UVbP/avVRB6HD5ITisqE7OpxBqmFgubPRo95yybL1
uet58Xct+AFPOSsh7d8a1Zxv65cKcp+itTrMP3Es2aLwGT7/Wr8DVfBqaMRf/Ws37crw79xk5Aur
LU+CHLRMFGCc207xaul9Un4tVDsZM/4pCOHIr45md1jXpYlsQJGSaGmM6NbgEcCzDsaM/Jg8sqhs
U6f9415JMpW+XPNsijYoIKd9GBBo+/X5E7P5yY6Nk4x017XsDCgmJlgZ6gWG6rfPhkdiBs7qY8vo
O34PoxDnTJFYZZLt4vd0ycuPHLa4cdegMlK/u1B51V3Ho69OA1InructJu73K6aekwDaEKjnLi78
nOlWMTx7LyJIA9Ns41ELfONz2NKVThY3GrHwJMvZd2MZMRgsHF0xwAg1nYuSpQnT/iU6BiISJpGa
/x16ZIPH15WVPaTGAWg12Db8BaPBrvU3usJXTIWDXGEERx8FZ88B8qz6mFOyOksTRPUWOlJPLMyF
ENYUYK1NORH86qZjwsddVd7EG3AtCJTh88dfq3QbbH1WUrPvItJCHC5Kc6dUVoQ+3EgrOC6mouA8
mu5OejUN7PGC6AyexDjPFTiwX/GbIEcsgIb5RFFvmjc6VQ6zQ7BhD8LbfVCoE9VYhrLq1ijeTAc1
3QkHamhX62K2KzsP33hrTu/tWcHWSxnRSvb4DwRUEaID++R9Eg41oC6LzDbs/TY4DZyK/eGg0oUO
SN9CiusueFmVNQ+Q4HfIwizoU66C74QS6bSM/+fqpj4puWTgzcGm4eTL1lF+AojuAtZnG4Hb2zlh
508B6//rsE+fDAtjeES8QeLzrFOWObTN9yL/guRCI/Gjdi2Bvy65aQ4NB1zSP54u16d3nGD9rwRt
BEqyVLSc1Zw/HWkOvxcEanWxUG79z+LNQov0tq5XvIIjvL8OgyebpmODSGezgR5m/Xfvremvd1YU
tja5GkZAHq283By7fy3b66h7n/jgUu5d72U+sK9ndgjjfH7nsds9w9LUJNktpyS3o6pJfFqI8VUM
qSrCwkPXmFZuEUo7j0lsZ2bXhqZaaprdxHEV4hjyrZJxlxX4ph/AbRMSenhK1z0lPBCKTClTQcWa
wLm3CqxcqhjmNQOxhv+mCeFOX1xw6snUwutN92t55mmCVTMi4FYJqU/lx2SkWgVsbd3IdXTdpHey
9vN5MMz5VR8IPtEby4iv3WtHMV6TDItsrBVAgWBlFM5k7rSMaA2z77XPqXwGERhMcQwC7tul2W3K
skT0anmM722BTpN/tlKZp4PjOyFflAzSxGs+RMtmDCoEGbO+9AP2EF42D0sEn5P6XGRRfsoKpPuE
aAKjkJzp5NZjXlsgH8y519olNO9Ca9il8sOATuVDoaiQALhpoOgreQAj6YibEtRFl7fE2aOgo8Kw
4xoeU2eOUh+NXrt/IukoLsQh5RoRjA5oxQtnY8bJxoe3lnNBUqf3FgFeUoqo1FY4NuDHi5gw0IAV
Pknd4zpJjir09E3DSJTXCBnYOLnRa2xY/M+qv14/qkHjiY6ssWkViAZGtFzWffrICs6M8DnbxE+0
cH+VqmLoaJ5CUYmIWsiS4Mt4zyuRYVOUi1AJxMsVLI9vTWF+vYvTQTyFWslcVbTtYHQCcCAYHW8h
gfwS009VOybfMPTV7SgQ206K+COVOKsKICDCE48h+IYQl7kRnjnjwLOdNjd3hlSQstRrmi3lnegh
Eo8xDhuTZeoWds6JRECUG5R4pGpxfGwAAkX7atFJRK1OeAKFHNj2kuKVwW+lIBxQcLbKPB1nFgVo
AGzcP+LSf8obd/sqajXUE+5YuBq+BQdAVT12Ro/kRGCHWqwDogt7Bm2V4LcF/D7jWB0d1ktX0JkZ
H5npsV+32wL2vv36HTTr1vE3IQDSg+Nq3DtylSDQDsV7lfNlF0kRt3AXRZKQFhCceCZ2LM0Ia4Gr
cvoxPb9xYmDC3A/45liHiyikbiP0nYWchPEWKFxx5rqOVaJccHOXI47eizz1fVD+kXOPwi64K0Jq
TcrO8GGcg7VqOwkQJY0VXWTTrUXW70ZNRo0soWz6hgwyYoCHqafYTwnB3wZa02dzuDjkeD3sVaCd
GVhi1jkOBCLG39Q2YSC6zi8vaAu5LQ+3IqO1yVOm0JocNUMcADn9w2OdWjTme7k8G2RhiRbekXRe
QMlf1M5kNF+QxLrckQJiq18bxvtbdNObmGeHptX3PnM1pYHbqXEFEqRTH87jDlZydl4hWs44RKW4
H9giPjzrtJCdQk4XWqtN/oaKjuqgcIF03B7kLPV67tf9dUUo1eu9eB2qQr+nrlUyIrHDd0+yiuwt
Tpkv6je/xnx4cTdm/v13oi7gn+pI5B0SKBvmcF6M2p/8ZVT93LrzFcocx6jWVhf+N+mCyrJhp07h
3t45l9n5kNqSC312n3CcgNLTgdsC++7ZSDAfmAXBeCfRJ5TS4loW91ShHGt8iQqV9Kuj9rxZK1Mg
2Rw/6PFDzEQmW7XowGMPKbXqhsPoHeb1qnfg3U8qbcAhx4riWbosC32yrp6q5cNP7qxs7V2GXPLe
dT5Xri9gIAysD5CYsrOdMrroS/E3xFZk5OIw7yD3HoC3E+a0nZqlE+lJ9o9mp/6csfZz/QK7QKp2
Ve0w0aTPqS4VtiaCHQy+Q3bkIwaCli2VJAn096aYxHlup5Bo7bsojcjtPEvmin8puPReuPRZCypo
eg1ccVkXiM8G7OvkxWjGILoGTnuJ5FLGL2er1+1NXufe655GBMUbgUTbVpMzTi7pzkskaSIn/NY+
dHhI0VHoX5B3w1UYMOTmohxgi7d/Xnvr4Uyhk17XrCGI1lhGwtLXcNVn8DuvuG/BW4igET3AFh2X
WASS/QjR9wVFg3qakWKvxaoupDnAbTC8/vCp0NThnnRMcrUGoZ6XbXqAs/UgbppindPi8GVkz05i
5rJuFj4cV6ZA/RRvJyQA9eVmEuz3nomCCqRBfMrHD7YoSs0ucTTh/ct7/b6hmCtAiKUySXNbtyFY
tWzDI9NuPuqp8HQtqTQwHB9mEJ1ke3yQ9xhziJeJd8Te9UxnxnEE29AvoBZTAmI7lruiq/0hcx2L
OUbxNrEr8PqbkxYlwN/WFZB6Q2wxngodliensAbH6GAnGEjoQC2GsgRWFVode/eOaEWvu4+Owmmj
GzDw9bF2NKOBuXeFa++uXh3dYeannnxCqLoobLy/sgfwqBKLMBwDv0R1R+fUqKw3c9nU5Nc5+idY
KYvOmQ7cw2DcFvb9mND/sbNN80brEJmT1WXaiOzfoOm9JxnuQO8iabiyAKQT9IRT+ILJe3V8Ow2+
J9saGwSQn3jjdbK7WqCX/qp8sa5tEnBWjgGMZ0SqPo/YtiJQrIs4PSBJMMCNEKKtD9gSI6FgCnuN
+BRnkBNkbudn+ryLl0F+Ma/a/IBxt9CjfCRm3GiphkA7TM4tGhKPwR6ut1beMQ+5MZQg8tAorSlV
0XNC7OUEFO2CoVs/MoEgWvfSlcmNo4ki3LKglCDPKeNaPzFFta5eLguXDp9J4ImeYr8R3QpcJSUR
BfwQRUXAHpsoc7GOFtREbgSQUkKjhAHqjNJZZLfX+f/3gVuls0xZ3hR5VVzEckBk3AXKwieKntCF
FCp02xMpV8xEzgI6+9kXnl4UPPz9nw0ayN3+zFTeEWWqF7e3rTv5z3blwz6SHESymjaOnARGlFEU
cdAY2b93W1dXccieVUZPg+HHwgGbJeHlZNGVdDq/8FwqfGEQKvNOzA8DG8+nGxYMnFyu4T7Pt8W+
GZE8XxrlWRnePa6T9ahcxjlOgef9JvZ3u/qaPgq9Iw948e8j6QGWA8hIjsovUzKXqtuu4lc/hbud
HNBZN95Zl+ce0QEPELVskb+aqwBgGn2PccBMGBSAnG3YMwah3pM7pRYRULeMiQb4CnI+tgXlhmN2
d/aJOfYXzKzxjIJry/QmMFboqcKK9rk36YCopnIw9N35goEYOrv+emNuIHdqtuo0KZV/tirXvUQw
v76Sm4IFE5wDTWh83PkxNLufbd08RlhZ/8vF8CdaVqsHmLiwu74qL+pplOt5S+5nXdluL90A/Uva
SZNAlIQOj+53OawojTHAORMaPv6kyil5qfFKRsM7QYKRJzc6oLqgOUMCAt8bFCWhCtLE7DlmzgyE
ki85v61+loA7/5gcHymG4MP+m8sU5s0obfWFx4bDg+c36qVwb90kPGG9mc3NXc4qbq5YXsYZGDwt
4awy6Q1PnRzjzN0ubgD/BkE7c7202IdEZdv2R9a80uAkynxpbxU/U+ayrwTBP0caOrfju+N6Kwto
pgUuzqTUnKqy5JTJec6eDBnp0HxSH/CX25n6yPXCra6ALuB+pYXMIH2n4B04AJFagPsJxAtNsbG3
dOUsxfOCtXXJt/GA0B/X/6nupsIx7usGMnCbNPSZOnyR/pmGZMtdzvz5e2s+rP0qkpB2ucBAbGFV
P+0TDGvpmOF5oFDdMsMcgvxNv5tv9uYWwXyeCyzs9RfKatS1M2E1v0dhhJVSXod/qRbYqf0DW6Nl
PvjgE9o+aY3+pdPExD4QmIVrgtHBFOCSywk7kSAA/gRk8xN2ycvE5vNAI24ne1UNLmLg3/4Z+9Aj
pKT0/MnEn9mVMTq7US0/RauTOCNWeED17nRtHX5KtKRXdAO7UGszSHYEOvfqV3m9UkZSSBSAFzJv
mU8BbHVhoxazWOaZoDvzjwXwOE56QfxloNHzJySwSNlbvAZ/TAyX5BAfJo+kPENbZovC1Y/PycsM
7DmwbYuVNEH0UpQoa9ikR5J/zw5f8I9aC8tqPfs0r+kIBB0sV6qDI2tvXnBfWDyofsstPRb18ZPk
Ncbu2QjFBUPKaHr6Fw7rUD1HTvZSWimZkHuqTi83C/8MPUvC/hYTQxfNifL2lrDmlOohk1NN4xzO
k1zX3FyFsNu4HF4mEhwzsAvYmJGaOwwBQyV03xrTpakzKNySADHPjWU94WA6+tFugfg/dxWO679O
1LNfMoYdtwm06MEBdEUD4kRPS9DlGvdY/K+sQY30kc1qxrzw8lWwnFFnp6HIextqCxBXVDpepiQ5
1XdDuxKfRZ1jTjWZ8EuNQMQ/TuZ6W+wYlY5LTKfBBWqsqAJ8HI66OQaLCreEkzP7XrwmkTesQNFx
anJJ5A6Cu/oAn8NDOj6cPMykDkv84klAqEUKm6R2x9S0OLV/1l0zzXdOwoB0wX8OcRxJnPgpTp9s
/+fXUedYSdGeCt4rzhgF8Zt1OnqR53PIZSxrOkyycofv3fYwQJvl0SXqoXU7aTg5+ignZpIMI7II
FNbWKBqOyoMCwxgzUJZDz4uwtWQk7FJ1uSGFVXqmTMgEV1Gj2CulkqxWAbzEnVkVTeOzbfiLYm/A
MOA589w3NsVaAozo7x3T/xGiCl1AhFv9Bx/3rO8t91H4BMM+eF/o34gOnVtM1xxKk/XIQwqX/nvG
scjoxEx5K5FLVEhpm6N665Rhn1MFmpxNtieAKGojKomEopqLIOgXyjU2y7KAz+vsRVJWC2fpNHQ9
Hwo4BpjbCTeOvw5exmp7TlRZhRmLeFML5aGxT5y1f8TYVNMf/++lyKwNNlf4ocX4/ksAmtaCgpXU
WxXkekAr+7o2/d6XnGg5UnkiqYxT4LXVrd9Juir13DZNyc346TIWFD/47MwcpFwVFIsQxxfg1PY5
oc/z2I3/cdPK24iFlWfAVS1kC9QNYn50E/KCOpIYACFvfHy7imLmshlVomZY8iW0nmywP7adl3e1
xtqFeskd6Eeiyj1IXiEliaFN0YE6OOPlj2McEkRZMOt1M3KOrm7jwpd5GidSeI5urjtm/6RW/WCR
rd9g8sXFKZvLZkQFmjb42M1+LxtrNFD61YIG0xXPPYcPkHYZtGZ73in6EbBoLZ/ZBwztZIfV1Vwo
RTX8ois3Sik35nT/phTc9lkPPqckkMOL3Y7I3d/2IFPyuST90OPsNXevf89t5Zg8Lx0tfCgWusaG
XWzvkMk8eNMfMXWUoeXqnfE9/c9hzxmLJgcqyS/L1mmmN/3d6eVPd5JB0IgZufAOL6y48JWlHjQA
YRsVUu/tqqDFrUNVSdowieBys0VWcfwSDwSEkU3OjDhy1gQEIaO5/S4DG7WKOC7liaIOPWa5gAyV
cFGj8Nnl5m9DXarr0I8WZ/iHyZHblhVPxBRWrFK3k0hZEf75eVb3PgMZpzCodJPk8+x8ZvqaTKK6
IfAlh+Pwp+p8rwfpuBlGDrsHvzBp5ghVqVLgSoutbStd+y7SJOjQPKmeB7idJlwPyHgQI5Nn4isb
11wohcRx5QrRhJBdNtYgsp1VFFtuzXRGW20hIyaSFJIk39Ot+oGluBoQ0pj5Ul9MNFyXIe8Ys5kR
dlVM7dNlAyTdmNurDX+oHPMMOsf8Ji18XLPoJL3oyAmgmCORDjf8/dcG0K9x7IT7lr95gIyJa7Xa
6Jb+iEvfb2Cm2xzrLmFzTPjp6DqMVwI6Ap4iYR2ibAGFHJmmDpuaZkwWv46P7tj+VeJyd9GI4evs
bhawFIbR/pNU1iTLUr0SclioXbJTSTNPIIMVOBV3+CuJE0rf7nd4pIBsNbwKUmBWOF4EnpNphjC/
UqR2cE3+9uhcb3Ji+oMOy12qDvnueU1dW13vo4IReeae/20WGmFJGa4GgrMSGDI50oBc/KqZDuF8
b6cMEhnk4WvBLwf3dUobuppL3lrVD0/5Mf4gWhwXFM1WQdzG0GHuK6l3piT9f3uIjORTMd20uX8J
3/ra/xjOrykaHXnDJykCljZcO3FtAxA5IobgNFG5jgAVcSLCpa8tiQdL8pRpXLYaLU6CUOZev+Q+
5/4/Cy6ZrJVHJ1dWoi6bsq7kztiHbkO24Q1fbkGjjt3G2gnMzUTrtXo/BItXf/eEqB0cbToSMpH+
/HLLSi8Y25kECDlp2bqRzsXg0x5O9QHqAB3ZDiNGyic4YDVq2i+acjiPe4rsevZpY4cPR4Wy55+N
qj77XB5f6pykfbi7fe3VSZXaJJFah7Vu+6xW4H2PgWcNIX+xih5HVngg8ujc9gMmRrKGg/slX5UR
jQvO+u6LM0iljTNUOi2Q2HCIVTtqFjNcQr7l/FV9r8JCtqRH0KcsmMjai+ibrSJgWoFDNI8G83kk
7z5K30TNp1fi3M+9CJmOLSATkh7pYP0Sc6Fr63dCMvCP3TznxLl5WdbVtMk+BdNglEh2lfi26vx1
nSfsbkplydCr+59Jjc3J8E65Z19EO9vY+8uGHA/UndWfgoz+Vj5Ii0t9Eh3YhWrYPFmcU+iJ9Nnq
PxP8NhROi+sAyHYqgzNy51nOcjVHuKDV9W15WwoTXM2OtrRkq6ajpkQOEFb1EnU63sRJA9sR49C2
R6ztApeihdHaAd6/tTEXuZgiN/elNOTrPbQso0nr9edUqapF+4pa839U/pfGhiR37/qzWT/ibo5A
JD3ThmRD7r+De77ynqDqEb0cyRoWP1TWOgAUK5LDDdvlWejF3nKPLn6gC3SFCCdFwLEAQLdbTxxD
b+PWkGA4iJFYOhWGO55MFP4+yl3y/I64shmRmGhZFhrFRXfrWB0ZJoM1DbC6rZsicAqOLAWml9XC
K8ByDPM3hiZ1P8+iYA/1qaA4GmO1XYyXMNCog8tdlRyJPzhTr8oTvJzgRdhk6RQBT5sQz+43PqYK
bILBYoj7QGZoQpnBqRPevJRUVbqyKIjWhZ11D1QBnDUzLgD2T5GjMDgUb9LAq4fgoONNXcfPqHLa
m/gmWoXUaPrWDREzyFU0EWpZ/8LRzHHRL7iakTcRwV9ymV1xThNFM4qB5BTl17GuHfqk6zU7HU6X
1OK0lIYT8TiFeOKdubTs+HzE677tvGMu6ty7tA3vYunPVEXWH+gDE9qqwweqmDLuyjIPN1zWt7gd
Ow18wEKgEShhtVmzWNKpCGumQSMHJ5bkSNfF65RxJh3FxP5Hl55SdqzrHs9cQlu/9sc9aSmIP5cU
mxukrB7eBw79JWb8PCmNXHbwNVzWf6+700J1YWNC8oe5KGnwYTHQUOHjOHxEZhb6oF/TZogTcOWc
BvAyk9/Ost6QJ8ZZfuTtU6/TqVMbHrKUoZvTkslvjMhelgZD0WvSL0M9FnzAIiJ54yi+AWF+RNH6
dvLUX2FtjkkTBQ1xO6x3nwzE+0MXd8HJdgbLdmVe0nzBlOjb3RNPprdtzaxDFqe9YLbIH+vIgaGb
AQP+gZqsB2yDeDE9/9hwwkFJvG+EURMJD2XvrOCxGfelimBI4xVFc/lqzl9PifC6ylT1uIdYW+oX
9tfOzpLirGSyidB1BOVIJ1ZFchYZ940/qUOJIRlY61dXWgmoGU0nf4zMV+mN31fjr2NtRkz6l1iP
Yp8Qpr20IDjGYS2M8upNPujmkNn0EbsXczckFJ9nZZeKcFAlhPt90Z/JgNiKpFJAbaEzOU3eV5nI
4fmnqv5KX6w1i1fPE1iiOMAC9id9q5TRyTOMvNhK9iGdrHhTVsRk5MLczQ85EN2T6+3ZWmYge9wg
tv7rmhIoPw+JT6uG9GTXudgqWwF/KTUgrWU8xsAjeCpoiXkdlJTMhAMt6rDSOS1lbAM/qfE588K0
b0KE6q9E2ESg8yeK9xb9moqLrcfhxRDxLTknMJk8ImUgWCzsodZvgffVMSPdc5MJVxzrwaE8Wu+p
v7pcW6A8h5w8MmtfIPy2VrhwKJG3RliZPnIA01CJ7l0kuJSdwWoMyaV6yg0DO3PiuvAOQ/jD2n2S
TLznIEMxnZdXlZPW5OJXFIhWFpcG/B00wiJ+8HKTp3VOr2KHqdmwe26rUshrNM3/VojQeZpph1IZ
kc2Rgwvm2eXL0taqnFNiFauFQHUuT6tGe2vr1U4U7U9j5nFX9WkVBAyxk1GebAZ9OVvs6KrybOnj
q8REoltV1/34xX6D3jNXyqSrSOv7P0Oant6oFVjFODo0m3nxpjvxhDv9F91bEPpmg3MgnRKiBZFb
StUzETvvggZakVL/bIiT2mm1Gw4/zh+OHaFpzo/Lg5SxZZD9RrBGlxEnJaBjWsxryWYWw6WRSf5L
2yCvdwWhPIiJip7xApXSukF+cou1fiJqa1CTjYybd8vX/VV4aIdoZ8fh71MIS6L3X5v4k6i4oKCO
SM2UacgOJuZfMd9NBokTpZAsThJRYYmlLwwK8ueqS+ETq5hzVlPWQicx7zN9nfL0fx0AGss/4j8z
oYU3thqntvLv/RPiRoXTLVSRCXD/QKcPAVeWcGYodUe31nij7wDtArs7p6e/EC5IBDPe2hZwvGSO
6BGSoIy/WB47hm3Bm5KiMlyLCs5x3Y9L95fC5Vwn5cpGXqpnrR7VwUuCveUw0JI5GVE+ziEI4Zm/
gCIPil97LvNdlxHRJKps4jxO33pDytSxMOF+D6YcgsySwZaUzDBrUqHEbQE3S1BD0qr9Vdck9olh
o9K0byfTJ0mEUyvmYAAx3wcT5WRoFc6ScS9H7VKi9rfLaHkr7RDGF2wHERZgocY2aoNkRBZT9Mhh
wfR+m9UiYZzAIMBDP4MN4m03j1O4vTfNJA5upbAO++6vJRK3IXYspruNf1556r2uU4pJJVHixo1n
YuMEnTnjWLz+6JejHraCyYaCu6AIDB1hafBlOq0OMljXgr1QK+anjIckeuqRsefyRP+90a1j5zf9
tIMTIfZwLaURZTMg3qMoLMYD+h+vAM14uoo7mU60jMC9ImnWSm7B39YhkzaBnbXe9pAX7sguQ9cw
fBMAwxiN6xE/zWmYS1C337g2ey0Zv6orrtgfJmmYl0l5TtYn02HIzHiVA8OdgnHCQodfYXP4l5Ap
6i6oyFdU9h8CkyaV4zGZnWXrjUGK3aSFJ2IcpZ9fVkmStv51dhQ97qQi8RCCTtjIzJGarr0ISvKo
BO/pxib6mzAiXSYTgtRI3+WjJHuGyEZCoyaOLXFs64Uz1irtQR22ki7o3GZ5KzT4tp8Lu5t2obeJ
pED21gTe60qur5n5+RqoUbelNwWZNXUX2/MqHAtMPzHmVD2GQ4rn5G2HI47ta9Z+uEpNIFTeo8QR
yhwu6rW4h78kpIPIPnYKJhhB3GYqIDQ1F6ZzHzaVzbUhC9tqmXkCHMUHNoMPp3C058mmA62W4IOd
900nmnIYgFqxKkZwl0IluPwx8fOOql9trYhGcQfGgPNQNJPiSm2vqKWrh2Z6PuQqZjnCnPEZDYrN
N3xAe8DFLXhku72knoMYSWkpShqwkZp7COMRKGtiWSVAPtHcKtaHftqgfy+WByZKqUJzJzYBfYta
pPGdVbfXeVKPb3FkvGUfUKmSNZZcJ0htqlI1U/vKdddFJELXcDSC7PAetJ79aD7sjr8gcJBWAC+d
bT+izlXQ5p/vHa6t+EHU7TBMaHMzxirnz88QPcZ6OOzV/hmLBiYf7sDY78Fc+TB9S4Fqjde5Ca+A
kDzFsvrmc37OKpR5PhGegJs27fJZfeUSA6l6WXO0f8jo0yFkBYmEzrbj/sifJx0IbI1HN2NBxjN6
+VhM/dA0Nr1ezsNocpNVVFOy9oOxMCWX6seJtRCcjLkVmat4SgG34gQWNdm2okMzTrLh/vBGIpuD
MjZSOQVlk+We2s/DamgUHSCDzy6SQpP/I3kGw0qiFZR1JhLB7FJ9E97nwDt5P04u7Fi9sLjvXPEI
hpgJBH4qzfg7aX4RN/7g/nVU5zbf/TTrOgqK9PEUFy6H1WxUORHYtgGkXDIcB3Y9WUKFt7KBXgzn
roEAkkFD4BBQ+5RdfEBcE7ycn8evZpbBfAkn6K2vtS9wJcMOm6mXaJaXaXV4fU6yuAGn8Xc/njRN
rgonS11112wryJs6vHRKzCdElILduVYkDbSrrDJ8jp50xDyQrNWQjLGM37qzsFbD5wbElOCXjE2M
m86MVppFaR1IKtVJ+GYZj1SCPcZNmoGudoTdcTc2g3pJvPx+lQULeAMfAKA0UjZSlJK7GEsbThgu
FKf6px0Vejebm1PnUBO9fioC8atLYRgqZXzzHVlxAXTGJ4uUEDp27poFlzTOwkMvVJ4VPpYa+u4T
2CKuCM/GYB/pDr4NjYXsPtvOF2lDxJB01FuPBO7TRv4QTH+DTByFGqYJ4DKW+Eb7l7Jl4V6C/aRN
6PnAIO3o2JiR+r094UDeIzBHom4jGRlpgn1qTs0iprFQUxf20vHeMlIRAvPbFEWy9BstMLof7KkK
C4EEkX/g85KnV+G5UzlWQ/0t4dTBqOP7ZfEDW1d6go5DeMXEe9RbPywCrSUXq28cDqvOd0ZY4QwC
XhsQU8mqLWHujPDKqTMgEZ+YFriyy1Vs+Om5Twd1I4V1G/5HC1XGSUhqC7f06d3V/Ghqcqm+iaN2
D7bfepJEqGAjgrfKzQyBms7FNZk4qG2kxP2DdNlWZ659gmFzNQhK680bWMrmzfKc14EJW1AwfDFm
3oz7n0oWaiThDk7R9yIj+WTT28ygGxtFzFHh/yBWuJJpsu9YaJnzCVtUOlDY2sh5ejHgYl38M6TG
A9je7vADwO5Z8f+I1eA3S/4PWrMMi4tHQfAUoKajphcdwu/nHw0XAn3FEb4jjpjpHufpqp2zq3pL
XpliFDu1276O5gZfzj9K8eMrx5ofDecH9Eit/Sjd/uA9dywJH9k3YWdgYOKjulaURetG9MwUxeeC
s8PJxV1cLQbvZruuHmKd+Y71zpUtM/HXxUcpxst+SmceF0jSUsDC9TMXlvKNLLbNcAZu+sgrPB2+
MN2NtDgOBP1Y4R/N6U67avPaAud8HkavmFImHyQS2YohToMgpS8zy4JzfEMnh4AvFqWo6EMz/azd
cZoNa4d/ty9C0+5QjSYPy0o8Og2VKzMWk0+NTbOF0/fXKflY33KJq1JJSVkyaiHrsUl1/Q/RG7LK
mjz3yD0hclg4nqiZNmpqi6hWJss0kda18/b6SdkfUJr+frShwBJnt94UbNIXQB2WX0Q9SlmEPZ3A
ZW4IVotTlqjVAG2tmFfimACbE87tuhrki4eUQ+LzGsHUblf3n0YKgsQDlfFzHs579YzxAMrOSrTK
3qnZ+yCQA/E10tR2xkWqb1BUfVYoTJaLWz3oqAOn2DodmNIBA4tO8Jj/qwHvM44opAG3udNBA9Bs
rer4uk33kfURc7FxfqNmHyR9vmcOaKHNnkROXVWHZpgjtkhp/RgNLAr93WI7nw3PY2xdRbjI+nSS
tdW8jl0KL/0mr5gOwUtXTKpISXEgpx/zQJrxsTg57CguWH/XeD6FWkjSAqqVC6P/mhT49ZMB1p//
XwGGcXFWalNGXBrSAOY49XvQHRlGEuvaIMLm6GI6KHEFaHef6jemfZ2PttsrNh+mogzkfXRVz0vb
hwQ+2R1+p7v0jQkbiVAFRK9C9c67W8c3aXvpTf1VWoGmUmrOW/xL0DL0Q9QfhOIRrNBDMr90EAWa
WEsg0CkbihK+CpsKrr10SNoqoeiDRR5kGzXGw76CczGiGhPzZAxQp8yU06FG8jcb2KpKDUctiYRB
4QHiXqZ2vjNnqY5aPABQO4Gt5aEgX6VUC72jv4GBgikZ7BO1LC+vjKFinDJz56eTFPmCWHVNi1fM
6E0hUmLvMahiTWCGvcS6wP9ASDh7U030UvmCFtgQKRLXgkyUyibUgngrsl5RvDAHXQVIersWK9Bm
zuFPa11HY0lcXuSGgb5bG5Dj5ZpWDHWrAoiM2Aj0zoXZeM6ytQkdryr4aGkMFl++p2+lAWQHY4Wo
hR4wHIhK4YitEmjhkSPp+zemoOcEScZdWf5pRO76E7mib4qpdpiTmjVgVnGo9cThjlOKsUVb5/ZR
K8u7BA9Wuh9XNxBjvBHpU7GuZEKyM0CzLz2/N6R2q1d1S06D4DHVmZ6HB5gO4KwmsOubwuP2XkRB
BlKD9pQW3BNjxOgeZ9IDRFjkA6SH9L2mlP8PhE8UpdwOAxsk+4e4rZe80YgmRzqjcUVrUHIqIJ4D
wgKjCl9+njVuodcSVUL8UvMn9zY1Ho/K7M2RnwvZFv7AzzHY8rqWZ7W7HADZIFEioBna35gPUEVH
SxneZMfk0OxmtSZoveSB4dj8FM64J2HxhwjaK0DORvXpBPsLdd3AphuciSdaKJa5Q0PZzVD0kEF+
3hls1vlHn77Gi/QRWw6k1d+u7B5EXN61mdGRfff/TTgh4Ue9+hdFs39HOJ2opvK0BLQ8sE6E6r/0
3j/GocIOKK3q2ZksRr1dDfaUx7CrPHY8oyNOw7lXW2UtG6cae+ERjuBclCrfIJucUn8OWGsGN0hA
0X1bMK/WcUshNNUKlJ1j0Ew+3DeOntHk5lHOfJCtXEQX+7z87j4PqKbxDeBsmgBtNIpvF+JGJpuC
1yo8ZdQm9/3tDW2LlCUqFWHamVIrVv85+o2zw549QrjXmQlWF8tJ/Kl+MZ1kz0sD+vvRT3mK+4vk
X4mNwUgVsextWlKW5nv+3O5Nu5G4rdrHjfCTWX3MHhO1sYUVPWvlveaWJ5Lu0Jpcdy+oOCzx5vWR
0vgi/kcE3C5gwcmXKyfQnQ4uvTZo2ciaX9hW3vhuEsZ0lovpZWDgvmVHEVRzaBslqpjVQVuuIqBM
NHyQhEL0SA/AJQFinsbFnMWO5Dg+aujod2b/ZVKVHAINRv4BiLEa6EQCyPEGvMHwbZHmc7r4kd5o
TNqI0jolb14576d1VW1bsz2tASveSEgpy++z9Tn3hbP9T8MqQGMv1Lzl2q0HleqkLEfihkbSJWBV
1zWG/HMIwfFhZekWQLjHUhpMVgKEJDmdaCLVbFBZc1468tV6FNBXZ+CuKgPafiPi1oMfPhMJqJly
IGiLFxP+M2TMGW6GTw6/yi/GYqmWSs0zk0HJOUfa/5o0q8qAlHt9PV26H+t+BqOPN9Z2g9zBY+vI
r9meTOVGYKUGnwbRVxzQnt+DMq8b87tNyjGhhWZFUvvTHw38Pka52V/kwPE8Vv8n1Bc8cAjYobJz
wRoZz7d3z8EosUfsSE9yftZ9PVDhEEG08PNBgEkpwWk6NUu11dlAOLgRatycRbYPnYErcZ+330lK
itHbGWLa0RYpA9MgtDBqAnfyxKyL5ygGLSRe1qJ3szheYHUJIcPmP26GJq/sAPpAsPlPLKkWKFJM
Y44adZ/2/tIrQ590cI1SL6C6LR71xsbsf+0ictKSpgSS5y7K0BZgYY64cMgRL62y16EvIjhILJ1J
Wh09zPUCtK/Maf/A3rfKwmEgRxm7Bxn+4vU9HNN7Ep2hmZKW4Ls0u+G56q3Xz+ctJAkbigQn8OAj
P1DO7kWIUZhe8prfxQ9HU/EPBVg7KTxgW8NJw+kifGQT/zsupSjtlUxld48ddX2zXmf8t5Y/ZEPH
JgaW1NGkms53ExWxWV599Z02fSNV0PjF1T9NyZZUptTmxqyeecM9IhqZGvLmF9kopc8fNWKxgYWD
Vi9D+0FjKJiNgLAySjYFp5hf1iyboDx4SyhvLaNsFNgmbAKwj80bUFK4A9qnfQ/41RlF0XXwj2NG
JvSOfzFcvw1KE1+lBB4pKAQFpckWbxTZiauaujFSm6bUxDm9IHUB02iWKri/i1lJ2i0/VTs3Y9Ge
faH+Ajl8l2Te2XKAYwunQNoEcDj3p6svkIJ3BFNDEB/HeGzS8Tb0P8QLBE6fWWVtEeUT5br2aYbk
jpExez2PyaszlMYhayo95N8ZVrYbeUkhVbt+R8PxOs5j32IJPzMUuY3ppuItYrVIRH6G5pAsoJAw
jPIkPyRFix18sJU4YXOXXAKPC0I6nOycCNCa65zhnqzcI+bFawLwE/7YR7RZhTkgZYp0UnGt93y3
7wRUAJ7nMBLUT6wVDDLchi9ifQ9Cg8PCZAIeks1wITxQ/e8zQWjvr0IfMWDic4KFKvMd0KsyOOE6
gQurLKTVu3079oq2s6ztsuCsuOrNG2uc08J5gT4UAtT9MVYJt89B/+bOVdPCRTDcFfZBPSRHnvv9
oDbh4/ZPpxGu/h3vd4zyqu/KzzJdkxb+C0fRrPXoBgUsP38jzAba/llazwCevcC4CoXFGm4g7s1k
/UD1xSeMl8lhAIbJhZopNZ06EyPpm9hTnGSI55QMFW/R/iyFms8/JK70vp+DncQJutt1njiwvoDb
krfWkrIBDKK4akh+fPRZMVIWYDEKErGeduCDnUEpfrMGIeaDetzfDbGNsMpclo82ROgPNBCihFY8
Fk9jq1uqo8M4vEcHy3sFVMlO2adKKZ5MEAboxj5OluCdyckrTn6beo6EMZPCRhJHU+jM6+XCiaoQ
4SOc8p5WDkEkkelhHRygqvgd6EDNFUO4jwCE162Y8vO+3J5vrbLpR9SRpFGK6hIKt3WNk9KO9zm5
oi/lLtHjXqfqlPbfUBoTXKNa6huqcGYWUkNNoD4VEo+o382gKDvnwoPNAKiDjZOdfsnCMw0Axcaz
2ES2laZGOU7K/u8m5wqJ4Uyd4Gv1jvkUyixwPOepgsz/VWJWsBDYOOD+MUGkclCdC3KVQ1XQk++y
gYxADFbd4/P5sMklQ7KSKIByTc3Rgs5885Gh736Xckb8y9fsHowkxIytmJiURzLBUXrc9IA2BAgr
zoBcrChjUnev0ZzM0nbTwXPBNrB/jqc+gVBSQDdSrSZaqmloLGLfU3d9T2cYo40y8avrfGxNkGAm
Ifi9NKz3CBaXVkcon9ABhC9vTEM4lfNJKo/VHj3fUIpfzJJ90Xa7AOT7aikRelX6tcUVEhLPrSqM
hzz5BOmB3ZQEXXvmloH0eWB50RVdAY3JpRXQXaR7cpSCzRdQbZnpgESXjT1B632hPpq6Eda2L5ZO
zdE0WRkUh4JbQMzO7kkM/FIB+5pXRor0FJvY4dbDgYRnKbfWc5iPM/yLwnXZt6/6bWiSZaK5vj7C
hrvBPkkDjgpWxGEqfCUL9DRDWaSjTAmnsJYDXi/eEbzfEx9Lklz2jrTZ3fgp3XbWiJXj46udtwwD
Ayr5Aa6VnEZkm+pdSFOEaBkMWzyCWBEtLnWU91vVFOsCeZgCj+nEXTewrmSnlCYIeOarlfxOBvk3
s1mGbSmsjuUDBofWv7KfkOIY+YaEXdHaM8/IWbLqFAgZRBVpBF/ZNPtX3T3/LlRheFSRPxQcikId
YkwgHDpOgIgXIhbkxsWnUVdpNfzzKu/R6eQpaRqRO7MgRThFj9SPWAG54GG7SGs2XUZ5++f+R6YJ
rJG4pPn4mPoDjPOLmbUu2ErCl/zLlX/S3mW0T/6gLupJd923FGm4kzao97iGnDiRNogLihqtIKk3
MiUt/9IDHe+IIoke882Mc13A5Uxg9u2kniD+Mkt2xOA4BbWH2sLvQPTuD5R6qNCochqCpuOpJGz+
l0ekdeskASebKapjWOVimundnO+oko6ZXylrZo7Zj5U+y0KJOSx7A8OSSSjRafZxRtu+UuO48VzE
VEetmPP7ktCWjS3cNCqC4GDFAqHTOoGZjn0iutT1fMncOQInUiKFVxd/NL/uO40TsTHHpShaEVpk
7arias+hZfNDMiqot6nmPZiVQcSJfxKFjs61DKEa98qUp3N34i2mSxGAlpf2IjRmPMFCENSj5GWW
wkMIqI9kiEDjQsoTnrH1vpzqSWVT96YFO+24K79+pCb8aUqQHaEtOpMgfr9jWnMBzGaLDlc//wLc
r4C5p6QVQJhqTCM5z7hOhoHuHY09b2q64IYSGYn5VvDhLFU4C8gmWIWFQmNJerGi4tJzCFmRbEOc
170VU1lZ3J46aVrGxWXNnRODgOGflNiJXLkS0Mwv9XLYhYvky/UBVyXmjKi39PGmqyTPKEu2tpCe
yf5yDsrNsYRsoNv9CHm1yagv71KL+Cb5qAlmHX9K3G8gSMFpgjiGRUOKBo5JxTbHiJKa4XDXKaUO
R2zTQAwM10c1DN9AAOg9SijamqctSVVWJmJzQNimQbrS1fs/q/5PDp0z5GcoGstG6W971Ab4OywU
A4Bszq1/260Qs0Yx4OmXCFo4zirbGTUugF/x/OPaXy9k8benYstlTTn1y9jcja3T5Lld4zopNW5Q
AVCbIzSlwtRLmY99D9eL23tkCJw2kiQ/3TASeyg/PrUN5ZNnTmS1oDSgAyTtcmN9YyekwBPpELTY
7DiSY7p4WkXDRmU7AQrOTwIzKtORGsQKFZZegd96SGK010ni75piAcsHqruDaeWQ8xbNQaQPEJbR
Qf3ZOGxpL6eE/vo6EjT890aOvvftjFNpMZIa8ig2STPB8RWYBs57kUSW+3bg0huV6nRqsaAEPOns
U3zHPuDtLC997C2hnpDnbm+YRWhfIko1GW88ucI4bRWP+mnrY1Z+wlhJm/i3i0duHIX+0U/VuU2j
BgsUWq8bfedkS/V2GEm2acTZtCTJxjC3g1XaqDZ+nmeV74lJjHqdkkJDP6lsvngPASGWIaaxTrfR
NolP3ADoRvL3vZ2scnSXWj5+HXSBje9x9EDCVc18e1xU/PjDqEE12qQMwVoSVT2JQjTCaFmhO6Br
tUUuyYD6SwpDJ+BOqnT3xTsAWtJzivnqZeX/Etr3zMZERJfhIFZpaMaFlh4t+xPGD4WCbytoBh6h
W0dzDk5+aJSXySFDeEIDrt5gCq7xbGjj/xXbvF+2ZfJtwz/lRZqq7lq5Jq6tgJblo//iRoHkAjWj
2g/Ug47wwFvNLDTXpInwssZ6xk0CJRSG8pHm43XzoFEuBdsusFc33Wdq5kdC/3k/5AtxmXVlJXm+
iNq6PQ4vNPzQtLtZY7KiUoseg77naEckh/6bd8802ocG8ijucaBz3Bmsj22/t6GdDTSma2ykJW2a
Gwmfgp6Ro9cubXMlgmypXZPkeEH2edO9JUEl4secpztLJvgUFHrzTf/bdlU94/vesPjCpwu1P2r1
BqlFU8rn7sPs9Muwf8yZmPj1U4+pGUu1GtPVcRdN71Ch+LQnlRGbZ2bFfsojhAfRgCOmm7ogNQeW
LUZInZYozhlmmWjqH9oDJEjAZJoKBhcZxcMgIEV56pmpVtLjwcdgCRdR50ARHesVuQUDHuRWKi8/
pwp9VFAICZ3qwmWIYFDooTWgDMamAF2hR4wZ6L7a/n9OKrwqwIjY8ct4oTEWXtKtpCJR4NeeYTk4
5XUH4aCK+qxPd8anai7kb9diA0us8OjbkksDIyTeVV9y+jxXz0wjYVCEI0UULEcfY6mbCV+JNz8V
xMyTQgK+VUj9exmiDagdX1ZGlw2hrQpaPDRJOqpIFuzFEhyaA8R0Z+g5tGPVRiEqL7dNJuwJ5LBI
y9/tKusxLbm5oG6nE2+ehHBQi8OkbC5s8yVE1R9hb22ubKDj1Kdrx2mi+AbDXpGH3oG85fC5EgfV
tjf4G+Bk2pb4tJbhx39uXRDrc9RSrg56zgpH61p1Rs91k5aoCoKJ+f24ugdjezRXez2+LMpbMr6+
1W/qje0uoSSwXsOkK5LzXd5BUGbM2Z0QI675NWKcyCrV0QViX8zkx75tbpCDTLt4J0gQmOT8ArwS
5lJDsHuchFdFktb0ND4ChKXIO6s3hPCp4eftbXgDqSYLnVNIey5HvcLIq3gKpIRO2hHtTzS40ZWc
Vo/A7ATBJZ0Nf/EmYiUzXilQ8/YJNPWAz5UlmJ2oCjxaNGM4CIKe+93h2MrouJHuGT4CO/J9s/67
kQDoylRiMOfXeKqLtosuGQ2fZJ/jjaiN+YHIzf8a++aJL9+g3XSMNfbyRKnDXbpZfRoGrFTygxaJ
F6BALZru95KSMZROwK6iXZfMyjD8ZnSs1rnBKnr/vHreM2Ck5/UZNXtruKmCPWXW/3NlBGES96sH
OGdbprTUYIcduhv8TDjaxS+ojGzhhcTUBqrp42z+N9WilWxPjfh5XG2XsKgAJhrnjadtKiS76+g2
KJFkynkKbJBFQVdfpCPq1iJgSZagZfslaDEF9TEoGU5wEDtIZhfG9YlnhxXCZsa4Os4zHfA8qnsY
vTz9RpJKhBej1+SMWW6Sxoo2uVHv1o+yPDLz1qZlL7rXGdw83KREtcdzbkZzbxaEdV0NtahK5oSl
2Aqbdgljn+2SxpD/n0VWcO1u6xHBLZqS9go5uyj/3Ip3jh9ColxshQrmH2+LC8uvEZyaWiFuUzW9
WnP98YTkJWBLWN51hZs+X22b7sdZn573DbCoBCPon+y3U3LyZ0TkRMIPYoqCnpKhT3ibNDq2bdk4
adUf35Qd57mRA4F9vFJuS72lPC/Tmgy4dXWrUTXCkYCOtwUJ7J+dxjpWVOuQVm6P3opml9IljMQ2
U4/YfVn8PBqcL3p9Orj0rv6rVnJtPXPhoDrY0K1vy1sTRL35TfWPVBSQWLwx/b1Z+/Ux70t4y0Ps
1dypL0kRznK33De5sHl+oXEbM4MqPzPv5zxVmYtMGQZ9ANKK27MTWnwdyzMNMaXVOFYj942tHZH9
Avq3MXdp3dPTBuyj+DqxWOC5Pwf0j+VuMcNV1B5ojipxtE32bA7OgYDhgK5XztDBaroAYq1apXhN
eAD/8fAI4x4dj4uM8kp7nHz6z8t5fGLzegXfn/PBuzHO6neTRdqg96kvX3jvgVF7GmtZIxwC66M8
2TwBaXsSYJXoAJP8jy2svvofkbxipVtrBWDkg7uvvvUaH/T4qn5Hgr6QXZrXNid4iNIgdlyUxgD3
PBXfpLlrcsYf50FgZClUvmQFG2w1Dok1eYo2E77RsdWnPNIAsa3i6/1fFlHTYMT6tpWVmg+cq3SA
OFV3qLhurdelYjOlITNgwd892+W3Hm2+yWoMZksnwYmxjk/KvHZLP58tTRHdTygFBElrRYLCygkh
S9xZxN5hyCs+G3a2JLK0g0gBXlDLOLDGkw6okpkiIoOteqiIekCjU1eJEcKL4FCIRjVCmmL7S4WJ
I5iiQ+6MbAOLk6Wpu+UrKRzvO6bXJiJJ6yhpXBgv/E3hnky8MQVfJLLlrJM9W9+PNugC7srYMbnR
Svl+jHSkwBSReaz16BlHeFnmWKELJdYcOKtA6g8p6NmTWjjBebPn4HvFkQTnquA2eyxCUXJCBLMk
ByJAmHvTEeFnpGKlgh+2BqL/u0z3XeEYJl7vk9VFFPaqLiYviE0v761acCN39F6UEs+Dj6t4QzeG
6RkTCf9MKSNinJkfp64aN0e2+ibTuGxQLIGPRsDUXvump1F+bWndLgAFVpEY5pD/k1umtDfWDp7+
60/AA8tHe9B5WxfkNMbQDzyvddtLCgGEv32RMPBtZiczBfPfVUNcqFE4Zm2SL3rNbemUR+OiqQr0
8UdKlCQy9vioOicBa7ZGYCw4Riub0488favlj7CCdN+ZvM9/38exGcH2sxozL1nsENm7OBKWCX8w
7ksVPpqFFIRSWYeZJg0xpG+tX6I9n3H2RyKI0g+5OqrlXFhx3/CepkzsG1Kk+N/Y+6WS8RVAXZvY
CR72MnD3dbLRsVabWcuCe6s82cyeM5zRDO4Wie2SVp3aQp9YW/ZmDWLw8s5IO7wkooFvBt+cDFZH
3KPukMSRwvGTC6RqGJ5bQuEG2I5vjCUVcqoLtsN/0xv3t/SQkY+sZ/kolO15L4vqnlf52q/fjWp4
809N3Uiifh8D1V0vteGCZzhlAwEPuOFtw6ZmMk2ex/0TerIAKXpuqgheNSnTAV3ds0gpgrgEtRCS
a8hWyCfeDHRF9iBMnTyho1229JrfulzRNcY/h51Vc6UCv8ILRjnhoQ8tuxY8OhVWzTovmU7oToHO
HwbstjHzIXitFzkRv0TX4h2FH44qhVBEomxeQU9DGWDmVKqQgwGGB9GXvPIZ+ZK0ArMSUqzSP64d
3Vplfo4/Kv/3r9MSjS6SYX4Z4ADvc94FkgaY1HuFNXOGDKMuHgQM5Ql4nhiTO4CQhGy1B+RfAV7P
znwyh1/RW6kwzTPBZaDRMdLtvhCQm8gVVRVnyr/ydkSeNIVbnPZHORxaSzVVsEaEzlOxWeszfQYB
Gpdp4WHJX32T+KMRee6ZQzRLtgfFz0Xk2+4uk1CENXhsHowDh+CmuJwamzXhIgu+6i0+E1gfpIAQ
LGAJ5FfW2ig0M5c3FwjHl+8mkpL2Sa+onpxY8e5Vuk9gKFGe8HS4pBBjjLoV3ks/JCmkHPg6b6ID
mbI2GfSR7gBrR6eKTaTqMWcPBQA+4CbepSIcXghnqDDvTLyYZwJDrzw2pWk6jBcN2kev2zetbv/o
2MSGdTAbRJcxWRpU1W3HGtO+vYfZFYmZ2GBch8wLgFu0qvoJ1GXY2dovrmssSBcLJxic/5jUafsT
ybKvL5zPwzY+8urf/BR0APIQA8BtNabj9iDn+5JiBWzIQTCwd+kVtA9MQPVvVZKjhX/CtzAcymkm
rZTXTZqI8QMkOdz/EcmnXMGv2Yd0KI19plYQ/yG0f2oWojLQ/cdAhza2Ika7ymlYXb9xa9aKroeE
J9DcSvQ7sa1uP8VyJ9hJfRC7fuoyoJcHbuvAlzNOFpjbQARjh13SWwtTSe9RPDbccLxBxDjFf51d
HP+UEmk6QL23blmMAUdY0zSlOOnLq4kHXbcNFC7DlNNJ1UmT0Hx1rGMGf/DWKoJJwxJekr6SWzIa
TESYrOkNbXIZyFdtv4x477JlmP5rQOJxfc8HeCFaa4oIj78a99A0IHFvote4VMBA3HTdRVRM/2Uk
RfF0wfIcblT+FF4mEOOnFi5Je41qnEa2K55nnEedgGfhXBeSwzUo68fxgpvXDFM26C00LtaP0qd0
n4XtnhOz/lYxKZkPTdWMxfxVaKJ0rpJLo2MgWXV1UONltLjdu+wrCmFnAKQVlL/oWS8T5guiotUK
8q5ToryGb4NqxYfkTjZZKY3YoFK7CmL4aCVPcUJJd0S1LtyNy3uUnhTgf56wT+rkzukSCBGBqAXO
z+3uUBxlHPop4u0smOL7+Y0jMtk3X2A0UmyinYmZPsJoaCH8uLu157KY9DKc/GBR9uzoUTxIOXks
YG6wUFOuIsNLPld42Lbbvpdu+k9Baf1jDSYXp8LeG4qQU709s3DzhQLigkrvlGYaMTIKDE2s8NGf
cgMK1/voQSThknpeR6UVJvyu3LFwh4RrH/q29GeqSvHERFIc/Hi3e5OEKrHBLf/uAReNYOVW1UGt
VYZSbMkOjustzVzYv6V8nKf+BEcnrjYOMd4iqAuUcTsDMX9dEsS8i2xnDnjBKPlTqHs9cKwHKswR
U6H5lwrVe83vV0aLtXwGQ89R30J3iiXiUvCXmWRBHQdsumHWO47cMIdseuF7ydJNYdNagB6r4AYr
Yl8NwgoPldLhCdohvfAf+JYt8HSSg9WmyVZ8oYL1J6aXDSfLYihLB/6VdNwzt06HhK7xyZZUlmTW
Yy5gdNc6JBX5xA/iKQJ8VmT1leO5OaxsRSHs1E/EewQHI6iFumkc2bZnxy02fC/txdzgkGTuIt90
SYImQ6MLLsN6xmvRpNCAUBQPjmW1R6YfEOsoTrJKtiGVZbiM78AFVfvJdDxFMLBGFECxOCIlPUPd
YNwCksjETxQUynMOogh54cFDXAUyshl7/af12NTsbiLKv/5ImzcYZPZ6LxE8lH+Ih66546nzMel+
O2cshKQOGL2/K76Bh/P4C2ck/OSrq0LWxhOqN9nZnIp0TSamAaBsf/UXNW4Zexqt5AartBmOAu62
IpXFYuM7r8CpKQkx0xGXVXcwRvHJyE0e67hex09HeFSeTVvUU3WbeYi2jT/YkdXEsRwcI5FkLrhc
gSXKf5WtWPWL7ORiZAx8NIpyTIL6H+QrbRNQ5LefqenezKwyvx757kS1iIPclf0FRLq/nRE8KrxA
X+W3pHc8GfaYUI5BjQ+jjDJ07r8WZlPo66iZSe/aDxSKZNVXd8o59I24QDCNfIw3mkw21w0h9Kj0
9nLpf2XG2lLyUc27UJmt2s5aRrcSMAsdnH9ICqkG8tKXtI5HxiF2Mw1tC2fkc+hcY2VLjiQNnBQd
7wCVyxs334rChE51ztRh6CZOsDTjQQyLE0CxNTskGbJnaEt7lV63q6+1BTQiscqmXkP2MwKgFq5r
0M8eYWzh0CtC5Pa2hzhYuspC2YLAbKHRMALEkSATI0rNiMOxL9vD5LI87zWjRdYZx8wVVOHW8B/L
HfFk4jIuMAfBz5RwMV41xbND1T8GvgWsqoPAsNJSGXkRX04iwGN2XR1T7jkNO5dX1fgmlgYhmYN8
QDNkMFbG2FUV2ymePiNV4DMPPFkUgE9wp0WY5JaNoVVyxB742JJpApq0ux7f1IQyyt5EQqCUNeOH
U266P6Tc3d2CkW7Feul3vilsZIBrv0f9rSMtH5iLZcjXFYYaAjxUh628ehvxtC8BJcRybvDDZaBB
zm/qknsSfsLM2pvNJZBs/sAJ45t7DfsSNp9NTakCaUyL6yzNnfo4Li0j1Skkimtl/GHcZ2AmnBYD
UNAdWEF8qvzwn+shq/wJG09dtef5udJqJU/OSV/XYPP3usNL3ynpfBpGC6gDcFNTU+dbZU7BjyeG
+NaLeGXSK/nQtFgJ4YyzPdF8YveBee80XfZwM+8VlcUsVE06GlGwh3PX1FbMt5ycICZtAxFXu+cZ
nAipAd1lzSCVHJLMjsyKGWnrXd7zvE9FWXXHDUAKKw5VXXMndLIgAMVO2ERz4zXbp/RBsrD31JcS
zCAOTM8NvQ8LQkc8/KhGPElk1x0n1X3heAnJ0fB4Vw4l6tRd0Xkm+K1EYvFFplb8YoTRbCIEvMFg
bDrhkSiQFrmyEfNc2XAVxSA0JtN6EViJM3WjaZ1GAY6v9mfMaZQmqZC/UudiUx8ot7JhymeXNCWL
QZDseX/JyszMiM8lmGQUs73QANHR3maSb+0sz6QM/AGaoPxr2/uK6Z+SfYZ5uPol4wlvxjJHMpFE
hkOXGkbcpyYWDbFohIFLq69GShVJMolLFqq1GLGSwNQYSTwi/GglkSwvotDNJ4dLsncQW4pnpObC
dcmxPE7qlyIIo12ow+nYLi1EgfU3/KUJ0BfcsnSk5VeBfzyEpIhrlbKDAmTomWIj5zKlZy8HXbPg
CGQBtEsRL+a4a2kTY1p25IVu/yOLfYExv6OSbk+ZTeZrTPEvLWR0um8t2aiXDbPexZxIc73M9aLw
bDxzF3pmapWjJn6y3E9Um5uki/SStwbiCJevHpV+oCim2tBA2eh2I1IfKqXWk5rN498JvQbH9tzI
Y36HJSmo+m0kjL9uigcBlyM9rsaWNNH/4ZMtWO85InCDyYYNk6idXqOkDASp8vrC6QPb6DhRVtT3
BXVvCNFxSO42guukh0fEMv4rzdsn5fO/F9cF61uj4Q2U7Nf1ElrNYrzD5tly0udJDcDxvDzfvGih
SAtuA0okDYbIlnv5KuavrAT7EcMRl07gCp7TKn2p2idwlsY2GpmkHpCn5LE/N9snvtOhytdQFar9
CYiBeQ5WSLYX82KUsGqhmxCpUR3+BQjljuZe3G+ynRpF4pdyqwFOda8k932Su7y5cdbvit6EVqUz
1yddXqms4U7oEbqvC+LFjPeiEiT450RM5KWHMRF7oJYmQnlyDmv/VnlhadRk30XZuCIKXVzzv7or
Pvv51dWbXK74e0gG64YSMcTP/rH20pVppPG0MPuJgHuKW7itMv783TD8oXV+NwLH4P0h3HO/UO5r
wq6NB8j+N6ZXbctbJ6lbmSUJ9Qo0bBxfXZSlZCpJkazET8i1IzQ1vxXjOwkso+ur43Ei/Gs7uwBg
oXH78c+uoWtHPVPbmYiU9n+kZ18Ve7ce8Pgk9xeqjaiYXCbAP8dqpRIpwcTRkJ3MHv1cI5gK2kPr
YsrynhG6FdheLSLpsD/Pe/6f7mss3PTZcY6q9Q8s4s49Xk5oCLg/m5IviyA4XuzTzhusJ50Nw8Tg
IHF182AvK841hK9ErVNQTbxuTFZFvzn50x6SuMVSJt48jl7RbHkSgj3TBWJJZMQZ16cCnqkZq1b4
DrUZ0paVP6fpcZUj9W7Y93Jo973Pr1UG3MM6+GzD/M4qssasdLAv2NARftbl7sP1+aecmc5OmDrl
2OQ1ww9MiMbrKYdeaFPhLMJE0imLPvJcOsssf18vUz5jIyXTZIOLdpRan7ZI4gL75i8q3ufyRoLG
DShmckEjJIid/qAVLah0bhEO4+HZHkNuucwd9SS3/W3AKkLVp7DxvzptczDMzKiYPGttNFKzGob6
B71DErXvvxR3qnxgXC195IhaVW5KXOZ/+PMy+P2334KWj1kC1NtmxsG3Ptk0PO32Uk8b1gxpn85j
G2pvMgEZxjlHh0Fs2lmrBioEHIWnaHHlAGqyVBmITvfMjWijF4iCAOivsIVGa3tXMRG8D+ifphsv
2SVCH/eqOxQXdzgJLXxo/VazeeNpm+Gz4HtVUfvlYE2cLDzeya/dJRPoGtbKU+YTpZDxYtDQB6M/
uN1Fe5JcLfC0K9m/OY9hhGwn2yNLTMrEuZx3HrFzjD5DCmpHn56jaV0/DOpEmPQaUdJQobqOh75p
A62DGRbkPB5R5n9YNRO8/HOPESe0ReEhuDsMFBt/nvOxGrIvW/w7ESNQ6KH9GmkKklLubT5KSza/
SngMVJPGjVk4xXaD7EaxH6UKGOZ8HyUQ6GHASw6JAhLBDC3XG7/QHMxhiXqBADfVZZXSwPwu4qRs
yXnUPZrSIlK/RwSGswxM6Nw1OcoiFk/ks0f+lqOIV3J+cww59k1x1ue9OqOMUXPec9q2tip1aba8
wwPci7D9ElGaR9vKmbNkuCwb2LI59Wt8DlpY3KxZgY4RNNSvZjFIrB/vbmupTMRmLMfK5P/3E/Mo
W9iuOHHJ2D4SODWcQ8y1dtXG73uGgMrK8Fc8Dk9Tz2aX1MiJkpAbKcadSxceSfFTJTJ4JJ0imgJo
B76rXtp4XvcarX5jivHTPgtj1YrE26e+8HiAMfvHp8ZnQFmggVad3hpOx9CL0QelT5WeujqFvVW4
SoSqGOuN/dbGnt9r/HFgGqii5Mjh5W8C8DpBPjOJUEnVRBK6kdwzVBVC4YRM5oDfLGHTs60KGHcU
Gcp9ooUFBtreAie51zGOFcUglVsEwaRjQi2RNlGrqc0Zaqx5jNFdcmxpyFyOVHAmfVMd5Ryn1DRD
PSOn7TLOF2sCbH68sH1HMOM4l2D9zotedL6zPCouzxUB9Tawm1ka9rdFbiLMTh2EkjDioUryod/C
3zbxjGYgAL6dt/uHzy4M41MRh2ut78PryImFlhSfR+lO4sNH6wz+Oo9QwtUKPI5fAJgH/G1Ve1zP
yN51T4iFi5IeqdK8NkmIj9Sz/qlbLju6eO5//GrnktqBHwrszfiJzNZJVoolHp6aTLqGtCgz7pNP
mnQqBvM6h2O24E0PzS6mFwUj1zjnZzNfMDzf8HlTQZG+4fBWUnXKKNh6FuBlY7HhDRQ/pLpUgREU
iTITI0w0OA3OU7UFP0q3QtYHew71JYaaaEAszt293D9D+vQz34hKcqvDVoymQb/CA1z3QMMu2QPe
9ECW9g1PvgVamLc8lT1CnuowjYFxGk/W1yuSrMxsaeXlH4B+52OEMRQKJa8DCGAsgLl34Rq8yNvf
r2z03QZNXxHqId+4FQQoFAHz0Dn4xPgild1Tpup62awVe78NfuUKq9P9hVwFw5EMwMpr0yavsmU9
U6dEX3yhejR6HuWl40y7Fyj9LBOSBMeRuaPYUGNrqrgXaLGgmA44xbz1xeElHZ53BKtZwiC1xm+3
HLfyvH0RHjwOh6IiMC1igTBl52QvpyCzSuVDnUksAwB2mXpzlLkufbPTa4R6fngTpU+nO+7siDDX
cQakpnIoo/5oIwtUGfgK2iFJcRjcOiGRFeUiBPH9gKaFsQUMFxagiSyOaJ3UkdVZ7ueORDgTIvBl
96hw/QOI9mLwlpJFTivIUQZAz4Cih1yf9x2nbj+RFBAj5lwvjFm+PD13lNLXZeqRLevjw2NlAdPR
Z9KsXmPZBIY9NGh4l38HR1r0zSqgZ2Doa+Nxn6fOY11JfR8Zg8n3pOlRkxe8iMlJjCzHDDBoFRbN
1r51ZubhiHCWqXJYlT1VEfI1dmOpfPg8efqlmpxVFQKue6Cis++RQEtdVp8TbueFeicP8xUZtAK7
14D3TwlmfCG+nWIuNEJ5fOwr9lvtY0Fs4IbFDfK+No4ngvSWL2a8F17AmlIrCEQNOr4j1rT/gkh+
WAFDgWjHc6BAztWMBnFdpfL1f2KkjLJrxs5Xrmw9SdyDpMMNH7abafhqyEukBDDtvwt0+Txm+7iP
OQ5N7Xz4GsaSS304CcMz/KYr0BB3TH5zbsIj4ET2vqTFiZnmvmR+1JwQqoNvzCA/0NgSVdQNVotj
OCQzzojd+3BEL6YIAY0E/PcIa/GCDhlu5ePq+5fHiYwlxOoaHQBI4+lGd4e/0/hAStkMlr4FaYj4
Orkq4mHqSl/e9ojwPxq4UzDpY9M4J4yNOD6zEf1jBh3awI++F7OtBBv57GpBts08PAPNgiGDtOsu
NIRmW5CLP9SwZZIxbpeuWco6ooS4Rtb4yJ/U95xrxx0Tz22TZUeg057WoV+mTn56uKjvtSpGG23j
2xBw3LRhlzhI21CSWM1uoipXxdzHkhtk7follb5CnphkYAnGFjpj3gMJP/p1Q/ox3UHdXWKZCEkN
SJjlTB8xMTzgz3n69cMBuO18vdEbTEPQ36RwPf2nRhrXvAR4BTRpfT7rBfR+jTw3QYRRRV/EM3Lq
eeEZ/KBQgRUMg5tHTxqapeY3S1IzGi5dPrS7WJx8XFo0p1l3Ovi3QEy8x7VZCJERLVulmycuNds9
PgYP8O/N/AzcOuefyC6sGY/lRjXPrFP2AUE6YLoCTsq8U7tuELSyPj40eixDSOq4k1mO+G2EWnWC
HYZ6oQYRd4B7+IqZI6KJUjg8LNvIPO0byY65juqRVAAw+fI/mekEE2af2lL4ARYOCBMI7CW69n5c
aOmfM5jMf6L2eKoGNmEEVzsnbDDHXCwfS8h2F4+G1cLXqH45O2fqWTIrdUPZiCLVdlL/b7Ub+EbV
XjGGs6h8smjDW99HxbsyHRjsv3Fg4Fihk3tD//7b6VDqW6A9tzwWI0lUbzwJxPmdCGunZB7OKqsa
gBVSnc5HIv+xqr3GV27sdEZEgXj+dgM6KsCLAzDk51/meYDq7v0Pas9d7P56puvgmwzp626M9K9y
B7PMU7v9wLfTl4dqeugiFI4zGuNr+1yQPsnCRw4Slu/QOOshahe6r+kdI6bJI0R/VdV5a+FcDj3D
S0cSHm3mZ4T2A25lLgWIOiNs5f44HaHR1dJIsqZzsC9VtQWQn4sj6cyi7RtDf2pkmxtOwonF2Maw
50u4YwixiTRc6kKtpacDiEHsbGNL+5iQjOE0xXA3eCS7UIL7tQnD4j6EaiZouitatOARYisjPJsi
884XwylLhArUpOsgCKkBoUJ/2RhIV4nbs4wYpTm70KUgS7hrtNyBd3dC5vwMEkb8LglnOKtBOU7Q
VORbvj90EAyr8nR5w33+CvkIBk//2ugNIjfClZDARkpfU5CcytteqI+1+s8WWalfnjqrqkmotal2
vgLgPh7DTj28uPijIByfx0xW3N5REgV812khw26rN2qCQvJ7pFWvqAADHx+yT/ie2t6GjG0Ss1gT
uwvSvubjFKdx3fJ/h0qgg3cioSgmtQPaAzOU71lQCz5ytRlo+Y8WkqhgMz+SS+AkElTsNQdpKC0d
IJE4K5RSdWSp08uD0AxemqQt1oQwmZJhAQJfKkUctVVd/wi1vPTmpBpD8v4YYChpdbp2C0l5FwtZ
Ju/AbipSHDlR0jYq8zxXTQpJvZL287uAQBhWAmPd/MrKy3DDB3BvQIP7/kL+acyoQYaKEQGvFP/7
NQADRwcVKkMDVO42lwTKijcq9dj6thsT4NBu3S7oAWazC7qZ0hufCHtUC4r2CCyoFSSsYH29Vus1
f8+SDHD1F0rZCRZHJ9uKrG3BVswta4fgq83sno4b+z1dvGefGszNnv56m2eQf/iqVXXeo0d1mhyx
04kulm0VeXbBld1Do3ow7C6JA74Xt20UhP7fyC81icB74sfB0pc2Opn+JqImcWAKaQOxHWaS7oDk
gGlkzpueYqYRjMDtNJ6OyWBD/FRBo14LuIOFQ88P3Cljta8ZJbqvl2ixJd4vftc5I+8bhNYt01IU
qIHPn3y2l0Xm/MsZpJ9znijRDK9CS9+zM6kCWvR3BKUPnW14QVktgi01RpQqsLV5JgFL2MW7rfJ6
IY8MlBrF6DEDwI5Rw9FUUrl36b2n/ku5eY6OhJchCnSAnTS6JfSDOdwfL1l4yoinMf199lBZiUdR
NFDqt+lUYLST5cOV4hbv3pzSF1TEu+jw+BHysun0KwrTYNyk9/DCAtwX/20koKOgA15AMrxSJCQN
nZ7ktBYv/so86z/PnkM+0NsWdhCeNibgXKDlBJRj+7VMFKAZGw2V+PWUcJhF0WWIbfM2BEKhPU6P
gzyM0aVeqKiyLA9chDu1QmCy9Fxq/lD5mdOuqnM45h1Q7ehzeM+bqGHa65EFUEDy7RbTywSGjWwq
ffC82Xnmgyv/81SPX1kuZ908pvxHxafjtpPEiG+AYFBBzifVMSMmGojAFoVPB7gOiQ4Mrg0lA7Bo
+lPH9YVcLtBaHXa57Kg8PrmuoxE1F0/Hc6k60qSluq9zQ37MwatMXC0kEM3r6so2lNcu8/EXNcaj
PXF40z14dVrOvDT1mz9xXiamT4/9d3AuVUHhjot0nT9wCPrJqC64nY3uKhSaIylpk5qo2noTVjw+
cd7bdBkfjnuugM9l8ILsnCer2XWqSFYV2qrxSlmBLvbJRpMLScpIEDBpagW1gv6xN03KfnfIJCDQ
Pi6UMmlQrMmwXuECDF7QAbMJUj4CNDy0jVJceIlI0llxUGpltmoxD4tBbDrf4hY5xfOkvVuwk++v
KF+t/5+8KBpR1Ngw8w6ZSKAD/EEINiN0U0jz4lQ4PPzfdQ96Jz6AhKLDof3jEHIk+Swmtt8NkuqG
kFqZHp86QD/gHA+MgcydT/akrIn2q6+mM1Ri9iIyr5k2JtMcCjh97Gm3JeTtMdIU3D+3A6nQdp2e
biUP2kTJm8RDGOBacT56MxgoJNxQzWKUOM6GP9GBJgveN0pkFhkE0bcQo8AoZjiEI8tZCWV43djj
qQshDLSQqvpClbeuwxeRO/ten/w6trOzhBvGY5qfGpGpJNOhKxKlwQlPB1gvWOjNaXV+5YC9FXa5
xQdXXjgSltj76tuIEcxA8bf7BgpPg99IKmGe4Vmlfbtg8wChEVDeVfdXQnF4/Jw2dRzOi70VZQWu
vWEpah2loNmB8NWTaegUwc/o3Ik4jubHjipNVDZNw/n6XFDInJISqKR4WxdB/2XJgdNPWcgnTiY1
+6wDGJQVwRn+V0O+d+l6taJutjErtt4sGUZG6gMZy4FiaGjO5MI4LnWgchYeuU/mYhJwl4d9kDQ4
aL2/D+MLxBsYY66duVNOuDIgHxzL5eYKFfsaR5G3UWSvYmCHeCr9kEq9JQVGaM6JUITcs8wfN4bl
Cou4pah9G/4QQrCqrgQlZj3/EXnzikQJHARhQk40i1voBPPMi3u7gchCgwA8PkAELKFT3qdIjiC4
qcGJL8gtyQ0JUmB5jRX1LIRWCd6YeEo0bNgUXUW7rbaNjiJ8cxRupfXUU92cny/ZrCuyEADc7bIk
cH9k78ZoWybO9h5o3laVVF7nf9XO2SxlRWB8TMGTR0KJtEbuNqIbJLrynXcJmTSqcvJ4sYjNpLN5
jhaTr5vvqbjg6IOjG0bWeZ24fN2rJqHShLkYZ6MM6Z20KZfOw02ecshZiBGR6f+O/nLR/jQNQaKC
7Xwc8/NbTslFCJiyJnWVAlCE+6DQwHe27DDT2a54bPRY9zGxwFvijFBZAjBR8zSOaQRejwrVBmB+
ClbCNN45pa7zeE7WtM0SBi7YlYqr0c93QT6pnICqHAwV+Qa3j7H5UghNoAARt5A5uS1fc4mLEKcO
cMDHu74ulsoksQiX5UlkiYTnMuFhmNQzSxkdIIKGVZ7JWlb1meplh8bXP2YOV+9362giTCwWkzim
sWQlruaM/f5/Vb34ksji/0zWzUzoiRcLAVuEC7ohdkzdvLUJbM9dI6PqCaVIJPPqUw/rkROOChJa
Sxb98V2DMnY4owzqgN9eobtloXxm+ylE4Vno69Ghbu9wZWUVJOFt8X4rvAT/B7WKkVONTcdl3ffP
bQ5put8De6wTC+1cR8XfP92urnRGvBYF2kRHzdS7WH+hpX+WGjZZGydvvIilYhjHOdlBIGaoi/9o
LQXjnvdMyeWPxQUBWG/Llqyknswv6nIbNBE0TxgAKU9ufqObzOFZL1gkE/RoWbD7OJMG3qRLlP3g
oR8EmMwBqov8gigXHqWDYazv9zdLu+19uQBr+brcZFivC1H9xucvH8GueCiQihJIDzj5VHf5GxFy
PoAgoeBWtKMojlkRrC5DlJwn8elno6Z3C+28kNZSqI0IIcSvniK90kuibAgiRG988aGgOlK1xKcw
O2M+jSLola5lezHCZJuaLMOlEHoxca3yqgoEDyYHlp47uKTrZGYMS9GB71Wuv9rMJiF7EO3CnHfS
AwoHeMsa+IgbvS1fZl6Uy/j1tjYTy+o0FeTaN0vR4XHJvpPQVZsLX19PxmWygjzQV0GbK8gcoTbL
lUnCuZoEE8MvcJSRlQ1LteH8nirUa17SJdptJftOLpqXIwCAG3oxXXraGEsNHapi2cDK/awAehOR
/Z/VJryNI70Q4+lqVmzx+EzXPh4LENQqTgSSoBSbOarMF763zNhjn5PfEGacy8djggZ3dzKiCjgx
ZTkXs8kLJhlmr5STx9ooSs44ROA6NJsPvrcPg9h86umu/kTjK3JLSRaDMYaNtUnjcb3eB8CiS+0M
bAKevSDvkEDtf0HOOkAa5eBqq2Irjr+ATomD/JqXAqOw3aIyNBB11A+Br1NF0jyoA8sBIwfJlvpN
gDp1vJhgVeCRVzR2pzIJsdZZaWUNj5ImZAVyZa/CGYJCvBgNO9zmRs+PYGlyQXWJmBLoSGFtmd9N
h+/dCcvYaad41hUcTDwIeqPoL7/Nm5bQyjMttnIjhXUq1DYCmI2au/Ll3TmOKxU2LBKRxij4H39x
WLmKWBTYXiQkgiCMgs4wGHCR7QvFvReH4OsxDZ0+W/wZSAU/GZJtD+aBgPPVuDTORTOg+t+CZ+m7
+TtL1WBOX2/1qZxadt4gi164sJG/oOpPABqJaj+LLMjN340dK0tA/sXG+w1V9G+7x3Sq6v4gClaY
gWhW0gfWicFLGg+2dzdhjfthudnr9Dj9qNe8CNKdGBhLE8PkDQrX3aMwx9QJCS1Ysu2Nc3ZlfzuY
O5TLanNsQ+YcWflBQTPLbpiBI1dGv7P0pU9YrnFirjxHJy96hTVzDn8XbCJDiHUs+r2hmLQJvcOD
t1EO2fI6u7Rpom72ztzGgX1anX3e8zo9T+iSUyRBqs/ToxOdRUjQKH11xIMD214BilPpFLAhSdnw
oZHctYSc9w6RQTeUqKgBY+nvj0fwVPC6Ta3CNdPN2Ylf4SztHToWxHmfSXp+hss4EJWshxqHwUba
ldyXt0cQktIfi6uN7kd0yr1bpx7Lm0mU5rAMUo4REL9+cTIjSipU8r3cD9ytz76tcJbvd+BqlnCg
H+/SKhbQbL5LQ5MZNrS7YDZjPfQl9rUXg4hUfZX2O+Q8DSom+fw862PUWzSHmuvMM5eWYeZQtbGq
5oLX7zoGmGfQLE8tJYNxXpqreQI6WEqOahOnjwhfKsR4Whi3B/Jon/ggX+6CyzBV4Den4UgB1Thy
FRYzYluF3aBTOVAqOedP+NpNwyJeqmAPFQTQlLoFcqzd7dU4ZL0ptyMk8k4kRvZpsDvHb/TTnvDe
QIHcLAF48cUj5U1NGk2bUB28M+TLPF8BMBwC6TlspbyLoWoVczHQsqcqqDLILHVnFGJMyzTIF6jr
+GGe0M2IOm3nEqWbiip1RtEDh4EdI1dNUpU0knQkBHw87n6Y4U18ZsEKkJohMKeDIvAdoFZOsW+d
/G/YYhHZivFSJYcdTbZSxRAOaP4n4Ajb5KVtaEFmAt3wI5/TNX0CctUquz5zZ3+6OeSzhbMmqmR6
mKQ/0Rct+NTKLXM/EIcoK5uoWNNRQKpXZ8GvtEX47nhR6JxzJlIMlQ5Og+YBPioRrGeH99AneIE7
DaE2m/sdmbLMdrlkXbhhY8Rp9KP8EwbEb6dgMlh3Yozyk4KNKVJ6Ev/VM6aFPcHVr+P5NNVxXF+n
V2tXfl66VuJxzVKVYtbZM5Vx6+6Vmj3KhE0rG1g/6tuZe0wEbvHtXvdgWma7J/Y+ME1gFjRu0AIL
9mATj3ethPWmdaCfN0Rdlsc9lOoXzkTXO7AV/B2qRS9//3LXRNZyrShaUtkiII6XQVzZEtjOhtQ1
oU16Qj3vqhfy2PUcC/rrVqxdHSo8rwDmmoA9gXZEURrnEkcoNj8GAQAVInTrcwOTZA6qYcJoLAGH
3Z87ucLoO5MvUxgYXD/3U38pXkcod28SuCCQu6+St6pgCEyIe5rizx7w99uwJLzjlyOaguKKLStH
9v/tiz14JwEA+ecu1n2605ulr6KksrcmLeBc0hJRsVggIUWUe4rFXHEpi+19qsyHhBtpUbABslu1
mb/zL+FLMl8TOVH+frpUc1HileTNU5V/jyEgBymujTnJ1ARsA/3+jq4WnBskC+X0NINuGDPaH3NK
fRCFsAy5Sam2e329FdLDKt/wSbPxtuJZSpc8vz1GUXLXSEhtJHuGSWmvWZZoEFO9tbN/QxJqJYGh
CPFjr5Ch2wnDz6ZNKMwlEfAFJJdtWbceEJvv8wzoBkQ7wLGq2r1HrJxwkBaV5k83xnojMmNe5Lye
vCqCfdpZdS6LfeL62iNwpWVPj486nm65Gkqvt2m2rDnXbUW+V6nX0oiwVgBoT5x5Gwr3MaB89t99
DI8yxfDrAfEQ9vl4+j0JwU/FMPk2P/a7mehm8zN2upWDKVMDfYq8uIvA3tUIptGWHKMgexubbVNL
lbJqUB0SoVwJL+W38iqLDr8xD8PlDaek3CHTjIpknHsFMgdF1QYJm7I+dYL8Cc9sfmLrIY0oAMEV
cNPO9AXlF0LMWj57LbID7SC6/4flMG8sqrNArGMNMoGDJFn0bxzAmmcRMTZGfgo9InJVqR/WnaOm
xL55KE+wcKu1fm5IUnk36oLp6stHm4f+8I93UoKB5ruYyIlUkhyr/fLKvnTz7Z/CKwf5ougvWjh+
m2/Z4zq3/ihNBe7wH7wpvXPO3fSA2J4IIz7OYSkW+o9H2gHF/zJf15kVlj/eS3yibILiwgaM6Sc1
gzm0H1CbnJI00eesJITSPhmlDjJ5/+DXW5Dl+ws4oI77HCam29N75YaVWODes7rouRbjVxVSCsbX
S0f/QJ+rKyvPYvH3qSuAD5XyoOHdtbQa9aHpPvrA0LP1MXNopxYs3Qmw/UTr/QhiMXSVXtIW5yP2
me691aH2a0Ud5MoAVrtGU92RiTqcpEZw/APAC0kUl4l+6MvtRRxT8tHjgE/zfCIOaLfU8WIwPXsS
C9Gezd2iJyHVsZH1Aa8XSfaVMPykzDrrJlkq8qYG4v7a5dNg8XTmN9xzG8MkLrZzZYs8Ubo4P6Rg
6HOltp8GUisgyxSiyUjKGIif1PAo8b4CNyce/wg37O4H1KittztgSW4xRcZBFeGGnRzuzkiB1LCp
4aaULcWn0Edisfoq6CdMkhd+zg385FkayGy0+1p0jQtJch3gPDuyZoJvEvXjDh+hORVKm642Dh/G
mET0itSQCuw4D5fHIrqQsT+Kh4PbktQi1vDnW8iHpHQD9dC6qRZc++g+gcFUcuFul7qQ+TeDHpim
h/IQuv/YwGmd8GAjqTH9LED1Ch2y31mxn3IjJyWfAqAGY9M0Zlh1xnjb44t9In68AZrwlisYuItW
PkrfYRaWy1K1CBukm1p2DBU2vVGMkzi3hTx06PwV+p2qwBLRaxI5b1Ix/mTNtlvw0BgUIZKJ4mdK
8BfGU0CWoWpDd1DCDWUYemSyvJfS74i7SuGpk4Zlp/LoPyD8QmL1mCMJjJ9xPWlqWiwT1eBnHsXS
WwsiTvcJbDfSDBqxvpCPc9QhoThkj4jTofI9AU/qtprUFW6urZzcvV+U5qxyH+bScwv54Zo1BLcI
l+DG6lCYlr5n/oTT8rcywX7+iSgGzpgByBkONY5AgwUNfIN084HURHg+TEK0P0BeMb22jRrgJHML
bYLSlprdzAe+MP6M5wtRx1cnlF5phLi8UQpXT1sh+3eL3FzozB3aHXlN1VKzTh7S1149RmFB90Iv
7YqHHTY9+umYG21YaMg6d3FiYpMayeLAwzDTP1MkajbR5QsTJKF9DkO1rG067Qg8dRwhMEmJuvis
RoWKHtODzQ0gkC4Vwdr8z/F0sxDGC+CDLkn5HJbaS7eZn0kFVgqDhOwblNK/c3xwtiAsIb/1fhzH
icfpBXUZgNYtB8EEQoBjRZCGqorD8Uriw5kYmS5y9thy9pJfw55rHgPOyJpSI5LxZGgczIRF7Mso
zoFK2TSovkVQBRbQdshmVP/RExbsUlMqUkTHfl+pxw/5fs87fe4+XIV1uVoEpWVlxinUhgKYrmCM
KDgbTtrTrBxwwf2TfwRdIvNQdiviFJ/K/nWNPFAJC4tb223BTyuQqI2lzH4bo6Tkk6OrYo8l0yxs
iC2rZ1U9O9QQ6E7yQnYHvDE3v9aR7StqHpU+C3YyMX/NHorQn2CxMRsuBg2kZgSjKk3lNqHk5Plv
QXNrB67hdrHvDRoHajZoz40GEVa7hLnAY3VVNTZqj6QZc8RcYb82P7/ubzeQUNgvczibM6ngKZ4t
83fSrRqvf8DWm4Z8iAmwM1llRRzvN1Z7rdptkKbUJVgJd6q8siggiolm+DjwczBLwEkvkHjvmSRX
zorG1+iUefWwth4GXasCgqw/dCUd/kqSZ4M9HeH0LzI1rzEG085E7ab6Kf/Rz2QpdjF3HtEqtRGV
a58lCRDHjrldA0iOneQdTHqXAiZnMP1htpTKnQwZtrBc43adqpjrcgKriJzZCH53knRoYYUB5rn4
9XQUljc8cWFMJ0/m965aP4MBFX0PG9E/cdUDNTPQbQCIEHMcuv2q7TwCn+6DhBr5h6xSaAvi1hzC
Fup3c2InX2lZCXDECpMYLkygeil/Iu+KFOikJkSV4zh8PH1zLv5PWrl7PP+gW/gnbHkYG2V0wHpM
rckqD8k2mNZ8FtGiW3/JpYBt4DZ8IKftg6nR0VvDCozm2vR+4Rln22AHcVeNhuVIrR5L6qu3iFB/
MoOL+IgsPCMa4pTgaXnQ6+3OHmDpWNgrvKr6jJZalFRiM2+mIBoyqTcfphbRTfMSKnYnN1DJidPQ
LTbIlhbBzdr7pHuy1nqOkDuCvHKDr0IKdxVl7ek3fWoyWjclXvevk7BuKPT34soCsLGIDasH2NHy
DaoKwsXBzM5bN0O5FOTq39BLu/EtpJn3D+rr2p7l1YCiIkBMmKFmr9xqr4On7i7HwmDp+oAZR/yw
MXr6WRxVNkwUlS2OnOuomoBSN41JXekQFJTfvST9M9oo7gWTnZ1r5KtbKiG5Smw/VN5DaUhJpxJn
9sei6S6qg1hRT8PhKeDZ744moIHzIXZ1AQMAQY9yFjFDiNEPU1F7ypfij5N4uAqOjpePbYKBRMND
w7t49joNYrCHEWWCDrkDMRlthn/oeffOwBsQPCyisENYfZ7O/ILXE9vZ9y6WJ+0Z50i3UjO/yl7q
oSCxzARP/6+x8/oCbIgG918e2A3WLEi3Ugx5oXcEHWYjvdJ/iLvPrHvUUmMPUg3YQG8r9sHI35ss
mrPGeYQGk02+x9W2IZqKwQBu3R3XL9qRRVsIMST1Teypnu2NEEFZ+WxP3G7mKFIMHffdzANailh1
MKTftgAfR/6bz2l6B+kiQ4tpIk8ftLfaz1zBzFx+x9DEtTRkxK4DFaM+Lvdsg+GHQSidZCmfztSd
9XlYlJBrmUiZQjcTlpuwS0bcCxX6Mq9DIN52DKWN0ABZOOd7ajCJ+LgVP7ufNnqzU/7JMgv/7Eer
XnelygOVnWxu7ekTWITU5F5oU+403e21D7rIaoLKKpuIqeXmnowDztYwcoxGgpQ4dWlZibzR/Emg
W6A8tKn/HgqBfF0ZIj+EKUvM8Q/mtORMcnx323yhJy5ab7fhGHm0Amvm+y+B1P5rq07+tP8qtfXr
5zgydQX/76yD9IZAvkbLiCr7booYoC6zeg5lvNMdxAbugpRYSzhhwvLhUwB2AafeKC2fiJ3p6X7Y
Mxr2z/NKgmHyR3t/DQ+8/iQyT/tO/Y8OraXucWuHak58V8gUpDK/MJlnF9X0d+9fHjTgPyComssb
R56ME+2HOE1fOyw9MkCHJ93jxUq4bQcekwckAuWHGsxGnx++yg6AvBV7UAdyyEtqsKy2VUbSyEv8
jtod8Mjh+y7g45SiA5zBWv8J9tfI5Ga2TsJVrw2Vqle2KlpD4G9Eq4M7j59+kvA/Onm7NakWSs95
PPF5X53WJMnJbDL5lnvCY2ggCUGeQkLqi4s6lDlCUNhVVTqV+6UKB+f05e/cZ63GA8zQJHwTlN9B
rPQB5qwnYP5/h7JOENM2XfNG6SqBVB1/xtW+zbqR/8oc49O32+jcBz+vhdTs8nE9voZ5WIVQHKoI
IF1bmJGxn0ELDEs5+HcMYi2yE69J4nczs5/Oulki2hcmzv5TQ2zFlq4fkL6GmfunApEyXkILBMAE
gFallS8/W8DH21U2YSF00viMOqzRDyYtqtlGDKm+Vo6T8SvUjkXJ/ej/E5IwQ1+Gzhd3ESi7StxE
fTavTK+mgx7V5bI17BLcrXt/ww11jB+ynP6p/Dd1+4yZNpRswbioFE2CI9fDZSljMW7mHPZjI8W5
UWG2Kcxjh9VL99Cb4a1ccYNm98G/IPLBLL43zJiMN9MyGz39XS3PDoykBii+6+2P4Dc+dd7Qp4wc
T7BKvkLAnY8in5yoxnLoOlPyCtM96+uFBCiNGZe0Fv8ZCwN4sWhV8ya/6I88poQMh6p5N4cQg9RM
3BnXoDbhO4Mb/osjvteBhrBD2jdl3NzzNTruIR0w76AHg4u77gxgbiGKsEIrB7uboqt/6oaoxdWp
FUnKW6SX7+ReAl6KjvMNu4wEVGhXAtsQlTaaeG+APkMY6xb7kdxu1Zt1uYKIeS31JYZRBi00jwLJ
SdvmZxVX4OiTkqyq1HDn1NLSw69mcwrqpGlaqF5+II9FATIIPtUsOKpHe2N4L2MCzvWm17Ca4onO
YuHU+EWSRzdiF2FikkBUwpuSY/lq1fkkEHhMVBnuG0UcRk71d5IjE6MyURRwz2/VeUd4zo3ZPJiJ
jCYGsKcD+JS1ZAAqOee1yX1qWMVFFm3BZ5B8bt1rSF9iUPSwFOtjnY3TE1OLgoo4Vh6Q4I+UuIyr
imfEp/KheD8m6yOJrWRG+f9FeDU1PupFvhFFN4rjtSUInYxOOu0/ZkAFbQGr5RwwAMs7zQtMV9Zb
IcOxl0y/n0ZgWppLv8Nj4oHyXxya62ga9KQp5DfGX+N9WN/AmCRAGFUbDHDaW10BBxhY8irWW/cA
YndC8nelpzdoyQEM4K4xKh0qRpvdnepn5dYDgyq2f7e7bXAvmDsGT3AOiVJcFMX+i0C9F5hbPiy1
kbDrkPks/qaDu7zQpG5pgxE/YGnZ0PwpSPeuDmOiSdcivPloWxt7UclElrgbisUCjDlsu1Z7d1Gn
AcQLpwv+75NNYk/TuV/oGNuicN1W5z9/4YPHqC1TGfFF3tJ42VAuBNkH9luO4sPeRFUdCDJjqZwV
MRiaV8b27fQPhv2t0U+L1HW+lMuQs10jDtqP0+/GJKNEPEfffW5JcuXd4tebSXG19jpWnTeSjf7m
qsjqXr1PfJfw6NsW7ETlin4/y7rxkf+h1vRM9x+lQrrGt3jYZjrD02gXAYbJggHh0vc6U47B9rMh
wXGClahne1TLTJiCtOjv82+3jp2tuonVD7ej+vU6RspYJ/INPvCio2fZ6QzvL5W+tc+4XTZ4qpIK
eX4gbxXC9tZX1XYpSPvH+g6aH+YTmFBODH63ZsnpctYv1yO94+ujXqxLH9nRJpboIPGHkloY/2yG
ui8x10EJJKz63iOFf+RddTm0vAH9CkCGCZUcxJeh5U9cNKnf4L8uFOaRF6HE0mfk33YcgIfGsaG1
oLTGi1eiyDsPo2XaujFYeHQxLiBo6m4Q5hTeLfKuKukdaEADNRRbknq27TxwZeYlINRP7nI1hXzD
oSQtpxCPXkFhCAYdy28G4oqgCZCEAZ+Ix1RL3zgs02mB6om0AOoUbHvb6Vebb/TrTgW/Sf0ObeEZ
NSgeE4o9hbfpjz4yR3APOaU/CnZ2k5G+tnBU6c/JuHmlp/X3YS4iSC1npNqCgpJeBJosoWv9KsK4
tgWksj1M4GPPJXNhdarFMbcRxTeoTZ++4WvgOzQ18ybVtuS9BgOfpLp4MeO5uJgiSODCqYrBB1+G
H/S3/GAGqT5gN3MP30ETYbHv/a38aweAqvHECVmgnDwNdsGhybdqxwBIF6kudbwf/r8F1IX4mGpb
wGsHUUDQ00Q7XyOtAngjmiGCbN2dnXFg5X0GuVwttT1SESGpQ2IVx3q3oba+hSBAIx+yaxkv9sKI
a/s/RxD+t1KgbWZ4dgKrNJs0y/uCxC2xxs1OdBO2D0kLiiScv19HikLtVAa3LP9oeisJFoaIwRNt
MysNdHeX+s77uLCZfVUNoiaYLyoLKv0EH4lJT2NipDYL/6W5gmwSpvzDXuwjPrX5+EdXcGJ/N8T9
PZ3rbXKC+nnHNXsHN41c9oqZc4azBDAhK5Wlpmfh8Plt4MCEPkT3OawvTO30iaQS/xG4BR0sgfxd
QTtnk5ZBhvV2ZwRbGUJDqXClew88eIKpVhwxSYck6W+H2cABoo9jcHeClqpvdDAFjIBBApigBL1a
BFbmhmIxDc6i+bpo3OO/1jtCkJUEBxj9JhxbZr4IbqvKIZFjfuMexDatvokvnVk9n8C//NuNiFk8
afc+wNjyAzp2i3nAbnEzWoYgaPaUjlWsqMzQeC6r+DiC0Ox3nfBSljN7AFlj2d2w9DZO4aRMBSlU
beyKluVHmqCW2vz8HhuCGzUqzoNM6mvWrRYaiKaOeFzRwFPZOugLMkyNvWnBvpi4rt5VFyGEZJOx
1IViOEbn3gE8nvA8RcbTFtIy2AM38AWgYrVdl38R3dXtFC86zP4JbFC926Uw6WG+4qpI0pS2dxo3
cQV9gDniybd4qQwAHkIACp2dJhWO4Dzm1XpYsxtkL/m3K/LoDGadXa+jaO4q2Twp8wQp15BSRzEf
QRSBgQlHXdCeanV/eR4cS4Rigy/H6e/98MhfihVfMJcxfhFg1NB80u8unzuMEdB0IxEHQqKu2QE4
he/glwsgUEyQs7O/NOlBuHveyIwa6rjiVDHN8TdB0gjGUpYqlD42MaCBLkRpn3J9x2dfJBSDj0ze
4mN+CR9kn0aDriH9HcT1qMh4bkQQZzygr3KcI52RjLBajhAi01uSDgUxywbnsMshbi0TYh47DGaZ
9I+ycK4bBBjYnFueT+JLnJPKYXBEIDgn7vK9jIUeiqZ4vxMs4UhjWKtj9HL0x3mf0xGWWOVKQ5ZA
m4bAVG24BLrmBjFSctyC+UTpARxeiMA8p29icQGdbDkW1BIBPY43YjO/KxPc/RqfOBSxo6+z3L3q
FT8+U9wWtKcl94CdBeeGJyyrdfeBgvFljDnFYiGJYDCTx4yXDw7NU65WTXzYf6tO+Quxj9CwULZP
ZOQGmWuv8d+lgp5pGpgZGp0GC/U6mo9BericorzeRgoC+dlU5orwAivjE58B/6mwXTIazpYgmjPj
aBtg7VNy8DfmbYQiafy5mmNJsKy86iMO+w9sZn4XzB6aRnl/JAFsD1eI5C+zC5hc+kN5+klM2U7S
BKGYf8GustO9yanu8YA0i/kihbQdS4w0aajXGwIUjx34Pead3Kld8xam8qdQA/Hs7smNElDqHrcw
uQIjf9RKkd4MDPK6P5F8zICzCMLwJeswwbpSWFR/EACaSKmhoo6XTt4CLleTmbfi98pDo0dyo6dS
K7AUGOZ4plU1IAHCplgDfWfly9A531oF523U1CsPnq+jXl/UUmUvy2Dl5SBH4aPgo8r17bW9/y8w
VbTpge7CmUyQrKR0+JFSqEJzoYnHCPEJKB+F1QD1F25NxECGvmGv0Dfc0FkOO7uBlc62xEznwrgg
2wK8taEYV7uhwzEBg+OlUumxiPYlT1pK86xfiuNFsg7imQ/IKG9uKqh4s4lVhusgXMrxPMN/yN/y
m52AmOdzZeiGNU99CdDntx3+4wiUQsZIsOd8+DK1YNDwPsFzVNWb5aWAAfHkIx56zwMSRmUCkECV
HpeUjb2MoYGCCBGys+wvGQUYW/rdJPNp8cczpzNJ30AIHDTDcNNZkvf22ucnpJ4MyTI2tR3FpDlB
UvYuHPXJnESeYrlZLJ51JdasIcSrvLTW1Iv1t7Q7AauZ78ZU+6HQjL1zDIwEXMIeTMcrl2oOyO3Z
HRtxbIRhlmEqx33F8S8SBCvnq9MQfO23X8Y5Iysw3LH/y/Ehz9ZtO4RcJnXRmK6tCTMcogwv2LnZ
whut5EWXxWwoiJjiVbQtPwXWP5sb/aUDP8Xxsa6UI3mlWbiZwBmk68al0Oh3BOfvqEIjFrTEi5NJ
kM1vf9LjJfxahhnrh+kQWd82CJhG7cHpL/SiiOvabMAnqhV94WFtlW+lJ6hsc7RvapSosDe3PQ9z
jXO+9YfdZ9KgHQGhr7TjAqoMqseWAg7I9+5gtUbnISa9HNbdGNw02IHXEQI8oCQzjIe0YSmprC/J
o0uUIruYRRwwBzdOPmktrqx3xwC6nVieEEBiZ3lEs1AAdvTCAeU9FJGbBmsvpZdkPSNOnVe91Gxb
DisoRrJJM4L9tNhewRv6/69t8dx7i7riy98e5H4aMPkKdByI34qLK8ZchuLjwhFWC3Dq1PiG6Gtw
mR8rXetv8jKL8KHPVXGjaLGMazWo9pTExZIvdxtaaFyJzg9LkT/jt4y8XshHI1HbAWDwzGZIeYrl
rtGzFMi3+holy/pfzi69SPDTWhY/YaD+wdFY6ISBhZQOdKNjX01xvRHJvS480ChBquKCfddAkGRD
s0evp+E2Xm6D4B9CcM1gxQ9QN2IMIoZZ4qZz+Y1qJJzmAnxnkdjlEgf9NkUGk7H66yLLdqohx0EU
bWduVDZHc0njC3jxfe3IYsDIYQ8/uab4aum8Z5fCw7HGK+97Aogcnmw91TJWYIpE0aRhcQJpBgBP
gGfua655WHJfXFIVczoECilXV5uuQYx3d6iXj3sB9+bmB+V+5IsBI8rkpVSMq2H7ZvO/oX3qJWsg
MmJss4Tz//DgdNP6eRXpmSNnM6gHTogWZbqrD4Ch7IOSehkWzjweSjY/gg+7vxlzDShYn1ULYbAv
G5nugh0GOusuQSMLNK9Eik/ieAZsLDkb6HPBKluW7ObiWjz/BYZ/6riVlcmXy+YPDylaGYgUI6NG
HWh/k/BvEmdxGLY0AinT2pxmMeXzV05AouzrHAdiOrPgVQDed59pAC9XGyAO0jGjJnd2wjVQtoFe
TyhIPjS6zubzIf3OHtNbBFmk7EKQG1eMlRJ1M6j4TRVfN8SqXo4HWWBSV0es9TaxDn7WHIPIi0zV
of99Mn86gtVWdmNsyLdwlk3im9v/fJs14LtnmAXFGpTHMXKiSYixqbgbWru1Xw0U9vg/HctaK37q
xUFVNvHYgSlhuNITgEKTWHApcPAPWJ7iwFW+zsz2QpFiWzEVg5jUjR4dayFH5s4zJHoZhW7LINpM
THbzfGuH8fLg6DYzpmKykjH1cOWYR7MyWYqEXkXjl2jAj/KiGBWoIbFZ9JYtzheeCSbp1yRReS1e
3NO74c2hGaT9EN7IBcggVW+JLPkpgijIFQNRGI7sj0XVUEyUmBshw3vAVVoX7HhNDX6wGp1al1Sp
n9oYYk3ues97scSjIqQvY2mJzTpPwopNVSXVilKGg60C1Tvtylc8iZL+NQhtaHobnH8/yq4hF0+K
v28MQrQolvFrYF3aGHerrGqL+c1qtQRXBK1BKg6BkG4LAHaYJcWBfvvtGpJzznsTHutD5fSrBL/T
sqRmpZqMHoHk5C08JccpUyvYrs7cQK0p2zX6HoTDy8MZe02C8W3qTQm53lZXbuGd95rDwTD47I00
wVhJlOpssOip2xhvjWEzEWxS09SwjJ56A6etl4xN73/f9aMAs8tUcFaZAPLcobb3ZrtgXDcCFPnf
TcENEQXKQCilPV307MOO4Uneit7LtkFqZOlb6jg0Hv3B2gVGVTw3UyjsOkYoAqS8r8THIdQCNTzJ
j4H2aLgGM+h1vjjQwZKcxhYJyi9hLWpVq2NjK8bzE1coVmHr2lhRhe0iX8wV8mwbv+CG1UOdBi4J
Y8yFrW6oQs2WBrlSXbXwJhiV7KW1B+Hn6H/CW56wiocvQhJLYkgTGUCFkXmgCfXjEYDun91cYnyK
ppyizVs0EKkRg2YwL3fwEgnJ/wEoPIJm6M5ZW6l39W8ngmemazYjjl6NzBBCCRwUsqGS0IavirTp
09g7XDMJNiQaRF20kinlgUgCGoTQJqYsXPWJMiDx6raB7/7+XTlKePlovyAxGqmMCgmtEPkhLPr8
JBDSs8/r8f1r+Dos0IwRHUekRM6UUXPGCwWrf02VGwcJMm7pcoNCTQxlwp6WlzY4B43QOVHyzch2
mGf9tgztNFHxfceNFvutPpyKxMarSGFtXq7fNdttoVEt1EHNzQIu3sL/EPuGA0u7jO7UJ+O6Sm3U
p9fwQHA6PfwSumj40aEHbOubKMXpxdOszb7gbSRPPsr11LN910A/+vt6B/+LC8shtZQZVTG9oRSB
QeoWIloymx7Dztd+DMwWBqms+zhrOetcEZRKQ2eIRxWdZYXvXuE3PvHtF7K9ybQGJ5cu+mZ9bNes
/K+Wt0pFfIhM+OD3xn/QvANlTUB9Kq4JOrIBcJqLj/z41fBg3ITg62rn/i+znYRxV5gQq6CchKdh
rA7ss/LdTzgP/JxDB35TI3H1Zj0kWKtd1bvsR+Bc6FQ7HCMaU1dQ/cS28lqXCB7YN7vrLKUw9+jy
W3ustr4y0UyWY3nejd/Fhsd3mc2ZdviuIVQ29D5nSgvEkBhiIRjTk1FlcMic9Z0jHfznaPHPLewJ
2BFbXKzAfj8drOqkQBIHd5m6JJwrckwb2/rFJBUhp17H0a89bK9t/wOLnWNtXLyC9S7btNxEqrIw
DSeGZygkbkRHgvcYVduO19nTFpmHlMIetQN/QYLW1MoXN0TyjWv0Kzn868rOFuiS4zI1zZYT3ocY
BawHytkvMokUSNvIzBEM2l5ZmWUMv5LArY6H8U5ySDtFe/srPTh9Glv/G8+K5HvVDc38uoKDiLrf
VaDw0uhMermiAnB6sHFk2ayRVB98k5Recw9FlN+uFcUCzCFo1b/jNVDUISKD/I+w+gywvcDTCKd3
hadI4ZdroWGMR4htGl8dLCxx3zHfi1Rk8Z1kmzVXb2Ue1kcWopGdX8bTaVprZy8bIFqTyoR/ScaZ
GIinS3b+tReOV3rrmGsaCmTAiRAS+02HG1ow8xG92Ax7DPtyJOwjUyzBIc5MWTJq2Y3TTQqi/U19
Z/H/oIEyECe3HzLpuXHxBTjBnkwFrJZboorRRWIy7+KTWW2o4lsXY6LYfcwVZWZFWricqBkq9PEj
tCcf42Sj+b5sg4RSDiAvQWS3iRhXC2UCmkPQAdsuuaqpjHIN8mftq/ROylZT0LmmEuLNANWycFFp
uN2sGIbRN8LMz3FHwsQ6NNbgd9r9m3meVNXSWrAwhR22C7mJBnntsf/ZtM2RfB/S9bIEKa/q4tJc
EX4+2LaVkyeXvqnqYtkzqkvmqY5/jNLT1yTC5G+dCDfErglcERg4PVjhMSlKzS4u0S1rdBtEfzuV
C/9M9EFtDdSg/nJlcVfn0pGbNk1Re42z9FeJMvQUDTeO1UyGj+Sahvwgy7phf9vETI5nBhVOUlyR
qcmncgyye/GmZcKZtpUFJsg22WvMaPZRe6f+TK3owiw30BfmKMH3oVnsvtDjAsmEWAddw/fS/w1C
lVQgh7DK+Knc6ohi8l04wmIKKFWsa784g0K6DgoS3wD6W1b+dN+ace4rCjIEeFu0CzxA4yOYuZuZ
T6MJKCShpaXRHK7Uzm0avnr+0/ZxvFJ4X7yyR0Ot0puSV6W3L0LpB/ZnkWDscuBQ9FXNcWzZylAQ
4ICzp1BFtDixnvn3ddp3tSmhw4JzZAspPkpUVvmEma6PBvX4EfLq3UsJhwyMVd3NSY4g9/OL1WW8
0qEKsOSu70q/rWzIHJ/qMput1msuCdWf33Kq8LQGbgiAoPfFzet8z9+Je9FZ+lXo+FF/5EdGs4Qv
M6f8nBsZ0vVLhPUur9gvWQZDW5RqNrJ8FQJ3dua9qRYdeNSsq6MvnBYiBiAqr7B7aavDVEFqppAH
NpCK5OPPjukwXAirFMu0GE6znguIhfHh0FN+ZkWlaEzIBBf9pbm7HI8Lb7ZWYC18nSzNsnMh7qpc
KHdbpOMGOuAA9RwhPV6dcCHuMfTBSc3Lxs+dCz3yujcXJWzGVEHcDzGsCiLMgw7KE+pHi9Y/3uKA
TckY0WQlk8083MS6Gz/5cUrPEN02pdT9D02H0UbYH+nF4tVAKx5hguRsBE1fhV957VC+hj7QwmEG
WWvxHdHoNXmqVk/450kv5/hlhiDMGuUmxA138aVQE0Gn4P7NSxaFifa1Vl5f/Dd2GY8yFOePgMpl
9kq14VcBIcJQSATT1aXKHuu0ueTa/JLbKa1j0yBTjSUl1KaClonunzRY3wq5X+Cj4hyUsKzEYhB2
9X5gTNTDQuSM+nZNAjS2ob8ZZ7IZXGUjqlhkAMeumFShxqWghgGE4auHNbfqZSKFYn+0wExjsUKN
lVNETnd4h2QJ6E/q3pcBzHkjRl6wBSDFvpd0i448vRyPCWdo2HEy2oa6CLNZreMQWFp9YJYG4nSe
HFGKL366AsN9cH7eZPrW9A9Iyx3pYpM87Nl8CG7z19g/wzKEYlCBF7e1hx/rg1G6L3E9HfxfDwBK
sLTUohD+sKrK2DElZrTmVqiqZTQ8RZhi950FWI8Nh6AZCQhDaxBTcOE0fTIAu86JxD7LenKRNsTl
LXYypTqL67QHZ8RaTlLVmXoh2KDAkGePpW/GzgOW+ZXSC4G7d3PcDysYklDneQusCYn1N8W4o0WH
jZoG+N8J9JBhCcbaI0XKk8s73mb50Be/BMp3h85md4VGBubd0kpKxKgPEvJNdHbDv0XyACyoXy2n
33TjWHMv25rwy5OI7MQXJmp4TdB3OnHdy/s/Iwrsm0BJNa40f2nRREiV829csHNZ7VGXT2a7sFad
Omm/cqNX83Jb0cyeP6XMo4yA2HK+WK1r7ewLt/fEhvMtWpxC/ibfEIgT2tBI6Ip1ntwOGrozAdYF
UmhDyxPviSX0YMMwcqHpJyPw4LIJp/u9jsBukCQnoqvTOKShCCFghSJV4TMAnVE4hSytzjK5bkao
L9YL2r2YzOeHjkIQMfGM+qpsugHj9vA+nCs7y7+ioZKACA/heCSXi2tLXGfphcW4RgP5M/DtNo4G
6iXElZxUo+kKmL67CopjIV2NjwOyLPzqZ4Z+R4AVDOooZ8qWh4j0A+j0Kzb93mCVBT2v5t5DRtie
r1g6C7VW1oFGgZEOySulu2DUnI/85oyw7MoKB9IYG8WMzD5S4u525u395+LOYwW3+xlLE8B8IUQB
lUUYa28DIC0E6CPdd8sdWeIlRf3p1UVzE7Cb3UxIW5k06tQA9BykihTGPKHGl2axVkqA3cnr3mxA
yBrd9d8R2fveoUItlWItXGpj3IVyoCBkb2CEbGqZR0fRtGRMeM/3KmXHxmuiQbr67hmbwRKh4BgL
88ilbEIhBc7Lig13+zkwKtfbCI0/nAKcU3xGkvClOM/qDqR8dYHipbTj4wKnWddgc6JyVkwATzPq
STwMX74Hirx8yQ5H2muKn2o7iycXeq2qBiy6WnKnR3nMVSmm0QIWNpt4pDjqku6jEfZe3Mic5Q1D
SaDnbgTEMJLQ6IWZEyeXgZJNX++FuuY0aTLsgMgr4dCSUfb9NnD7w7QuaL/MkIC2/Ab5igtkODEb
Z+nk4QIRUWp7Gbwqu8X1Cus1k6rGXaJeyzQM9YSt3W1BNRhHE0m2ifE0hJFzQKc8w+rjoMYwKBtq
itT1uliAM37VTAO1UwPrDuBYu9MRqjz3opuJ7ubgXiQKRp0l6AkQ4xyz3HmJJhdHkcmdcZ2IVVLM
lCk1UpVt/K0Uzy1wz9KXt9ytNCEdNVloo1mtLhGLb0QUxSQtwzjNrv+lbu9p3xiAFziRz+ywFAcU
JwKz8/nE/hsDLMfqqP56ehPxx4K5cir9oTUhzvLr2WKVd+qJdZGq39PGEb4e+8J3uM9iRHERhpUU
VItjhlv6OOfXrX1Twek+qE8EFN2VQmn1zLLNvEulIfr1JcqNej4Yb4RSrvp/ePJhQF/+8meA81Ob
P0cPcLIExZn0S/RTKDFzHAd5yl/roogtfK/f3ZoaEftdGKjK5Oaclo7L/cwXsxJEbm7UJcZSst1A
5jt1Pu51Gt3YWsn8w0rAQNxYFtS/rqtOXf3rfy9qrznysZHJj5Q4ZNI9mnvBiqHLFdTgBj+fZwQY
LC+L8z/wm5mwiuRaI8RFUA0UfmjDFLOtrJd8BqfXCd3qoKqRS210e+zuJkWL16qEkDifYo+/cM88
3Xo6g/o5bMcLkwcZ6qxWbC9GuhPtPQnV4dMrTrJaaDVg2PBW7tWCTtgRp5g6Br9oaFWQVDxctki8
YUfyzJKcg7eDnyAwIcpiLz5zCg9TiwLc6PUbGdjPin/x0Vkqm5FJ8TEVs1epnhQ3A3nr2kGS476z
PQgfi8EcokffUZYNkoN9sY6uvnJDK/IDN2GS0CRX8VSWT5lQFA5hUXbrVP0UefUQpGb7ldiIMRtv
n1i90ll3ul36oPktnV8S+p+feMXQu4rYDrQATFtH/KiHVxzS0BxKBbPTiJ74T304uLxY/MdGU+LS
mXlitFhgoN1XVF9dQSKMV6qVQaIKFqJCpnPC2p5iXzowgnshWOyxIoNW6dOmah9NbplGV1IpNlqP
BYEgxslJVLMwWye3V/qjBWlH4CgVfP0FnP3UCDH4OEhnTVM6DnAXVjrVj+ZJkITaY0RQRyMUG7a1
q2Wyg5v00crR7w0QdiQJk58R+Dd+e+YmShVCEKeinQnfZTKR0bZX1AZCZlvB6dILYER/02FYXJ5o
PhmOchrY5XbRQ1l2Ep+9dt/BJBoYXE/zCwINdfiXgF4vJtaOFQeQTbjWGEdxyTOd7ZrsGKtXpnQO
BiQE27klYKAZRpt03txsgJ0Pe05xDK1qcq4pK2vz9xcM8t/NrzDle2V15Q9Qf6w3OLeZxET89Pfi
S3WfgTNBJQrvA1fC/xejQPDKIOFOXNdIRYXnW6R+jX9+V3c4sZnl4H+mJnKy7TY7yR5ZE3ppeuFZ
xVgH9za7TNK3pQ3ZEyaOg4eTwB3SRnpVrm21uUu2TOn/uj4vDWpcNnYb9s5WTstDcUcvc3RJD5Ml
GFJt3RqH2YdCiKJ+DcU2rfs1T90M6aBnrbR9dhtCuh14xKrweGFAmwXuQZUbrF5fx6L3b+mC6FXA
hMYs/llP/B0ZXAN3Fg6ECFgQ1MWvtuBdHhYGfvg1NxuwPGNOBDdhN+eEwZZEn4k2Z3P0r3wAY877
Uzjg8l3VcW5TOQ0eVlbxaavrA8LW2PEZxRYjVeRne5bfvL5n8sbPpVkv/L4LSS6OeWOktRhV5wtN
CGoL8PNojW24Jn51TiYgCwnqnl6aI/Ci5o23cDmDGmTIE0RnbbEM5ag3o11v9eJ3+D0M+ad9Gc6B
/VOfspwg12xuJk5mazx5EhI0qgfRu8PqIK9aU7JGIvrKyqScJ7yV/lKlniYtnpAQsTVoyLOjUlhk
IWxPJa/nJaLFGDKagGlmWtt/jqXcXgWZ9sfZInRZAYJ3/wbbwfULD54Ce6+dIBTE1M3Hlrt+eoij
FDuXVeEboJXyIO0kS/mO+J4wSvlbrglXRu5bQyphshz2uKGxOnNMGWqxDcULBw6NFILqnROMkLot
d2gUCawctLSP87h334B4LYCG2NL22IlyAGN7B5thKC197IQdr4rb/WAspdR5aMPmlf9LaltJjN4m
P0emL6xB5xhY8HVOdwFwW46JTZdy3awN4YT4iuf0W3vzo5hO2I80ut6kQeiS29vQhG3WhaLczlmb
aO+LTX2B6J5yWkBe4XxjxSvDNfX5q2sonAU94fftYxP+5d2Oki5BFW36Xywy25q0DLkgMnpIQCc/
v5XydWoZP03m9TuBh7lLFOykn5N4BO2tsN5UUB2Wv9maF9RopC/hIaMkjlcH8IN5306Oi53bXGR2
G3+RYJc0D2Q8iXPYxebqzCpI8887C/KavUIToOZENWZ+iyHB9TTMLIvJgMWZIErKcPTqwQtB/A4j
ehAC6g3HQzJ6Xsnjk3uxmenmVNhVgA34GvIt+jpWWPM/2S2Vmsm1556kgJUq/wpzqFcpB9rw5Q+K
8mnzEglUrN8MwT+wXLajg/jMtxb/m5TdeYTmPJwTc2kME+ngQExma3ZLsR3PzwsmFE4zriZPdQKh
I3pH4tCXtTUBhuzCHZOQKOSaZ35/wMcbRhrHyitoonzDBnRLKCxgPMTCAkFTsf6oWy/LGVol/TIb
Fv9aOtPICPo79VqG2DOcZu4WAJJtg9JlZcgzYNjSMSYE/Yuj1OoK17urwAd3U7b2ZY72YwDAqqSU
mCPHb310IBTVQ4v8YQGEmqn4xwHo6RIOaoF0BBvZO2Y6e5ClpnqedY3etr/+qli/7NYZNmUcQ4Hm
CfNbWaopUSI8f/uuwu5d43FxGKs2+RXKRseV0VSxf8VV8WTMmWOm9cKjmTNqhHgWe9jJAn8D7fOR
0UNWcg6YjjNGo9cnQcUEtnKTkqLRKA9unPk3KSW+Tv3j1mZlj3qF/MdceCQ4DKR3VIdQqzqrjBns
hDzo8FgCUv4GTUaZAy9gyrEfmEWCeEyFrCpy1MLn8TsELssPMEhyPTbLPDgZwqvW2Rg0j5oL6Um9
XzNUd+WmZrNDNxF1TKjZn7SfvJJ17I5Za51v6zAxUBWubtsXeU3JIvUmsJ9JBf2fzj+Mbo9jRdR3
5tX0a+sLQYVrk6p2V2dkfv70BOLwsU6kTwUpAk7bsokFcJFn/8xjREP+ZlfwAQf5F/3DDnuPSrIx
ZXgK+GWukQ/0d8DnPSoRrDU5cVvZkF1MlggdaIcaJLQhpftFekoaTJywvpjWdsRWOkjCn6wMUg6J
/fQ2ws07VpKryPgFwTdFM+4JCQPnW9l/mUwsuwaRwdXGiW8fdy9w7Rv2bQ8iW2Xv1vQv+ZjkpnQa
z3icNsWd+RrANoxYm10mI3ku9cRIRlGbPRyhvd4M55i0HwhOXWCxSrH5kBt++sXvT+Wz2nISZhbq
Y6vCd8DwzJDb0/MMrwdAgKjqEo0Y3aRNF8M6LA2fBct0/6taf/+S6Z6u7KrGJGrT51MRWACSprSk
/M43lL4WC9+iq57gSNYaGQmgNcaFl9rmkPPYxplZbPq59JpH7bMvUc5dCk7QAykDTwb5rsMmIz/D
xfjqFP8EM2ScJCpcuNssK9c1vsT2RouLzjJNsI8AvGlhyAK+4tFpfr2C6jdl4EPNnUqMrsckqE4K
dSzuQrGyDsYxB6FxJ7QsusMXRDQ/bFz6CYg6LjD0jHrbZk6O1pLxqHzEPQVQ+Jch1/F5UqQnjQdf
1Cw70DqKW4uiQc8fkS87z8UZzj1bPMpdk4vEEzsXgKuGpiAz5ACOizk5BzR2d3BOOTek/XitklbH
Unp4oKHy7VWAx6zh0hne3yXJu19F9Uoygkuxlen7fFlcUK9XBWOgAOuVQJVU6Y6wXfXY8bsfEHsl
lAOpXUJq3tJjtPiBRycjI+0v/T+MTfjM9Jdn4kOf1YvTZz2saVgSQIlu/hUKCiSBFRv0pCVg6oIe
PhYZDhKjrOl7fF3XhdFnn1MQ+dbuqQ72vkIiurVo34l1b1ZXu6iC9FM4NBJIRNwkQfi7yjW0Czc3
YE0LtZB0fEYDa+rjO4n1JWPgRm+mnb1rnAGFL11AzVXZC2JOeHvRS1lLialAQvt+IdWPjp4I6zcL
HMWWu/9lSsFT+I58GlNf3Agqfry6HzyXtDFcFwOKcZz7krnR9JbJ1A9B6p21INyarTqcfNEveYzX
4U/K3uFFhXG4FuMQiD4H/iwvvedOsIEnR6FaqSDVUo+Iq6AbVR1VjpzN0aTySVjD4fENmSzEcE1O
kfOcOLVmnElwI3AfaDXv7Rb8K+fO97cdv93gDdZj9RTpMiwqOjLeBlTpK4EWi9PKnKt1jkC4DylV
KRpVrHS1ModLoJKe2sZhmatRg+4shM2IXSA5g4u5V5AcptsN4OykNl/08k0dNvPJEjgLffZALw7l
Ja2eZHU9bRQvwNk6fIZJz+s/qOKeDLHIn089jsLH7aPKbFcoOB5VU808HafWjtkllwaiQ/5q94Wh
ALpQ75mqWl5K0aBfPJVTDjPGhfK79VCYrpewIKtR0YmlVG0jNvjiV17IHef/BvHbTMQhyDjf93yj
1xdBwSiLLoOw4E6me0hxK+N/BhoQ2EWRrBApmEg1A5EaWnPBOif1Amkfd1xhSfOs/HhODt3l2LmQ
WYbmYdi+uwfZcoCxwvkVtnEQtApM1hqL8+QlmGlouiKgFRcyePUtQd1/ZEisAQVGaShNJwi9tFzI
qI1EYXPj/nQhFvvSbH5mfRqk/T2Z0BSfpG7c9dnzH1XfXqNz5tzmgwFwEA8Ij5mlK+DhfJffzVaP
D3FC0+x/kCClPEjvzJLFr7VXKUP27zXJ34Z66RlmihGV+ptmhBxJqYSlyhDKYprkGI4kn1hd9aZF
L4pcKOhuqVPjBHpxW35EP/st0mWXBBJoZ+klVKD/6mu5x5NMMbXqd9nc1yFtaHCRHTwLi5LNRp3w
nzNe9RcpMhAoZ5EXpBXbRoQkSP5HrdRxA55lQb5v3+VAnAn/3BFBQSEYRQe4z20nkAimfKUOWFn4
VxJiLpLRcP7VJow6Uz7nxrGRU5F9BngkKCODWTrBQIKIEsjj3fq+b68RTYDC2tBBp+IyxoglL+D+
uSkObeeXaOz3GmzPI0bBtvesd62nKxAaRlulwqCUTcjgpqcz/y9sXT0mfCtHS01IKdkW2k3xKlpY
5u31KmRXjLN49axlmSqPpZlHoBu7YsDSuJS47buWGgoP/F3q+J6rHW+RswfoKocp8JqkyxNYZTP+
fKr5nRJs+idADmE0MpoQtAm0YjXl6d3s5Z+Q1l50lzkkJa1lUAtJFwGYu89BP+ClTnEGfy676Q8L
4SfTLAqVlKAMCIeGBz0AFh2dtgnVvi1+jg4DdJbQABpGOIgl2IOW3/EnrtvRSQV9R8qBcGwdQnxl
tFaWM01Er9MPWRFYVUSFN+M4WvuoiDPPl/sN/iveHm3nTcKgoUEHHe2KFHe6MZtUP6LDqvPePh5h
EZaJSYtqc2m+NwWb3yvSkRmkJO7YUa3uqZ5kVHQrAyAKkNacQmdSkMoB6kEcETVnmOGMbYA9fyQ2
Ya3/o1ledHJUaBiWdXlw6GxjjG1JX8z/5jQAdefWb6ftolMJXG7rr8AfBn6pneTrakItVe2u1Tdw
64hdO5aEgXyZd2yCQcXoBhteKoqnWSNS7qWaYPXDcuwhi9mBlrhFrFPApi2b195qbez1R/i21hKb
3gymaivC0ZSDmT580i0IMl/Wp0zhfXmTpOBWgfEhA9EH1cNG1j+tSGeLUodVlzXZNGgP5UybbU+d
95qr2HJjo2Edrm7cUStbt3MejHN+Rn7AJWMWiZHnKHllmRXVtXZ8tJ01M0yx1KbKrME0PEcSrcqA
UQrRApL6lGSb1XV70Bl6n9ziImojpoW4ntaxfjTrAWV/8F1sSAmiDsLUEoooTnVlsKRJuPfxYL+A
qRjyyE2EogDh7X7v/S+51p1SNOKMhKKH44b4xfmlx61NVR7Nq5wN/vCKyE4QRlnjdHaiNu2arwLD
oEgfe9wh5s27mmxyixkFXIH9+nVWSVWA0p8Fc7ENcV9ORUgb8R6z3xAVpl0m5c485J8NyFjXgke5
W/8PqIFAmBABPQPSHScLAy8BBBWCCUZNMr4z8H9v+18ECy/HU/JODyvnGp94XvjQtYxmtZ5eDpcb
suHhzB+ZUrw8rU99XjBrmR1QgQd60+KqTWE95F+IvPqRXRY6rTUWc8sfwvL6RqXSsnXXvTIBtNL6
VYCtimuX7E/mkKMIOWWQMIwvQtHHoC74dhn612vzrPEhRlW3PpgJXUGthal27Fv1ctmAHEsfKYbb
pscwGKHFQuhElu1064ErS6kTQdQtGX1IW/B6kN6iXEt1ykWACOqTnEpJ2SC3m1pyuKU3etygjOBj
Fx8+9ef3mnyPub48Vlt4bVhpwSnf05lUMEQIoi6Td4RGO5wdqweMpxFnFCfsExUaqBbe98Stho9s
ljGyeYK6JCF9OA427WWxaTUm+mHAUSZLaouvYXMP+1WeYdknbDnc0NR1CQWHTolvDHiDKe75NzSV
OYBRF9jBKCVJegExdv/ixUaZOBWSFZnoZh8XfAQStnZi/2BvJqWNVIvfPbY3bQGLH5pRTYsERpZm
0NGVZ2Ua1ULii4+Nxz43skDPZiizysEpjJjg37vyCt8wkZep++PQ4wGkcmvl125iILjDIp/gwtyA
OIidg7qB3AlkdeP3cESPHOsQ04YD7flvvQKaQMi4WSdkON96MpzpftFo6NipFJfhg92RPGu72Sq0
keU+sfJ/be86/zATj/tiWDOTG1F/dlr5gv9gMxJDZHvAPuZylNsi6d1ZS5ZbdkC4tX2E5/R62dBx
xJutP9PByvOV7TXaF8UzVGkDipr2hkl+392p+EUmdE3UDQvV8PkrNjsAEmp2ljdv4XuUEN4sMq4A
oAruBMSvQudCInghQIaOXC9VTX75bycDGexa+OBn+iMEO6h0s9w6v+3n61SxTdSR7nAkzhcCJL1B
IKklop0UdIr+IAmlamAG0tdfySA7RLZZp0KTiBwlFOFyqq2bz7azQ6J+FXPHRsS/daDYSWDCnF3v
Ckh8e4ymoJXffib9+Illnt5+RUgQABzLKRrAFVksBM8sLjLu+wQ9xCSPAce2ORxbyJWW66R2Nnv7
6g2A5eesDwiFdU1hfBqLQG1AMJl00KY+CLZdT3fJKOBnIaSVCKy9PEGVHQSuObgplveDbB+qfhEQ
buWsEWIoLp2jc+5ZXeZ32yXzOM1DxVjt5ueZ/MgX4AoyURTZf8/PsD7hthvbYPwKv17u3GY2WT2u
YZ4v7Ob8gPBUW5sxUYNF3jhSUahbrTrCtWUu9ZF1Zl5DLmej1PwjTET0B+s2iDUiFNfsN8mQJDIB
m7rR4Xe+rJE3CGrHcEpPcWJytDHbXMajfBe+it/HpYxTdfiBbavEKbzr97uxx0POaKVfVesXOJnS
Lek7be6r2qFEW6DLPk7pjr3IYODLRW9sorqBcpYWZCMQLDSLx7UvYOPLHR3aYpOebLhQDF1GsnuJ
0zTmmkCGG7QrIA4uC6wsehPnDanuKWTKKYw+IY5RLkuWdm6ThekOkdZb5igGaKY/yXNoXolql4Jh
3DmTNxMnh7+zzzKlzetI6nTyhVjw7aFY7g5tNU3KWgol2zDpnaG9uukPqRjsn6aObQ3oSDDVWCoi
HiCYg0s/OluYaWF3fRxyFXp+YT6tmpWsuH9wvdAvGlxnmNvOT5k3sxhMJyfOqimWFUwACuUOTTp5
mVOIGkMNJ7a5sxh05+XTl1WJVx8NvSd8dJeyfNSIsI4ri/Aif1b8Jt4W1YC9NYGrgOlsrTCYgiV2
4G17y5cjBWefGlJEXLPNl8A2DwFqHOQndqO9ev7Deh/otRqCtLMB6VmFNC9KMDPrO+bODW5sw7pW
wMJ9wXhyr/zxIqVTp3cszN+tS31PYStSb298pomWPtMuTHHziqnNH1X4QT3dO/F2pAPJNxoloiR4
ivVxPPPHNq9hwEMQpWDODPWFAP/OF1CeXipVFP52BNop06LDAf2raUxYV8B9W+Jgt2p2QVNNGj3N
+Tn46/NbB68g7pFGYFRzIfJV4swqqcMox7EEAdyptGNjQHdOEIQ8r6O6LJFyECBZcfVVKcXP+WlB
qMpTeU9jGGH06kDZgNfUu3Uc96gDPvZd6XmugDoJKXWojAiqxiUWjTSLdKmjfkhi9dSIZcTs2GwL
HR8JfQSMw0AD0bXCIJ8jVuoIUk1uuOHfBKpvvA2snlo0hpDiPkeV8O8TgsHaEmMYUHhKoQB+HDdT
U5n5DGqk6GT6ja5wyhe1AB1Nxmn+98Ar6zow136Mf4xHhADhc2Idwlv6kFKwI9Mjb/NVGHFpVYNn
B8ew3An2KrVO8w3bUfzcBM+1IIES1s8bnx3Zx2ofli6Gjg6TaJ85I/u8ZUdI6Y5gBKeahFk9D+VG
DUY5+zgtWDupxAvslZAP3FpCL9+dd3jYLu0f/qRdPea3ypyj6dRgnf0daaqU5AxLJO1uwJZYudxd
VwoTRW5mYZ1bkS9FUhgaavYVkEGJweW8iqlcHbFbflTL3NGRuOG2h2DVBAf3Z1EaC+qOvLs0EVLb
kijgFV4xR9GNJrTPNqyEWO5Q0lNjSRWYt5/buHXrqoWYa4V2fZSmnIEjM99bVr+KFEs5h5KNLkBM
FZVr7P0hhV9Lvjr9U5w7IIUSC1kXTKFx/d95EYgpkU8uc6580cp29bFIa25uiD1rg5JuBMnCxLDd
SpucnByGvdMaVxA1x2tSZzQkyJdnMfgC8iyLHKxtN0mvIePXfNyAWMrH40XwrNyo0owLPjMVrehs
hGmi7yqH81j2bgxmyf+dBo9fyZKmbz/Hd6VUkpqjKzr+k87Plm6ID7R2qXzM7u3EGpOYpJlOUynr
B6PjyW66TcKvq1oY0lqrarV+Z2/Trv0LureAC8QFemzLaLwpEsWYAgdWx8M/XS7aXYBRqvkYIVS6
n3TFnQJCyZpHF+fk3ltlwyUoHZP8Oos9UDcKQCTEtsszNqkJgGoMEc4C2KEYQtRy5riOPVe0KSgp
ZGDQToQFOXsK1EAfaSc5zv+9d2uDVQdDDo0V/4oXmnn4jp8arEvo0BKfAcElW2FtNm3MFRqaCGu9
jhJ+JICLpif8tifQXsreTXo+mM8Faq24xH90wQNBlWvJkTCeAOg2gylaWAK50pC7F1i0bGl7snBn
LHG+U/WZihqslPMEUKZ4nLo6k56eoTYEekVwvxD/9RZS7lZwZXsa58gFLh7ymq2Tw347ptZIMGUG
XlZ8zCad6pW2kejEqLByAc1+IY9ZyyrSqv4DuvQC27BsJYuECSkPAV7clyFc+hWwbe9jtihPBiP6
OCmvDdFiFIQpFxJO7cwR+BSdePHcyteQmAhkNnGpw+SEDhHDQyumYWfiQLffv7iNGmWcbM1fZtK2
LOw0B0Nhgey3JM/mMGYPfkV6dYM+Yty1+VjgDlU9+wpsWEvE8tSg4HRpOIl/WVgijrsE8gPIiPTL
jmWIrA8mygDaYY23MjdO9gUz0dyKKheb710ee2n8zD6nlgAL8BU+C4Bg43UNK1YXTGuqYzbqil7r
qixymLKm2ioqYD7hTT/C39d4/9xNWILR0ZnIcvRdR++30IO6Bz7ySZ6gfyIVycWtyrnKLTpsXiBS
bI6HAr2pYoZALbrON+W04z03RaobDYHFPMSNyzjXb457IOqVx7VDMjya5ZAQkRX7T3+/9l0BLh3y
CtzIGROF3qTRA+8TEom7RZTUZxDIP/SE6vOncFSGjE1wwM9557TlDOQrAMY1dftm/qz+2Ku6s4DO
PUch0x47y/NxWj/4APly5rMdcXt7tAns+IPXIrHnfgrWHNsGlNCSOpzo3848UJPGhgNQ7PsYHoSt
W8ewXrDdV5EEYdj8YXiZIH1ve2tiEY4HxQcADbrHAkV7xbz/yhHgR17yOm0n3HH3Ts/2wIqVdGWE
Cz+u1xLm8EAl/iwSUKGbXblvNuAQWEz91ORPpIQEatdbfNoEoHOYiCf+dcmozi1VeWXftBZeh41g
2K1MBfuKIiiWYdakKp6xRVqoCcv8tcdbxEEFLqJV9TEKqjZFUDPehE0vha+LCBruul+WVCkyJGxR
m0xgiNxzmGdOXEyicfmTz7wja1mqTHSXRDrF7Zk22i6UkHDSNj5M2qykqbsuiSREcCVNYw8RUkiU
7qS3jeclHMIiN8gsq5JO9uud+ZeT0Rg4V4nyvnvDNs444dcjTBa30p5TkFJKxyaGXOB/CRZKLioB
S8HQpdBGjeobt/fsgU1vdJakNJs6HZBvRrVuSUOvzz8hKP3E4321tUtyT8yjhPO2NQNJh7Wn2yQ5
GO3Pzx/WQwaEiTcwwi1on2ajKkUhEedfhBZBSFkdnerMu0REJuYkXH12v5JdhlKpkse/O0LTym7N
+4tWypAzDhluY0Qy/5MZDXq1U4N2LagxT9181oVB7MgmMK8kFTSUQGXRUTW5IYNudKaFvW5OeyiI
ocNYt1dC6BIy1VcFTNHT9xlv0OOj9h55U58NBXwaNxp7AfLaA8z0XkvkEhWkFpN2tS4Qs4N1dE+V
Ulz1d8yTj643g5OaTtSGxGvGZTFZb1t2b4Rp/hJSQZnZ/ghFJXoWaH77Yx6xLFOLEmV8pK+ztakr
bnkwcwZGJNfQSdadTwHNldMhK3dlbUE2oDbHl8/PwLQ9oqzn/k3Q2ITt0/9IIz3PkMlSyFTjOat8
vIDhaVvX9vjb8JjwXudbU5hhHd6HOc1Fj1fzNq8nRz+A5DJYpCVj+sfNX00Tk072vnd3aNbp0war
L+Kgy/Dbzcj4phVA5WsCnreh+rwruOxhTb+9tb2up+PCmrbPaPsjFXBUZ3K92EwIeklqD/7BcyzY
+7YGC/nMM9lf9WJ1BT1hf1p5RwSN6sBy/jJqY/uHF7rul6xNaiO3bBnEPUOV0gAy1VJSnur4VH1k
2yBaRoypyOO7m3sdSZNxNgf3RcMXtaldhksF3laJv7gU09BU+qinnbt3ejTANy0+plT7p5LXzzKO
7lNgCy5eRmhvQ+OTU6CxuAM5+tqu092Qbg5qWCvjLY4Va/LcOBetVIAYHz78CTVS7yXOy6/Zchia
KlMbSkWMYIH41aamzXP/bovS07uSqFcj7kSNpT3h7SUUlnjSNTonze7v422eBq9DdP5gBFDnY/Fc
u1993kKQ6hb0U2DKnBD4FmW0rzvkFJD7NDhrWp8TTJ459fL2xtobw9WQ4t+tAPB+6LFsr2XlVXcW
cYUZvEj3VC4mguCbmRPPK/WAzzFCMRduJDtGduGI6AF8KfGG9L6SCf96gdkchzjvMdFZL2w1Oa18
yIyZPh/ni9QXxbUkaVW09U6ODn08cboRYzOwwdC1jyEfsU6w7pRj83nzOIx0MC0Rj9qp644p7fHN
IFqhFSBElsvRsCoudfdw4OJzEsMVkSLYLEqqNeU+rSn0s8TITCXFwFPj0J/NNbbPKhtxbbM19o/m
Z760BetUpOTEXULkiqY9hMdNZJzHJGltvTsgJmxA2S2X797V0bzMQJOrihThAHtPYrU58fJUYB/R
jmLBlXgHKdyOB7EcdLwtf5QXnNWEnc1kJ3yRGssdPBei77CBE2Gusbw/wf6z50cGrM71XVTOr+gN
NadpfDBxurAqzL69Lw5NMsgMlf/+D+sfbLRY3zrxRtRK3zZF6V88GtJJHTSd+lZkACVvjm/vapN7
JKIBOKIOgwuQhOeS+PGCRto8Qfa7AuhPYBTw1/a7eoozI/X7og8GOsO+MT2vZGiQV8oKodFevhyT
eBE3IL7Ey9rS5QfoFKR6VW8ly8rRU+udlVloguieNbklQIE/ql2pf1i+6cVkIou2KW6la4+StsMP
/amuNrmNX0DnSnXvXMNnDjBK5ZsuE25wkTLye95Z4L7dsBogNeOmSe6XWhdbDUE6qZLlt0B1nCxd
tCGdwCUWPQpFjmbJTkNXCqXPYyk2LoKPA3AAcQoPWFmPuwLPtrEIO/2RGrXll1aQ4TH2w71HNjTu
GO/hzMegbj3PEGA09pFML2CxkbYdxbXTFJsAmAHhWopwdHvAN4Dj/tqFHw0DyQGvpE4UX5BvLZCB
RyQIBW3sEogL6C9er0HcFxZ3Hj7jMED7YLXFCB3CBf9f7lGRRS23X2wNOnMK7W/imc3KKDLj8Yui
Rh7TlfXcX9P8FYFewZxBM1Z0vZICzX6tRwcEX9rBIm8sc5r1vGAJVigha5q+dv/hJU8ErTMkNztM
5M4Yt/9c2TWyJYyI/Bbvi093P9+pszyxWfyuotAX0/dt63ghmN15BLI80eQ8oaxd9Jm5BYdd4jtw
Y4/va7KebRsPv1LOCsuNaQPHkIo//VXM2o7qt1sakkenkx2GN3yZcOqjEEiKLxXahZCPfPblKRe9
qtm0CiS/YDB5NdwhU0gC8HT4vKAmrP/9Chs9XdCgRCPcJa4cxHnG5lZAftRXKp2poCCizZtOJ3bJ
pmkS8YtCdmOAXBSAfL6hBzR9bFwUOirQ8C0PRUuzaGRZzrZDcP49blJoE4mHuUqBdpFvp/FoDeLa
yWQ28vQhS+J4Vt/AUCPBWY2va1p6o1W43Ey6whqL0E26YjaCO5Roe9eJGcgQEAPT6H6M8iIMhfai
F++hkpuvdTRzNXFTnlDR0ZfmEBXrlCgI1CAQ10AfoQhodFRYFsKkE01iag/jglUr3nlpxIv5DZHA
j5r00q8rxfhaTkb7piMUUDkspBqrFCUmoQV32nHq0HRxiVmGg7Jj84SlPN55krq5jj1XdutRi9w9
pol8tbBMF/J+OgPJLK2gSLPyAYt4kxV+au8JUhwdfVDpMRXRnK0wN5xB5S25bvyXdyPPL3FX68ku
fE+80mAoKncLTGEe4HuptsJ7Mkc4rEYnfRXP5ED/OJe1AQqgv4vkfBhuiOWWoUJpkiiHgCBzwrja
ritXSN8vJDiR5Zv5IF00LkntY5EvZ17/qpMLEjd+dgIiHrTPAXR0nOvx4g1sDqE9L8LF/vZSdB02
zrVTjcE2MUyg1jYi5FYOshEvYzEab0dtkPv03bln64Ykv1tNDsc3Vwkv4Ml8ZX5reHRlKPT2huPG
eg5+s2vGyku47MUhPZWyZNgOXWPgSllbCQhzGvUNRgJv7SF+YyKVsuXiehEbKk13ApVYgWS8yhn1
Z1J09xelpLr86lb5eU7vdxAVtGKQ8vkow1IT5p0G+lotEiJEnuU3Wd18s51RuRR9MbQkBqJPPrjJ
53f0IMVf2bQYODaErPtqX1cOG5rVNMFUp91HVLFB/ndNDf0Kz9rTNKp73sIHoLPh15Qc4oZPfuDC
diRCs2dwFY1aHIt+1BP2vE7ieHWKPPgjdkXmZPNOqDH99NsYskxrCTLx7Imd0xtFUJofjsNPLtpb
zve6d7hvkP0dsoUgGMChMYsQisNlziZvIBBdYwoNUpILvX5LDorZ9sf9GDZ9XecpXL1BMyd63gg3
iNdPkpC5kJCBkCb9dXFfvNOX0Wf5ktd7H9dieFurC+eKGx4BgwVXcGoA9vtZ7/nsG3JCJFqPptTm
uLiftD26/reObnVQciC2ktOld888xNg5ZGwUagFfVX0DXdm/Mt72jeyNFV7veOtGvruXagEs/Q08
EPo+Qy/WzArCrLJ3AIhGYzH3Sn9wsv5F52JRTrsgeiBZJwi76Y3aWFnHHK8+f/CGpg0mJO/iMnkj
o7Mwo2yFN/wnVoA4WvU+nHbPvQDd4lHwHn6oeUlyiwOwhTR5hQzIWhDl+SgiU+JDtrM8QGTUEhrw
W+oI8nV7lmdimWbjKMMZ6TThzZR/fmC4QD9eRJtdapHRumNGgppbk+xhR2K6rQjUsDUJrWroKj0z
Hb6S2cLW9jMzCtwLE8nCUnG4q9mOeX59jH8h56DWEIuQKo87+psEngzDGnbbDKdHWW8Sk1IAAuEw
mxCQwyofoket4E6XG+OQOtEIm7mv3ut8V3FJFYZWErRMDeGyZ0Z9y76sr+1i3i0BEYPPhB4a1HEF
CkKwvcK4374vLm0KB+Fi9z7fv0u7UphNmAp7RdXVgWHyu9U6DXXi75kR7l+dhzKTO+WcH1ZfX43g
NAFMXNoev5KX+D9jo+HCoNyH+sKNBEkpRta8gaUiKETO67b+FwA2/PWmHpcWnXc7XTS9HN5RdsxT
z6K5hN2yJnEGpdqiIUE+2aQIPenOmNktZpAYzcbMGs4o+HSCHHW6lIfSZ+midlqLcAuQFg8exASp
RuG/JiK8NpnZeVIxldiKVlHvxE98zCC+hM+hSAqrkULhaib14owLi2plsG5cWJ+w3Nd5j7CUh+p2
iNAOGevIlvvPkoB3soFM/47uIjOGzfw9in2mVjLEoVCwWTTkI+2O0BPDhtpTzaQAu5f1m0JToqWZ
s94kqTBqL3qiPOM3NTWNysDoV+3Hk6z2Y/myCkHgfd4HTvx5kQfqAN3P6Fbmuq5RlW7QmeBCkHjR
jQLJF4mkHiJefOSfj4rUZW1n6RtdFbibQq3ZGUsQuiS5JFCJdsUB3/KOiHaCi6EHQyYtdc8Exjz6
kyvpANqYuOJhKjME4x4yOx6LCHbtkKEjBfp+fYbPQGWKUuTAPwRwb3THkcMabKYPlVSccDJaO19b
u/bezLFpq7GcHsC2fV1l0o9MmqtOqrKTY8mR5Rcz+adhxk2c5vAasDYgCDDssh8X1DdDgReaEOrq
S+Rj1ZYEob4nYtum0jVXJorli5/mSM2HlliekChPjIQeNOR0hyz2ktlyTq3bmbj1qi7dvj5Lbmao
dH7dvy8S9n5JGSM4HBb6Bia85Z9bCcCqdSRtddO7ZG+8DZXyy4zCh2SB9L3MjkrkLn4zbaYsfjrk
mfH7FxWaRAFTn6yeYdm/zulShxOY1XCaxuw5aB1c4iMuSv+8ZtzJsBV22rs5d0PrGugpdvqdPZM6
D5wbULno4NMuB+GXIrXUxlBkQFqx5VDIqlWD+ESWwtTuBOhTJHfHq1mG++wTPcmFBaxk98Dt4tHO
qdE6gbLj+5SBF3BmoMM1sewe7lVwxK4+qcwlEDGh4ve5oMsqIRCcfZFVoiGxtjhICgA7zo7suFIx
adneXw+KcniEYh6m3WcDthgsbdcLK2C/PECPNzloIEv9ME9gvF4a+lWC6xgJDWCmcw+r5BIq+VaN
ILthyKKtYJJD0RS5uzpDmabcPzMZHiYy/Gf2S19/aj3u7CVGrzXT0cZxPde8NEMH5d+YXbn6za0W
skEbqr9Tx6I3+mJZia9gdi5ZKpbC4focEQmkMS/UpRhIVk1LBgUq8CM8gdNm6V7rtjEGr9cW7HE6
YYkO7ZsvIX0jAbATnct9dEn8EztqkjWwaO2v0PmLzRDPXXzoMb+nUpeXwkeBYV9j081ujhlw9Cw3
5Nrzyn3WYGIbCuQsgpWNUMRxWpbmLUwtOpivRdaafMdxvC9yjUL0bhWrO3pl3fkXbHR3qPjN64C/
7tWXLMKs026VzPt9p5I5qdfZ5e4d3kHcoBToJkIO53lWTZOUIukvPr1M9Xw0IwR8U261AoAJa8EU
QRY7FZMNIVurs8ogqoInt6BbYnbs1fqLEIV9IkZOCQxufvHf481nJ5jY3Jt0qI2yBbBWaDNz1XjC
3lmkg71wPZSqf9fDeChu+Hbej4ukDjlSDZll8ZXIbbEq9UWeGanS48c5oBcltew0epRtI4lrGedh
3aVrjJkd1Qg3oU7oI9J++sLkEQwxFjt+W7/NNiXVjIq/EISgMCthm+wfv0lcCQH6X6Rxpe5Se2Sp
Zrceqe3GbmnPv5/lPb+GWE2Znbf5vVKk0IqyfTxk9lSVuvQh7AnxZLpFp5QS3no7pMkE9M6PAC3W
0QJIF2WSjatszrlSxwSaNq9scdIKLrXQ++8JfrearLk9cMBwi4ja/gVLKuWQl+FoqsyvbK0+kX+C
oIrMGiOMS0UfU5dpHXa8sfTNCjt4uZpr4zScXwuifPMfbHUg02pM+TvaPWUzazI0VCCzj/DiahZ4
4cRkng6GDEK0dRSmtquSm8HhaDOfOFLc7IJYEJrK6cZrlXEhbBloxX/jzUW/UFLBGWKB38eUOFM7
iJwKiue2Sl4KyRN0OR6ABx/NkpkMtbEpDwg/MlBFK+1uf9dihKhpg/GKvnWM3/NvmiBPnpGg3F+O
iO9Fjrd6d95nOD7B+dlHHtJCB3bWfCuURHxLl6q3LaprpjGTYZUhJKP31l9/DwFXTgynuSvpWVX7
rcx4l6f2DajFsbZQqEBGrjewDveFgG5td/oROcu6yqP5Ro/ghLKEMuZqW2M9j/L+QkKl/xkYtF9Q
DonsXmydpUw07EAK4zadKxmk2hif//WR/7XNHJsMsBT1a+fu5bUa3xr2QdRi1PcI8pPXo/Liyk2A
jx8vAFCEL5KiBet6qIbIux6OnPAz9qKXEVQ+IWWireVEIH3t/1YOTCD3DJEM4oc0dOHF2Rb4NaKv
kpnE5Y3kKR3CBjs7kwvMvzF+rhE+OlEtHhlOe3Jxt9ZZX1rVLhYXbkUtdhQFLzAIbhS3y3N8o5Wk
gST2oo0hWfMAx7giYhljqYu41mLiIMuyJBhMWKgKSknjiH4O731t9QbSm6hooeYLy5V9M1TH5cbV
dbnvzcuDEQdhTPnqwAgnxN1gFW53Q+AwNBsjd7fzvK0vKOHOAF3ibPrMbzaJI0ddcaEwHhoJJMLS
elSL4Wz5PDiReRSi4M9JMvrQ9+6Z3qhrdUPYSSmnmkLdwiDC7K+QIk3Vae9z85tYWdTfZR+M4zTy
hdnPgVPAhvzbPleJW2d24edW4R5ljZ8HDRsNSWjG30F1KRsqUXa/rKPsbzm/vTlbvL/30uDgK4N2
5kmLwbkMA3wsradLbVUsi6Qjwg9znB4H5Detipx7wIDvaQGglxEcRBG1ItO75I1zib+JzT5hpP8h
ZzC70LbH6vpyqvbAwKyIbdC5nW0vQNIy3MHovC9HmC9C22QmhlhXuz8jb0fPE+QsnAnuouOKj7a3
NiPE0sXlKsEEswjx90CdxuQQcIHxUYYkf5dHIGhcliDeGwKMIix9OedENmonFtt5v5tBe7yO1gCc
kfcsnlmoUx9R+ENQFXVCl4a/4e8a1Q1RsgV0qwVjLijrIQlVfAJPiSktQU2u95SHUuIZHaz5xhi3
uAp2TFYRdUnmMC8QQS7Meh5MUHMOvLCt+qTkIpDXWi5nI5LN6M5zutjCvBzldDx+LDuJHU1q+DDM
dYl89der/LpO+lwimcw5HyKafta7q3n9kpb/zeG1/10NdNiyDayOtO2j8HC+2u70467WAvy3pWho
1Q2tWreuY1CzRucE1NngT4yR9HSA1Ld/P2PSEcRFyA/E6HbwnxuZrMqj9T20e1t6QIQzvmYxA9PT
mEkXmlPUgfoYNMD6uFA18R548c//FQq7MBRzXpIT8r4AdH8ULknOIKJI9iC0ccMw1f2ARUeBiqUb
H6t+LXi9cR+bOF/jCTcPTfX4EI3pFwecspeSWjMYpssAZY9NYLYPaHC9Qz6SIVGNL/gQ3FDVItK0
bNxRs1XnLWhUaY6F4idjdyPJKL4HfWfn2grMNHRVaKqpdkAFCrbIeJShONFpl7feVu6AyRW8Cnvb
2Sv2/rKhr9uJwTfZPR9H8WCkYtubXC5ZDftfFz5QhZzqIeGzyMQvKf+F1QQC+3HsuC5nUvUMgtDb
ULwcM07hEIZl4psRd3RXETN+FVCRdzLdhHe6snUG7AkoyLMq9WqQpEID2dmSoMrQz9HEEXCmuAPD
tunio3yWGar5cjEO5eLQB5lZWavFvxSArtRWltjsHGljA1ZCoL2YQMvAwBH001KZss2Tn/fKQdry
jlXiGSGZ1hOT0u6aKZGgQJgrxG0ktpd75K5k0G6seQ9opMwEZ2ZnEJIiDaSUEUoDzJVXTV3tlwrb
lEmtG2+cFysvEgBJPz6BMdgDvB0nVn5q7uZvmbZv6TWGxO8Gad0yJtXGZU0zs7Zb9zBISNbNNDJ2
J2Fe6GZtdMy7Tuw6iLKosBajRdlRJmBW6iKx38VDbxTydnwm6i/Vdlz74NFEGJM9uOYDd4zoyA2j
jeQdksr/sBZVqNzX/1/zWgJ97U5IVmqu/wjtHgenoajsW9oZOrDZFd6JPEiV80HP2ZjdShZgwkUH
vsAqsNFbamZ89IDdlyrZLR77CKfpug+es9w7DKcWy/OP26HUI1TXQ7n+gn3d1VK3NrA8ide80XUh
TLKTLPI3TkuiDpvO4DeWa2YbaWmKnNof0IOWmW5I5ls2LxpPUbfqaV4jSPagr2/hOHShINoNCZmY
jgjwcBMV8lnw1NcuKu4H0yiMPDjVl8pish01Orab3UZHc0cUAXGbqSGjfGzUcKPcbSrU9kOm+5Np
qy2/rrD4lnqQ+LLzDTF1MWkDSlk9CcPgYbOK4cwGnt0Sl8avLO2LFH98o7GrQkr2nvdepWmHYR1L
52zp++hFokNvacdMwqvZzmkw2CBxf4HtXW+1yMiGl7cByycyCuwq5E2qsAgGFhiGfPXjBm4wYc9m
bqX01TvqKRkqCfcvbYctI0tU8gscXx6DXc7LCA7obADRTCVWmIps0mvynC1U8yde+6eoKpNboGjZ
8nVe/6LNS5zwKaPm6+j2M89JDjhxjl1ndMWggJpnp1797QTolK9mzmd1G1uGLpw0ODTdP2YEaVPJ
x0K9ZbpTur5yeMnJc6dp2l/VNAIiESrth8GvWXWzFL47cUOf5ZGUF+ErOrmUXEYaegcLrzMH50S4
2xjwNmuGQstgT5dg6XMrwWS2y+owCf8LgD8cWRhqbaGqpKLD4TVOr9qNtp+kivdocWwLnKu1AKFK
dIJImlp5BiJk2xrr6xcYMFuMGyKDFQ/h5QOy6y3Kg+H9lzcJLrK6K9fyMq1VyDUNdfDtssrrnHl8
SF9O5UupBy7PdehgyqaFMNv3H4LJWpydNLUTuT5ODswSzzo49ihOopxRTGoWE4dNnwhxVvcU5PLA
WG9ppj+/xp0Uu/T5R4lDNARXuNNG837f6MSWU5c6+kQq9ENa6XpG9HxrGw7PAVg5QqfJe6KK3iCk
PbRVTWcftMk2IwND6b1+1jViMAZSizhSBu7UehE+IHZB8Wy6aMwY7kRCw6knKTkKP1RHISRtqyva
6fmLvzicJsCBjKaPsSeNFNsxqEb2ZiGUWp170pv8Pc/DfLux2gwa4UAIe0rMxCSXEzRs4/n/sV1a
syrO9OYnYOALbKkW446H3yR1r07aQggam/v0rp/7IGk7QNoFpp9+UWBtQhPb+2TW6PWUHBirHOqJ
PrnGiiAbwVo/aklGPT/uY1yUL97IfKP35L/lE+u/FM3/DC0slvgrNXHsRA+X1pvgoftqx7YnkeWf
bjzDcL4/Agu9tuu01CVUcTlZFXesMepAt49+xXPB6ApEn+UACCUBIqCj02006ebdN+DTMIo0RHb/
2c6pIyLgjdgCEHO0dv2Ct6VvufvRKkwK6L7Qelchlpwnw04vmF/22GHxGwF8rJtH++UvsWFz+wie
qjf4Gt192aXwlUVnwl9zFzlbT2GqkCD7/AajNXvWjRjXjpmsoxruxi87YnREE2sX6SkJY33Ifwwf
3nPpXuY/zGZL9dcNq32UOb8kdvUJ1RT1w302LBKN0Jgsi9b6xh//yv/m2S+QN9mMrS/j0IIMGHVY
2FvvNls1YfKF5SiV+X62FFMRxxmpqTS524Cn6lheJ442Y3gCyMxhQ5GltmacvEFIvRimKyPJyQRt
nm/CsadyqZLHm4WdTFXS5sz9tpVIO6i6p4SV2BuDUCC48731Ag9PrTldxkLWY2CWWMy4rLZXODRw
6ehjD6w+4m+jsAqS71FiGCAPdLqEAQ3RiNakd90W02pHi9GzzWpVSawyDZLqaQgNsRV1h/rBNldm
3kc5tDnxZ3i4nR8Pu3HwC3qIM06f2H8M0mHwF+WJJ3zxif3D77QTj0LeNi8TNxoZTRzm4BdUKPKs
NfKTpkTjRXpSdDIeUzww9ST7Png9N/nPX1sbURT44a6nU/9v0SPD3Qfiga+kKcZ7TlferU4VGpln
Xrh9+KPy9iFF4QWNN3734blt6E6As/x1tR/akAIchp5P3pfkucGhxV89g84onQgfyFSP/TUtVwnP
qiTV4zDwvmSYlJalmSbr/6TTiY2vCLRc05MMnLDJDKdhMPkkipqwA9MnTm1xDVNgxSzmJE/KqZse
octA9iXyV9PrzVWeLNSIHTJa/C0Gx9O2FNUwf7TLrrp94Jaxg5Qi62h5NJvYyM6uBuGB+WdmNy+o
LSZ5zajcPRAVWuXVzuPVomQYSoUB65d7S6senl/aekjTpUfJ/GZmHRp5342CZajgKcAnGKX1+xwX
PhQ1q3DCklsN4SyWnVCwFBrHJeO/T4wbdkP2V5Qyt7a+scE77+rNl8kPQ1q9k+/lHVUGGl1+PRbU
kJvx9lMz40RH/8djUr75UXP8dtUdBrh5Km8td78HCucmZ1LH34M/g24glmsz9bnM9QeWg1/0zcRP
qPPZSbJ9jE7uA5I3ExR+nc4SGQcoo9ThA/5jcl7SH6w55iuLoZiMHAM1WKdwyVumyglbtp7Z7X2a
IYzR+YYIH7TUbvJJKk/dVebWJPMCnmgQHz8VpZafE5NfqjEOgROKKG0DIyEIz40ZKisa8Zrq/uWf
ln0CAsTsZjoz5tSEZe1M+MxKgMf7XCkRDkIYZ7HgjxUOquXRV2FX+mytni0rhXdjNyQY4o4//Pod
lR6MoALPrB6cmAxWxFVYBGT60FEJqTAS3LJfD5BPfsy2OxYk5jlmHxQCyO9pJgUJLDZtkfOsS9fx
gOpo7zdF17ox+e4gXRaCLA9cxvD7jGyAxfE6bQhAASK1lVvt3iNA2H0Hoz0X1zBCygY+lDtKykuG
Wns+GFii1E4AGI8M6nhbKJWSj57UmJN5Xm1KHkJ/3DnPCMdZL/dwzMhwqU6lB4WV67DfSinwNRA4
t6Q9CGHDckUV8hbaA9R/IFTOpCEQ7LSiEh6b8c5ksQmO1ynXCKMC4JHcatULmMz2utIkJkcY68SS
Ih2HoK5uQDA96bFE+lzqrfp8aerEotBshIn/uED1dcr2EMJOt/PbWBTxZttByGMHJ2gtyZbe0p1i
oyFR5HWLsv4UT4jfIVx6T/FBOKW7KueHJ2WPo6AWe8y3c+/ZjhxNQe6gV+2cOqoX91Kk1M5LHT6L
0fDFp8bxzIJjfpdgPuy+VvFZN5ek0pSgxI+uQx4q3sFcQJhyuvCXOiFqTew33YYWwVNus1ffn6SB
Ta8JtdEIgDaEsncxWuGAgo8Gnq2Fy6jmtvhiPnStY0NHS93isIkmhH8OlxiyKG+gAmQXcIdGadYS
IqGV0momDB38vXGPdhMlneZpvYhlILRJndlNHb5F/nl94rxyJpqd8yoXE77J+NZ9YA3VmbBUWgxO
XNOnaYR833CZh8TJPdOhE25zoqSVNt86YB3d6ATALp2wM/awixXCu8e0p43UJ0KMPkzZPzJyb3Un
AoTZi23RsNKdfkKcZOhj3+0DPlkAip04GPLBUmvUwkgJb6Y9OkQGneuMcTOje3YMTJtHLoDvZQQ1
flzuuor7N/0XdFAHivIxrs6APLz+gQJN9GonNIvI4mL/Ts4TNGgD/M7L3ksNix6vXNtDSBQW/dme
sPSqnGuCewepDyOwm9WORuDrbByDjdzd9ayz1JHjWT1NteDBWfywNTkJZ8iU2jbQ0e1mNcw8qsjk
oAl22a/zQi1toZgah5AVecIN4pSKDFqjiI9GzXCdz6WWUNyuu2W2Oa/hQLKtO7NaHBhANRmm/OL/
2QZlv2ZdNf9e6bIiXZPiet0K5KRj2cw9dviXzOgJ8AAM8z11KDrIQ6KVzT/m0mo/yYeGh4/i18mT
V7cJ3/wzdEZ05AjtNFDrIaNSIfbYg4q6uJjPCtJomBwVQ+WpD2OSZRHvU1QY4jvibnPwYopk4b7P
+sjqY8YGM0qZCLC+9LUTPmRWD2gMmgHntiyLvGnEctcn4tLj+igHHMPc+A5jwbwETAxPkXe1fX5m
jvCN1cVnox5It+ND9gwcVso7RfW/Ku0BwxKpEAWCDHy02ZE2J2c7ipprRfYisljD8hntMirAFm+F
r7nfIetdp9ejaUBzQqXAIeR5MLSmDJGK3QH+jPh/lxMjSxTuRPilfGYpOjTD2NVkU/sM9J4VAw/X
ZC/yKX19jBJgKPLcUiCFB4kpMuRTvapKGvia0d9ds4fGHRsDqHc1fuxchfDaPgy66iPptzCwyECs
uOWXjafcvMIf1n11Cg6ydLrh1XisvSKm1i80hhxWHg0D5HPQAYE4+oNlXUbPF82rO4GZZj3cDDKb
7fFwz0VWrjDLnkO/VaDEfIa4efU3zS6U4pveXS3m541WbLn7viS7Mbm6cO1A5cuxH6eJSIsMALfR
xqZNV5eDBMxoqSvOo92YRDxZ5IeVXi92xTHvit5on2qImu3URWpcxttm5jRacvBdaxMIO8RW99XC
zAwlds7V2tvNzlrarDqUQVTI0lBlhqYk0CL8Nl00CfABQSRavirR6Hoy5PhUWJ88BJ2XuUKbXIRs
oicAIaEaE+8RJ7Q3F2UHpZpb2i2f77bdzuoEE+MhrL1B71j55jNl0AoVoQpLdugWsahC007vdkxk
vCD3jz5i+MHXgQ7+q5nop2DCgJOq1MliI12xjm4tXTlI1OeXZo5o/4FTGnvoq6JbE1DkNHghFMrr
vc2gJqP9ji5DqIqhmikjSqlW/2H5y2/tiNCdfx4hlxX8T+WL2PgrvUhHsjkN4MIrKx140YyMKY14
qUiJWU04OCrnTTYa5XP5pITjTR5ilXVLuaXbj6xdR882+1Srp0hYlN1x6p3G6LnmBbkk208u4geS
3kb8ANig1mw0uBVvVRiA7OOVVonOc4pdNbjCKJ67MxnhsQSygkmDk4bhFa5on/M1ktggjc4lnJGj
qMpQB/Gy/EXf4gjFaB1Vtcn/8sgq3MxiM7RGWLRhbesHT63kzfGXsJUa/iDKeINO/JvwPks8/GMw
zWFvJLHn8QdQmyjGmM1YRPfkRoN6LgPepN2CpdWmoHfsUI1OYc+yC10jr9g8fS9YBzvT4PGN+0c+
7cA3UctqLK9BA9vdqqCUZU41rmpUgOac05cstF6+rvTQbj/cA3ebD/1oZK2etIR9U6NK3hmHdrPc
STnSOX+ACrlQ+k0gMLqzGcnh9bpvI+unlH2YWCsLDbJ7P+x2rlYE2a8jnMWhAtYYOV9zvaN1tR6a
aaQHYe2Iap6raYr8RW3/N4gRtUsM38TAcyJiEc5p2f+bztyFdzdvwYwfCYwKpKf7DJp0kqKWeYXV
C2W4azlwdzRzRX3mEBvEF0ATZF63E2FFadSTgAFcwLz7sWpeD5yGFdazsuEoITsAsJ2uYRwL3zaS
34C+K9DeElx3GAnZ3Cpayvr62B7FxynF5EI/cCsXQNhLqX8C/Lb1MyOUW/MxVrR/3CmuxeRAhD5K
yNr12PtWEIwadFZ5BhUWg8BDnY27HCrg8M6rJ4bg091urjwhfZ0/UBS4M4z2LR3+J4cP7Pax5hLl
yNGXJGEm6D3+HaxkT9RXdkXIDfW04l+E/Ggks/B5A2+bF/y5u6ctnexDsU4aXR7y5nSdz0ViUp5d
LSrntXbayGyG07+I/zaz2N74oi1mSDbmL/pPY3PDSyUxbXQvgiTmqokXuCmzYFw1sFVmPSq/V0MG
8ZL+SY8bMIfUVVQTcSpIPgytsQ1660f+gJHZqVuCC3CHFmu5/9FGcGG+rF/zW2nAHPjodMJuiFvQ
g/lKoxpLT6q2taVuyNtIOm6fDdCE+Qytsg/LxoAkD0APeBKywB1a6cJAVISDfiYkwUPcnPHn6gY4
HjC+5HlCT/2E6oV129C4d1P5oN5RsVtH2FZ6NsXVgaZSF6kpjbixecAyZvcTS+WeRLPbsENZUl84
hbAkhkg2ZE1YglgrYlyzv/acflR24FAH024Ei08lms5nbdKos/CZeTmJMj475VCqrg0tnvljOPDz
0AqDOuwX6vbovnoOZauq/nxCLIWqddljSgU5ed/48HrfQJtWHuJ6nHM8ZAk0XcjjfNxsI2gfE3W6
tUggHDN2wdT+OPxMWrQ7iYtHWMyrH/w5FV+oE+WzhXJjXqRz4reajLY2gvYgU+q2aM910+ztF3Ho
0CTyZngCz+uhU830GSftPJ8ZNR28Y1tgvca50gujM9dHOhfcluYgKo7CCIeI9eTvq9mP6PrEOhvu
47cytqwsUZy5oBm4DxbxIX4neq2BwseTK8W1U64rMVcmP36DCOo7IYWkpl9so1S5PSOmU3rRMuM/
2sdZQfqYV/nISRYhhB/n4g8mjn7V7ZlG9sn5wF9oLhKwzUuTsrhalYrqHATECaamyGmxLELbMRq0
2hQksr+n1C3gCDcM6Z6SdVJbqxQnT2gU6fDtUWYCoSvsBTvHOdSEXBSLbRsNmNU2EApoCoa5n+Tz
NwpyMByXYPPjtru/uil2xcLte1ckPhSeulSpZJJVbNH9ZYgMMCCQU2saUoK9vSCaG7iv2RKa5bzr
AKs3Zc8wsFw3CNGwowhxyq28v/JTfRaeeYYj/kZrOR7z0UIArxva9oW6B6WR2td5HyQA0tHQGyTX
G2c+iHSISg9xZ5Js2tswOgWXJ6S/MngmxMYbysHVKglIZ+b6ldIZgmT+eGJXEJb2FKvJ/EqGLD7F
ShPstvrhiMH647iO8Rs5Zyhblf9kh82DRyNgJIbGLegEF1KwAcHdD6CaTJvspgc2TAuqAZOJiIKk
EENCy1VG//EVgu9iIdC6wBhFRSVFyKKcniHdoRgSAwX1+Wu0T4J0miw55NWpPlCPe24cLgPALyUp
L+ibca6e2cw6RBb/ajy6U8gPZx8R9V/y/2GWx/M1r3qxzRa6YMvIU0xuLydTPWJ57LC2J7+4vaU9
8MW5hjFrpEIEC9Zs8BMAfssmzdyiS6LnN3lGNqDxqoUUHOP8cY1Ou/Pq3DQOdT6LmH09gchMnxD8
PrCBNylLZ2iUB5+EdD8iKW36cuKTDSA3c5fy0bCG0FEim0MrLSKq/dsGXX8xhD55cF5VAfGV+9hJ
8q5elffnOQ7/YNLe0Nat8sFDv8HuxZBUBg6mRV/gcFC1DmGb1dADAwntXx/cklq+nyogDho94H/X
4R2KFePYRQfDDwOwUvGPCUvSBDAjYAmjqciKqslT1ejlcAH9us/pPGutisbbf7JPvKMJkhOU6NFM
pmgXzr90CRmW9v+OKfkJ+GmhiYUFfJj5uGi2A25qDVSzRcTL+Yd+TyWsLlWjQcQaeHT9BDaGZOKa
1ioyYMPX3GEKz6Zsyukvy/CffkbRm0LzWxb5GZYTt5dwDFVVNngFOLbO+QYxe6tztlxFsmuu1CJK
uJoj+W8ZLs7juiA4AWq93/7aJAO17CBXcd7xHIXGJ2NBrdmYbnwsifltIFNWjfbIG45fIlPMVys/
PiIQ3XbW9cC9CKnq4ZUHfXizAEb+eNSXzXM7v/wdLa0qATXXF6l1xatqbNsFkBzQ/3MMgWLQX2lS
yNDImfUTtcjtQ/q7zv+EfICf82yBeqfdyt6pCN2sJ7gymmANzMeIhTBhgcvJv7wPba1BAQR3fumq
jJVDiWw5Ouf3tyeDDBcy3avQKqxalLAhJxjr6Jzl9H75h4ds3P2ucDEp23iiFPcv5Zue05GfZIoZ
NBYdYrV/4NgRbWxHlUwGMG7/y/ivbCU9IjuGOJVh00atLT4qyDaAx6UEuR2V2Ec7fxWxm80uNkgN
28kbo4A0VxLDRVFrVT7EBBDxtcwFteGOit4XKqn6chF1ys5J/bZ2pJVyrgsnqMX3H3QPQc6ZXrbZ
/EkbYzu4svCqmobdullZxJxkCsmlFaHYPIgQ47A8klhSJnLQOM6fBceAGtRUmVyMeGFvo9XOwpgV
0fo5alh6ZLuzMYxxxeCKdAY7YLZQNLGsrYXE7PM/zFMNiH5OFv4agvEwUZvBcstB+c7W06AECIhH
VGCb0unAVZaKNB5TJvAcxEHPYht9j4Iyfvm/MjZkIPgqSHY5dCMs9i5BbxKaoA1cCttG3YR6cNMZ
sC7jhOluuQVZmW8xfhVTK8rhYEI+GE/I7FLEaHSDoGccaVlre0Jubs2gDDbq95+ApeFB8g86IHxN
9cMhCs90T4qcElSQAE4GTwXUG9ddY9Nuki3/rftc5FOm0KaqluoDgRerqB8uUUhvmdKIKJ4jKBk9
rN0uKF/+JVYsCOqFrFEwtxfWvb8WXdALqpkMfHnHuVu5KYznuLfU06IeoHtHQ/iVKf0N3F09QWy4
KDg0O+/8HtcNMQOzGEFMZL59qtDzUu87KWfgdFPWqsfQIF33MLtn8A8QGGxIvltkP10LhonN4ODT
V9C4TWl0GCfePsOSM6cGpy05ZzicuFc8aU9uv5zi1CQg7JW2yEi9mFbNGNCs+G0SaqxA2Y59Sty6
u+MKPeCQy4kIAnk+1TQR25T1BX7iN20A065Zq3HZWKZKlLfPN9ZSkWMOeokW66yw2qWGlDo0TpzK
7gyX/asWI000AOT10TUYTo7k1Ms8NHnRgdmCm2xeVc519Zro/r/yIAIyo/1rp5tbDpqb+Onh05L+
qdZXKhUYfJVbNh5IWYw2uVTjRtIq+AtFzr8VTmQdQxDzjPYyAzmawmss3Xovld2D33UL483NQ9h9
/MF0Cg3mKhvwE+ST+oPduTztvCPUETVnOt0pbV9IXknXHNbs3NnNyGUKOXETw1kxvBznwaA0keyX
0jkCMYOKARyLKw2sm/ZqCORkwBYln6tz8yzxEiI5NCQ9fg6noOt18GTh1IlndFDaiHvQPWQq/2+z
MthAUMFMWz2w6wULGorTk38RlWuP6RtZGpJRR2QvIqp6M0i4dLBT14FJSGB8aoRS35nzlHuN7j5F
jiPHEQbFvpDAhtsyourkzuPOuo5FHykQdBfVNfVmDM+8aRSECKHCOGZ6Y6ZdYl+ETYrbQwq9Ujc6
O0J3fjbvZTNmjiCq0g1mGLwUt3tk6l24MrDZ7gxDNZuYLrGPVjbHid7jyIObnh+Q7ZIVQAB+ds2i
4B04BzPzoxKJrMAwYc3VwmVwLDbpzE+P4zdJ12evfq/tC4+X5aY3nQx2DB9hkho0IpUP6kx2ACW3
P4JNkP9A2frbGaYM9mD1pU/xTEoHonPUf25fwhY6lq1iDHxjyUk6R3WZIszK5CKf27INQba0Rl7t
cNUg0JWnt1rNrYrcgSicg5jqvJNAWW+0t+eYczU1fI1ssuNQ/LMzak5Ik0uHYALzSMjkw6ltDSOt
I2YZXIC8AtTi5W/Fncx3mvTb2ZVpcGUQducCBAzOZ/JCiy9KjvWHyeCDDQ6TQOFONWSWntbyHGDb
ZSoPEm0L2wM7OTt3XviR5F5thv1JL9cBetLP0G2YAPs/zp7zXGyMLkx3GO2NZSlfKGV79cESv0Uy
T/sFYyJqF8fFHNxof5aQs32g/IIdz7hhtSTomJj0ZASecDDJFt8AnAQ7OpgY3S//Cj6WHpOXBEXx
yFxQuOwFOOHagUjfVmN42HYx6zjL5si/fwTzJx8bJmdnfpwFSdXTAvxoo4vcVyBXj2MNzzqKZ2tK
X+5G3bcluchWi8gyfDhNBw8UdQ0rCdmdDipcaMJ0av9FQCFFZj/zU78L+piDZ36RwSbkjTrqmvW6
gRnlPdC6R0N/0ZQwTVydDsbekxF/2Cj5+9NAdX+IkFt4o0ZYiN2HKEtO/A6tA8N9XzPAg5jNCDln
S04N8cE1VGJpThf86ajZ9wRVzBl6wNBVaupDoaS8K/tbMgGhdWmQmqJmt13TPcPFHZLfchwO/ZEZ
4Ba8UMzBY+X+UoJA/OP0uHeS26IaM2XtUUj735RnT/sKuoIQS/WZIyRDeybdFISl+7sDC6kAAhFG
5/iMeCMscKQRuD+7aHbK/NwKX/obAp3rfja4BH8rqoh8/suIJ7zofhH+B7PfL2UCdSq9Hjsh25MD
+FgAJbi+QDlKmSaaf/xV/hasecx/GOjjZveMVEAeTQECLrnnPqRrkYNkmQRyNAyq/23zL72n7RRJ
GcYd7yodixmgQF502DWQns8Tyr75A7J1C83DKtji6kOVmBdSn024fDpCrklpRhL0FreSyL26VT+k
3GZr65AVmTsSXPntWVAMGEqrmbs6ziNo0kDCeP8ZgIRMU19AJ8cXsmC0k+2O6rUAVCZo5MfoaxDN
XeN6LJUiouRH4n8RFu/psFBPH7J9sD4g2A579qlMe9iytP6UgnJDKIhnOJ4jVkYTg/JkJe+Lkipk
RntBNMnlgm0za82l4+Hqz8H+h2G1OST60J8vY4ofMGi02xRCkYEZFmdrCl2XGcCSr1w6yZZg5SIp
vGWsia1oAetiFuqrLt03oh2/hnUeVgtJeVpeQ8dR2uJ8sdZ1FxbIZlIVbe/9JpV8anIBwTlW51fi
dfIoYLnshciOM7ydl+JGZsDqRy1SVnMNJ3Rz1GgvKI/l4pa/iaJXQ3i3zw0mLAdIdH5Vqodut3sU
46jD2J9N4jivS2FcAIDw+R4jkSkU1jiSkLVaZqNnMSQxZPIWoXjwrW8+o7BbdQij4IMOfRQ3dt0b
xxnyAaFGgEAb4gGMnKq/BiCd4xH6PXLVQjJq87K9smX9Mri7FjKEJRaHYT/J0Youu3p8/qXRr8M2
GmqevkYsegEwDw2J0U9xGnpxbh3A9HoRoX/YdvOOqrZjKqqp4VymhXXpHiVInrBEYWRsFCZbPAfS
NvSlf6V32XXLJLhGAhcSRrOEUhF8v7QZ+7dNUMmHBn9nKLFa7vWGvlQMVY+pgEgCCYNZxYAzjSdS
px2DAXZmAK0BkhlmFhE4Q6Yv+/Fg/HRTPZyRu5R79aUyQjkokwELbx5xgxmiZHJB+N/aHPJcKgHf
B/jFsXq4+dKwv3TbIUKBZsjGwf5xcbQRkSzutaBRbQkklygFA2bHTpp0x+aQ88vX5z+oGACn0ytk
uLF8y0iZnODnFlKE7FpwrgSHp3h/ZveJw2ztRDt3MsxPnaJtOaK+HB/l+ypEyVVea6aupQ2N8rBP
n3FH5hJmRkTzPY+9N9rYukcH8/hK1cUmanRWtyo2uesT8A9rLl3+5pXWpjx0Ttv9a9TuT0FrUrNF
nBgbyr+5n3027OUZvFVLjAfD2TSjBynmWUl0Q8qZiQ+e9X+D1aNETf8PWNJNxQ9yGH2A0/aGEzmq
LdNB2SQxn4eSJeiklrEJQoeJlUeRLbtV/uY/fqab+x0XmG0nA/0fkme1dzU2PVwSXaJXGjh59UxX
g7lUn9QukG+lVsVoYl62x2CqZ1WSgC/pkbrZbuJlupcsdPzCiLmzD1pAudcCUfcaZUewEPQ7D/8f
Ko7da1z+HuFjczIA65+/llKz9Mcb/1ea3iBo4GysQHjOmlV/vIA/z8drXONw3/ZKLnvh4W9k/Rrp
Z5JJQ9tOKwk99A0uI5bvCc8HqpFOZ1SNlg4evn2uODH14pOmQ6MwfmFASpvgybsfgj9s0zUh2jyp
vXN4GcjKinHy4BkTU/JsF3GoVdvh6krvpTWDbN4MIETeFIMEcv8uZUQrdu68cg2FJUBxglcLzLEA
uAr+Y5fJDD3F9FLm+3TchnJwa4r6R+mzYPdBO9NXTlrRLS2Dh8rAl1Qs1Ib5z8/3X4MGlXoneebM
Ou5kgQ7OtG7RjYUGr269YrsQaDTQQuu91Hm0kHO+Lml1ZsQV/VRrEWG10d75/+3S7xYy+yyLwtIw
MDN68ocevDv8ntxKLmG86PRPDZ5PN8/1KNW7WZBnwrFRdtMbF/N+oeboErUv20KuMrChy9hN782G
H+Vz8O8vJIDaO3ZayFnkvhT3pojNmHSVcjQvkHhi4ofLEZtA0Gh5uoHnr3aZIiOAHuBZKJFxUTgF
zqxklb+JK5WLz9JIQZ4YPJHJkChLjPFlyTiyrKXYmN3rhwNh1v/qoz9r+VwIYUG7GMbl47PxHq07
YBbYkRCnwXbp05IaAqJNn0DFnHfMysTUPdfwUbjnslN6wihe7M4CvP4JtX7+tTHbhiUJIgHcQD0m
+K/L88zt8L5GPLj9EhUiNA3BvRtfzRaAUfgNZDzKeTHwa8yM82Yt32QImWg0ki0g4wtym7ITxT8m
f2Vd7rElK1ypHBH3jiHzU9vueocgPnYzvMQCyXDXQPs6n32Yp6uP/pMwRXkpM8ZYCBQljqfUn9VB
LLpHS+NjgDNN/Qda+F4qQTQl34Z3YTAPsJdefwpkq3YTOigGVvvTx+dcyTZGxdg4Tq7nbP2suU2O
vtop2+QmRRiCTJf9PQ8xXAORHZapd8YVbyINmBhq3ld8W+/tH8ZuVuaEaSwIhcruFcicKvFyd0T7
ZOm8VFTmpHuTzp8jL435X45bOfwHSrN38bdhlI2sRep4bAjiFRZxuLoUCD/4wdndoPxprl3soGAH
jQXLKWDqwKVICk+a9nX9pQ4Jv7CLrh+KuZu0LcIJJvBzqCh/Go5oYT5LGxz3v1eEWxTeo9pUB4nH
D7k6+LPhe5rQyu9PPFefs6V+jCPXLrboWwbHG4zVz8IDdF0MVKQS/tCVznT/wSiwjWJMPmeYLn4R
S69EcncFKJ9lTvuWXAlO58B0ABYphQA31q84+yV1gpoYj1mjd9v90BgXBEmYsvpDo3QQHrox4QGW
+cJAamPQzjk2OcdUeSSu40BzYywY2/IYZjhRWOF17ijHCfJdBRBp2Kkpp5+r6gK5ccfTiNiK9rTE
/coLDw/4foLWORfcoEdMrOeZf4ra1yakHVpEInlwW3ZCS7vcwPmYPvY8DfPqUlqXCDlBvfNkYJvd
WgWwosR/GI7pOjtwjgNtuRx6Iz/rNwERK8L7SR4AX14Ua2AQHeIhTb31WVWflayVOcGrSmuSjQGL
689nHLQ+usjLY/iVcKUCYwiGzb2Qt80v0rJ6N2opxN50osKdWhmN+758gY2cTiqOcgx4Yi3G3NxK
ezrcXsDcnSVse8hEncBCKMIzn7z4zlT7/55OE3hOIdXo/bfN3Pf4Bfv7H4yVuY7olS4CSqRyyNup
uaaiwMpeIfhWfvHIojYibpCSfPpPg/MidJpe/c/5wQbdTkD8QptfKTaM8Mz2oRPVq3qg13RZhGST
TbYpcOR7Z4IvVpgazWA8GhYuIXNfLd7tXLu2/spBS3LzZ2i2HCX7cm+rsRxH4fMfI1tMeNO617JA
37iD9ZHYLhnUg0F+QIF2f7qkCykRD+8NBoHZLLjNJu+R2r53CP8fh23CY+FX1QCElkaCDddSs/u+
/O7OCIuVocRN8SlAdeqF/AsveLc38cRRthmXI2ulbxXUo8e3gkKcWV8VVbrdB/uYU1di34Dfgx8C
sgBUoXHT/Qn0iiK38MaDZTgi0T1T0BzodZUuumGi1HvDCDecxNfwaDDFyoWTFdl6HOZf2Qvq7feN
lUmFqXCY+AvWuN3aw9yXLgdYl8p1/935jn6SAN23eg2yciN5pbzc3DiiBCDUBaPqh2pA3cfHU/ca
hdkzTTNjqWMCOHPW13maK4HDSE/Maj8z17Qr6snkbyP+v91ZxOvk/KLMyFebJmv5DyR44p2yE9Tb
u5M7Tsv7R3gtH2wlix3cWr4xAfH8dTlheE4qrL7XCA3i70PWith9qCwu1JgoLaqzxXG81Ce3CbcM
KcPsykY+5WjAjqIMkKSD8R3A1bpt2Ly+ozD8wybnFvJv1cIfPvXpt71Ci1IlLR9VL1L2vdHz6O+7
wL3vOYMhWXQiwMW97xG9oAQiQuegKRaV36F8s3Qzj85YXgaEoTTdJrW1OLojnIbpgDLhLrQukUe5
trDdKni7Tsz8a8tbMRBlMMO4SUSQtgIATKysKJaEdSkP4ivL+I/5+PNV55PsIP8+IxqFMwIFwtWU
cRH0St9JXxEb3ZGUAmxiBUkX18//+kRmfTX5ULF906OBHpLtnNM1jpd412jhUtbh507VHLdC8uOQ
m/57UGnwRaAFOz/OTIhaEv4GAWoEPozDbI3wPnpuqjVeQn1bxX5UAuuCXqZaC/NW/50+F2ZrieRT
QbISQ3BB6KU9uFKxTwTVQbP3Bp4GAMsgS0QCRmwqvBQKm3PAmMlcHS+NhYYN+4dz4P543rOoDiPj
zpcSHpM0/FnOVC7NWHIOCB2UQEA/674biMbtDYGSVS5ZdO1Mb74KwvkqLEtWr8zQPB68t/gSQJiu
sHXF8cyYZRQvREH4VWJtXLogIUvoRV0E5wwOxf2NgfZrH9a/AfUiUs2tzWejUtC92jR8r89nT9Hh
CPONCJp7rvgpdaD21Y5DcuQcJHDCzFnlUm0OtA9QpTyt5vY+efEP0OHxkhXtNzU39tNiIDSgp5UO
kDc2nJXd60rj7EwDBCtMnQW/84IDlx0jRn6ImaiPQaaXF1htB3AQTAe2o4e56DvYo7MkGSwqoWz2
x/NKesHz3FdFTHsOQEGpCvpOKvPVPrn73k4kixp3CUPfuN9K9KSHpGyUDhgAWDU0vC+WY4wkVKIt
LqqXAmQSRFxjFUPVrOO8iKHS1CpImgUnF3OEPAgzPivxKYbgaMRKmjKGGLBInlzjA7aCrqJV7KEW
ZSUr8au3IXq0XZV5wxsYtIYqrAJRijL0lGS3NQMLKeqD0Ozx5tZLZbALe5ABxyb67iT5TrljhxtN
hQCTjpbpOEgJfsItc3Gj+yHb+XzqX1HU1KObA6cxroFwWGGEEy+wxP7PBzqdkTeCJqEHiu7DfpDf
L5DWjdTdKea/IBqgOC3laOm2inO5Bd7XCctZrAmyZNITUOdWpU5okv3RuZAcKah9GDGk4vd8v72/
I2lQ8k4gkjHprmrzTRS3fcaLVnZXCNYnXGBXOI/AgcPTAn2Q2KpzPlwVFkx07oXX3xDkCi1G/qb9
qNXA8AzVS5Jm+aBCHKzHzjM32MijJC3tBnrsAg/EIsb8g/g5luvvtAeX3esXD96HR9tdQq0YxC24
z8xNzv2oWODOVymL75mdHiFEParL48lDqV03c6jgdnQzRmJ/+sVpwYKHSUp+F7XajUqdxvsp7J5k
Y6ZjucsjBdyq4RrokDsgB08ooXLWWca5eauqhktomroe28YY3mLHPBDNNrCuFnOZBAc/coU+45/X
gQFDEF5NP6+u7F+bgjTbsF9jme0QobacByIe2bcFYnLIh8IWRjkW0hCTuJKudS2QEl0FQ3Kh79C2
ZNrYMSyHR5zNiIcUC+OiB5PsNy3nc9hTSXklNq3G7MZnJ+VnSKuKHgqSl1h8Pe9e91aIYtGm8Jym
JBao949eTjc6zAbDKgpvvo+kR6a2rB7u6SJ+ojVX8Cg4sbm49bd1leL13v0jgNjgYiRFrK3ORpI/
UdLvzyaOGycJEtuvFsWXAGmBhUDLbVXvkeui+j0s3zSEw8URnG2qsjtL4vFtZJQOQCwp4c9todjU
kRnAYzJPYgk3AV/CeBqzcTQh/sxFtukaK/IGNgkbudvh9byWN1wCy6GrXWB/y8O83UU2Vio9URy9
x7gbJB/QpCm7EasAqQ07GvR4EAkRXWcvrGaCKm4EbzeJe01A3kVSW4wuRb7e47szqd3PTaiRzqpZ
vMCd6T0ZOqoeWhr1LtPGLjO4YhhBxwYCPOCqVH3q47iYWOVEyLmE6Agybojib0U+ev0C5MiEsS+O
WJeDtCjyHstpMHUtM+vtm7veLCcea0GE0bDqZO1DLpsMpmVKfF9q2T3hNWDVecqlV0+IhQctOJMs
Vfh9QV8nPY5B0ESBSGhKj/dbn6HBQC2rJLdrwRfBB3S3ecR+bB4v9c/2BygFheKxkdtqkSMTWFnO
pMTCUKTzS7MdXnjHH7Cm66y+cNl/nsTYYQY4CH0LmUEcyQYJXJeK8Cxr3naG1E0fek28TGM/oNTp
yihPwgbAJja2/uF6iH0jfDJmbmh8qxuEnaR3VXAN4oK8t8hJNjpqhZ+3m3MqYdlY/+3qa6Geakbu
8AcBkP2aWUh1xiUoEVEgcyaMjuv/5hLAgmFVV2W+hqjKVomL5so5n3W7IMmKvBYhd/2xGZ7QMfB2
6vJdFhXEpeZUymazL9YyTHoQzWu7CJRwy51nj+Y25UitOJZWtQN3bwfrOiZIF0/joKNObXBGieMI
GzPLapvLUm/AW/l0C/njuEnXYK1dBWLwvmJfUgdYKFtupt4wtOwJu7KeAVZRExp3WymykrmDtHWN
ysREY/GRvKNdEgqGAnyfZBsirQrcxVD8xy/C5rh5Uk1JPhlMk5Kyli/k1pAJACoX4qG4cJJ/y87k
LszCKlwQ05679GZtAuSUunYCJKhX41SztCRE97007gww/jvSfgWVUsfIrgVMawl7mCMAunJJkdYN
P+0s42Kd0pQaPK43SfrImIaPP54U6gY880nvHkSt/Uq9LqyCmAQUlGa8NeGz51cbjBKatTiCZOUc
cMZ2RaySTlPfJS2vyI2UU3rbhHSc8S7u51zlwzkHnm5cheBnC+aXD8OEeciEDjKhSN+3fIfm/Hu1
lzfQN6ETyd7hPlIm6bTo56DRZ3SQpvMInpmOeT1l95T7plhC03V+cIKLqvbJAKEmuPFsrRAx9qw1
IUT7qE9F0qEv5qyw/zxeCCkv8NaFCgd7xUlqxhPVixT8yYkKrEcTvjWs+z4AOjX5KldwlgC9Utf0
/1JZ/oTm0H1ndjV6Nl0AWP7Z3r6ojCI5odp+om4VGDT+GiDOCB/E7UD71PFfOJcN5TePjy5xXk2W
wsjsuBeZ4d1GS7OQQ0PXu6JYYnrnnphOj7GfKsAPQ69FUv42UZ2WF4CxCXQrOOhr+cfpnjE3uKh9
IGF5z0oK7SBMlpEzvBbOMo80PkT2oL9H9g0WYCYU2tSplKQWUyE2J5sFE2tMBgGVm9mZ3nIu7OF7
E33Df3aagDULwxfUrNHPjaNliPqgAlftQceJJMlWCnhacwGRwpjjKscPyHBxYLQ1tJYmLZ3lHLev
Ir5QGgwjdpm5KzbqBvxQ9DdTAAEz8CG6jWOlm4kOzK88klJXXd5Vmd1sBCbAVEFll2aJUD8ZRiRj
ShyCI97QVV2Svdc5Q7+mpLhXPgP97HD92kioZd8wPoZ4sqg7P0GoZMT7HP25A2iRCJM2GHaUzJlH
REtSDtdCOoPIW/K2RQH87l7SKSFGED22j/ngbWilNr1gX/MBhaCgWuqo2V9nYIX93U9bq0UTptg/
4XbiM5cSQyZDFjWQNdxXMeQLKIjA8kaY+fvSju1Ggm56FDVeH24LUxPL7kwm8Ufr+brwGSgmEOcU
yLuoFEgIieR1Z2xshB/GFTBmSvjjnJlt4TAWpCTkEX2cUt3A+khprAiurAk+qF9kSy3OC9VKaG22
P8wp9Gdojvs+NTgc1FHtllqJ76gHR/e2zCSIF3VEMHFaXXo8rnY7IhgHk2kfUcQp8QuZZV/8CIDg
f61MwiaFCwKpQCPL74LpYQunVRi45v9QNKXsAOv5RTWx8DVx9qGABStdAKc1dJl0m/PTMlu5fjXZ
IAcHt7r1mDLClxpL20ArEMeMjOXudEIaa4eMn2abmgxPtw0mb9WtiZ3AGTvGYdW62UMh9HT+aGjE
3kthlrEHmt+mrf2pJ5TEeCyb892rL2E02NSk2510WhT3okFTJTh945Ld8xqc5gfnr7orvVy+qyuz
FS5QEHx946NOZKdXaRAM3S5aCm9HdpaXFLmN7xtn+EKFbvpFK57bEf6ZW8bD+KezKB0DruXqnZjh
DxTZ1nksdGPUSjEJg/Lcbt2MHj85eVI6sWNWhyqiyNRsHtx4Heilra4ZNuHrikYKbQt/gF+rFdo1
N9grKi/+jMCk5PyhanX3sPdQW2N+JYXN9251sNfv5G6tsXJWFj2IspAzz/rGCV7U6YrMORCQGKlk
/EYlzUURRq3uiAP3ecool7VymujKaDEGg9aO5qGmxvbDorByk5s2hwFswxP+g2WjShCS/PBxMFrI
P2uP+75cXYigYLRv2KjtE8EqPwGNLckWMMu4+8tihOZCX7xM43ElbsfETMkwcL1+q5mPbh4p8noc
+A9dNvMWQsRaPdKtVmf5xX8XJL/+C30PTnmHX3fbIhSas+Kagt3wbF+l1QuZiQ7pTlbLfMP9tVhn
YwdJvYB0rp1quOb6f6CxPfoMPJIuiy6xogx4KrhEVGUtY5j7h29mMeTh3cwjo/0tGNyvtoj9sD3V
0NfPK1sxjFY3kxnPnakBxDIRjBpEfcr2HZFloiUOAM5lxqUUkswNyisFX7hT41P0QNYr1rW1DlR6
MFfV18q6voIp54+g72vTXEmIwpz2mSV8U7uzBAwPAdw3JOLFIuopI6PNnDip5l/GZ9uSitdWG29b
fAAHgRQRHjGO7xca0FpNMhHGSyA06v+ZGVgseTwLdnXhgTbfPMWTRtadObsvE6GmI6sFyfQvOzyG
tvB/q184LSUZft6P/KicptrixE4Z31puplTgXQGChho9ZAVxanFvPvAASe6gZvmxifkcBrHqBQVw
zOKXAMlTM8iBbh1tCLYlFleLTj16g8cp5PWQrNkiEvXgQKPO70hzxLnVX15bqiKtPMufRaOw7Je1
CBMVmdPy9CzV6YIyZo/d6G1T64fuHdAR3Ldxu/SOubdTlGsCLn3DNdqOIoNDqPXVK5U84bkIPv2f
BgErtHp24q7SEXBOHxG7jGExPzbL+KuaUeInYwn7GKJiG511FBoGogJXUIpMdcwqkzrzcW+QZhTY
/Oa9/b4hiyXfTQ+uZ9R3IxVTEmw3dKYOlO3N+rGS4OrnQomfO16F9s+hQkAXNFuFdroNgEGEZ/5C
u7BVFn/0/T9/h5VjDyORHmrZ/32tBRCqr3ZAV3Yu7WZjZtZLrnAxehwi56u94qiRq0J9zYu3XeqM
lD5dix+p+1W2Dv4mOyLnKnP4BlmrIM1kEpGfl2ZF7y9OTGUE+3Qm6pxEEr8WLQIWcM1LBcizPasR
E7WKJNiqTHx0V6aH0k6dTr9q0h1xBTtvoqNmvikFlFgsoqcRnk4F/yjW3lB6Cid5R3hpOkfRJ7XN
vGQUePqOf9j7K7d4JWiX99fnMmQRFBe4/bolR44MHCrz/8bV/C94QxDqWTN40KYWyfvVLvEot0hP
pu4iD+aZgQNn71qj5+sdqZZcnpw6589cFJhVp5WKIdUqfZBaOrhfbP7nvs8id9xTSKVce2mJCBbE
Ct+U/f1yGNSmlYSgKm9i2bml4kjIf1PrG52mjULLK/hW5L9EQQwPiASZnqvB1RoUWK9Xb+L1y8Xq
YMkosxk53NrX2pJ7Izfp+TkUJrpqJos7d6AM9mS0as87QQRniVqkguUrmUsLRFeuQhYnISkv+6bM
Ty3fJjCBVZTGTwjXwEfhXcxCcGu25L2+xmkoozNVXQOj/sn4ehCYSxt+2J/mqV+QRSCmTvwILr0C
Wg1qRZ6QkqFOt+WXx7g9X0/GbPvThpQ4DGubbHKXp4NJ/JTZxRRzwZR4N/9lSoc3FyRz2AQIj5F3
JN28hdqHzoR0+zK81irWO9K518wDfdj6ySTQ6bTbeIsN71ZWDzfioprToDd0alK7QOxPFSyTDSYR
eR5OyOyVSwBQ0OJrV3miPewzwb7eds0YRLyNoTBX3KX6uJkQsiuCwOsfzbN+mp+utk0tKxMr0TwM
bJmeKOcNuN4KnC3VRf/34Fzt3BFK2eNPS6pvUu73qzSpBWsUrhwGdYnQEq9vraeKv6syH4PBdlUD
xGa1wBPrkR1VPOaoYn2qmEfayHgJ4UXG3u3ZlvGThqqexhTYj8BIGFfMxmDzWq9FGugC/xkYEXdR
Pe6tjGVEADD48G/leyk7hn9/Srl+GVp28BuaXWH4VHbEZ54fgeI4ey9DEplNHg5kuIJGQJcezamg
aXmyw1M8IYTWjJIxeJVcHipLV0Z/DgslYW6oqPpMdxQ2NMmHyOUXSlyZwfzdFCAOqf/zTTEvg3fj
T1GI8qhUIj9fYt/cwN7oHWjg6ptUrk5FAB5Xq/pe21oVJ7mip2hMEUHRbPKuwvhAZ/ywdmTiwnn8
jwwZNCXqF5OeLQ95QjO8IiE9MIs2+UWd8uru6A2B2hfaStkNHx1pO8zNCbyVUO9aTRODC5xy08XA
+RhBPXTJ+sbrsL36m0pOEnWJq5UqWx+hncbZWw502XIwQnGIwAJyJxoiDF67ulqTiHQiVMAXFc9l
kWj5d4CvLH9OjAXgfDX4XvHpiDzrLYgDY8Z6o+lvMzqoUj5gobt9aRX9Y/3zPGANJvqCcU/aqHHv
nDCc0l+iGsUO3qi5TOYBirgZCVwsoAQ5w4HIw9F3ywG99EmvXJdACBFgpS16p/1xUpObehPrYOp2
Bbmz8WXKEFCmbFhXFc8UTN5wshjIAj6pz0+JxHNUUU7q/Y0IEGBNTdC0iRoGitcNly8JLj8udaE1
KAG3EXNwpym84OwIUobrINmANZM5hNK5xW1yDxo2qv28IXW1avouMQqmVCwp/S08JZ7hhNP3e1Bq
8X3uVVl6kcBZ3mUJXvJKIiJkLx6rLSOZ9kqFBLrl8BbG9Znf0oC7t8AHs7syFPevOlsqFl5JgQIe
isL7zMsSG3dY5XAXLGf6rgw+ADfmPi9HQtT4LzEz2nqQa6CLccl0BVb3aqSb4tnfJZTuPcio5Cmt
Lm7CD8jYHTwcCRebOZYv0tYfvvsf9EEgKPp1gUQj5NUkhZ5z7DUHeWryEnkdZ4NZ/UohUZqaDc8d
KqS35Qu7GfkMjpWwmbkIKzupDYixGvBRKCyvPL/rVWdVmojD6QSkj4kLoq3BMy07m/UHwfgYfPhs
fUIgtm9esBtiCSxT3Qu/cMNzBVV1X+jifdV0tPCbWzgJ7FSpfuQkulQ2D5I+Q9kSOTIRqvHZ9gQW
Tjtp0tI3q4Oe5qY/PiwwXJcYOCwaXlW+pZ+IVBc8WoeJe+UHc5/8txPiK81IatnFH9wlXDWXKdFN
d4k5t+OGHIx6ib71J5DtA2E2bUYFs2ogcPjidcAsnlKIkNt2lV3/Rn1Hku5MT5nfY3583wz988iJ
Sqyp55jP6LVImq1JiPwbR0DAaL8q2qqQzXl2Uj4BgkRVxJo9qb7Z0IHCSNfL0nfBYExJMrFg6fWz
As0NYAEzBJuX8patz11y+6f7gsrREqSxQzPUqeu8orlVJ/jCSzp5P3vmt7NClReUN8VoiVzgPCC5
b3Zf4GIi3FVyjjhz+64gWSyCY1N6LUBILfw/MsGqujYGui/uzRZGMwX4pCfHmo0vviVBEXfdSRww
1Ed0nxqTo26hKBwTq+k2p/o86jl+nAZmWfixFKFyM+b1Z7FE3GaLqJKAu38Pb7ckWq4qEQ3zqLkp
O9UHTi4QGxybsIs2CZ/fOylTp+P7dW+xgOYq8dxF2UlYfiKQ7QB9aa5mIVeoDVbEFnW2pb1OnxZB
GZkXBvbNdK5LF+4WPZW54kqAm4g1dYZ6/sLlQu5G0WbleP+jyF94CF8dba51q95TEKW8G4S2hfCT
k4WaJLCSUuyopyJXVNyxgcLDmXzrb3UwEYWDcc6LCV22fZfwT5qlexXz72QZ7mXxT9iTAgU4DKF9
6OHluD8OzBq+gxuZRnxLQO2bf6zAfnmmQhcc8Vid1yl0EaetdNXmKv8XZMF7eP6jftFX2QA19KML
q2RX7GIL8yyLTaHYFi7ofS+XygvHaqDvpAAvoTN52zT541JUWsxumB1VcAulOHgXwMODE/1pUDcd
uvO9XWdhKOwx7XzZWj9eszyesmkxws1Sl4/FRPLkb/kU+BsjGgMPNx3AOdnfcfgXXQzLKPMnuKGL
OF6Pu6c+eB4iwntJVdD3LIVzo77d7Ht+dDcQF/lkAqujRG7j+s+ULLbWQ23fQjB3NsRqZHABs/bK
4NEfxGNcBDQwq6JUIknrPfdeupwKHH741dBxX1Ln7tV2PmAep0ego/jd+UBfrzb6j42Quv0gNg+Q
o0X9g38qZb/69ypG2DmgYRmw/YrqllXoFDAZYwsolp9Xfl53KgApFAk3ZPzrSVMqNzVPnDsZQU4O
NzKoUfes8A4c/PUzHQsyqb4BzMqRbfdQSyadXx75BfoEOnktBlgcKwL5x58BPsZ0/RlIvaMkXjQ1
qLPenK4ljwuw9d/KWIQ3uNEppi9thuIb5FM465KSUrIpn1u9n9fyx940F7TFzEBTuSKKsKHtzvfp
ZwnPfzXnB5Wb2GdaAOn4q3VdI66Ijk9hUmzHWz9azY+rKAupHhPsVq8aXpRodx1IH1ntZF1Wz9BD
8G3Z1qQ/uMM1DWQNZSiqDrYv2IjSqOEU/8NVhklMFfuZATi6jae0AGVSHxMwPeCVogj6/9ALqwp0
+05jaEq7oHQzH4PRZU7CLbWTejJrq6WSNrRH1kkUyuOVsjIsf7j8ul1z76UfS7LH5ds+B6h8nLgz
2FN2FiMCu8K1mVipc8BtY7hZVJSOQMmVTBp9rkv3PO6XLbt1sVK5UCevjFOdsL2GkcPLA/QpTGGP
2BLZk44t1ISpO1vG3XhuvoRB4CLmGp2u7YdpR7REkb0cOFGBo90EEf6zsasMpcogCHcUbBpdoZM2
eR8xkjStTxWIDSNx9bhCkzMsE/8VBk93PLRXXb+pApfX5Y00ylrpi6luVe4nQGRHG3DojLSHGDJq
OyQm5wErNf9bATYIvfzMZrv0L4CnnYjz1ePta5XJLnaEt5EC/92xU62jypi7qTA0OH7O+SL3w89H
kswfMP2qv4Z2PWCNh4k/+d10mLV3DVg9zAZjYNj4Mduh0SDdnJjOaNSfm0wtv0na2K5VSz3C3DqZ
FF3TTSfPXiWp5y0e/GHypJ7fLFeVOuOjGtdNJljozmQUMtF+1EfxZ3N5P4UD7HCl2ZgojGTFmmbO
rH0gwEywLr+s/Box/Z2VC7RPat/woUybsv8L7cjkvpRzsKwYztl/SF8ZCGd5tHgGU5BkHBTzqmuA
aT5diMqzTlh0WvEHqf5kQ8ESjSfdQhUv7eYsVZfFNkHlTqlWEYET1rcCLyCcV0a11nL4ez4RH1d2
tKEBpOqcaaY4PKAsZm196IeFRQDetMBLmjc3UCPwGX2TW081nCgUxKjTz5Yimp5CmgDUUdtn5ntI
ex2EETfwS8lm/mRaGZJffXyC1s0YH+8nDZyy63l7RVUTaS1LSCSo2wCo3YrvNzKbcXyoph4RudWF
sFrOTnqa1BBuTdkUmPuupY67nTGX91cQbVdqmKwZS3RKTP9GeRIHz6pYH2zgofZg/C+Q2Ldn6iar
mXht7zEgREkMf8kc+YquJ3MNhB5fLMuM8J26iKblpyiYBI+PAPhw7SxazIsakO3XCWTQfmt1iu7W
JjSWKEW9VZkuE/d/Bkq3s/PYpHJfFToDrH44FFuxsbHNQnu1wjVnxICZeATWJUFW8kQF0y9YIDCb
l0xdHlrBax7KRNeFmHVzLeZ5r4o1oNjxV4oAF4MfTkfUeOtpHvwjB8b8K39cZEX3psW3k50zO3YD
DQOyzptG2cJT4qUb38X3CDNpHXvLbVgXuATnbLDPGwykKeI27iX5ioxX51aduK6xDVbGZFG2Ldth
cUYp7vYSKADWxqPXV7B+lJWz9gDQdxPMVEk312Mis83thZfDKHGl7sCWosJQmMNzYRvSxfYgqo8D
h7ir2IQSBQdvos5jwzE0A1708v5lPdZLRtM8GoKFVQXZpP4+guIIKU8px8q6N63HOg9ek0M3Je+J
vt+vh+iW7AqdTegIiHHMKD83sfMFgAggx2iq/trdk7WBDzDWuLdcr96/N6ulSSgqw+uSpuOJNuT5
7SgJTN3RWpSxTTq7ifEKKWdjgcuyVp6nhkjT3xKu9JGBOdpMIJD6HOJOaqnG94wPkOnbwuMCO7vx
Pfx4pKxuRZFTiaqN6TSSuabWx3nT2o+FqobaKCQtBUDX9MCko+4ft3gFetkwcIAmltNz7KHuOend
WEXtIt9NooxevsVj+ldH3j0TpgYXcLpaE8nqgf1w+Knqm19BwvaqvSdxQueaWxfzPVKfaCtl9NkB
c9fwqWoV0aZdLQ3HQJfCl9YfVtOMUupAJKBaoQH0/mRgFsKtRPaiVw1ofeMnc00Cg6agG20PenC4
BfCcLVi4nJCbc5Lae1MWaNhy1XmEyQprEVUWR671PYY+zjhXDNB2yP/RaV8KGSSYFXdw9DBqW25q
WJTHUNIAHbS25sLhxKdKu2sxPB9YGfqLPfKm9eJhvAW7eF5Bx2jfu/z/4dQ9U+0oh/3357+SbP1l
1kzZWSlF5lk1HmLFwt2g9Sw036DP0Uy/t1ZoLftHQ+si/M8+5Usp/MQ3hxDR7EfEBc9iex3UfU3U
rxMcKGuWdQaZ68HY0Jv9sF8bk6y/Mi82LMtaR7dGXQJ5S97NpzNAPRasJZy9v+gQcXZ2ARWpuP74
jpEXydFkl4daeSJsVPHHLX/pO7CyQclhdTQQt7/YnHSERgAUg99yQDjmEXQrj5r19gZdkA+NmMXd
vFBj1iC6MtGiCT3/qmrT68E2UWFiNSLbocVeCiZGPiVKeyXWmF8Xin927/I8BC9rhUV1Tsg6UpyX
0a4i+sZANV3OHG2Xt7gQ+uJN/+r8dJNz9JubkWHKKMRMO6xu8gC8AuFwwuhgiP5v4KzoeFbq57RK
/Vdkofat50aZDFay/8QgCl8jbqp9OuwbOKuHMHPDuwRBtGZK6uh5QVlTtrOGXy6nQ9XlZUQu6N8U
mYftSNkWpJsFunZW3wjEzcgqEoY264zGAUEWok4laVqD0lox6++qH6PXe6hpXjvm0bwpSKZCOnrF
bTPKUTuaVpQHNnSu7/sl1QgiXO5bfSNlprLi7PrE1U9xVYCTuMrA92R75xB2Qk82wM/W2jkwj2QD
0Agy+O/G0czdxnbbZJg5HU+fJvjbe6fGk1yLz3Kpynw7TL3aJaQvRMpBzuTGDVzxySAqLV++DojW
SSmkiLpk9yTj45HNISxAAh8c7FrZ5Mv5RURUt57CfxHYqdu3EMR74FlUbK3wbqLqYI414SNsNTqL
MRHc6pXcmbIfJgLVBFvOap5XHCR61WCE0GnNe6P0JMESx5QTRVhbmjSAwz/4ntiNupmUKAQhe029
y4vUyLqTxipMei3KFYzd62lTWaWzl05jbqs1E+y+s/YA49pkpivE2N+PpDHjMr95G2qcOS88qyRO
c69/eVAUyKsCUco7VowAp4dSymSrtRaS3OCDPWO272IR6lUCi/4pp5MQ0ET6U++QH3hp5DOm87sn
B04CalbQZduyPbIVVJWswQqXZDIzvPRufDwuwfke5TFU8Cg7xTsWufPfb8FdHvGT1+NcA8qgLLlA
8y/mZGqiiCB+55Nupg+sR3/XbQx88A21AUz8vJzYGSxtXyJH57PMxsR4SR6yzNkHCckESxBxaTMN
pBR+s9ZePkvviekubjhunMd+lpD9mohOwOJ1oOJuzAdjIPlIEs03sFxLDVBPzWJ1D53I9/Rkxh4R
URPmzRm7gvB+/K2IWgYax7eZFXc9zrv9OfMHCJvhbrZ5VvP74gTdtWqgLbYAQf6ZsgqkOUOMMviZ
1JTej05GOKJohOH0VYH1goMz69fdGvBu1TrCkV1aJnzmJvktjGHm0wt2/LI0ogdV5ly/gK3iXOFn
TkAHHpSSuXqcxXEiaBOgp7xhs7YAQMtT4UV1wz8DjHuLG3Qz3i6DyZdRrMYpRuV4kK8TeRqN1aEr
LYlKKNnG9ML83fFlqRXVMMe+cb26FndxQG1IOMDFJhcS9pU1WZmRY1BdmnTpMirowKUEFhj8aOsM
tvHjfgisKwp/Q46CrR6HzBadlRJGa3Khm6dLC0TH/3wjlBw4bTLH7guyhOAfUraU1PQbypu345Z6
/+0j5TzLxmEMXjQHIrGXbW/ZiVp5s0ST7bfQkmbzrQ/4bRgSlcSz4DxmtX6q9tP1SHzokUlk1F04
bAiCSjFSPeP7/fVl4GxgZ2W7ASwsXXN6DRYa4w/ZOAS26sRB8qzVRLc7q456RrIfnqgiksFKiw5g
WY/5ovueT/K1CNmqAmEy1Ux6UMWekzqCveb96imInjTReKey1N0h/H9Thx7aFx7UzDxqzJK74hLC
T2ey3EW8gFob3CIVAQ0Zm00K81FJg5QX+U0IglTv2Q7u4HanxzVSOpCQUbOqBOb0g21QbxpK/S3G
9ECRiocCHrkOswX+8VJIZ3xG+alEs7AuohzN2ammGapISrE5S0FupyMwnDyS4suu6kU+ILN8INJc
hA4s3XvRV+isCsKwcVU3F5WtZvAc8ahQHxKUqHAZ2F9BNrnfc/2mrMguLP5YmJBBOt7OJgkZd2yS
xpbX8kPTPJpSb6lMTYGM2+4Hr+K8x47JIu65p6Yn7TSySWXKiqkIEFqC8Fp6gXEQDEktTU+eWwj9
GzfcOs9yi7uiyQu6TlcHi9cA3mbw25WpCFgUhf1H7SQWFfm882Fchw1QQimmyFq4iSPW/UadF60G
LE8KqILzguXRarGyPh+Sk4KMul+O4iFidS7nYTefq7IuJx4SkI+Txan+fwFx8qV1K2Oj2T6AUIcI
BgOcsVoQu4JaZgszDRjXeX1VTWL8/rt0t69E3RpYkhCucDfBAFgCnaPZk/ufdwRIPwUs+P+Edmlm
oBUlgTxWsgNugciIG67kbqH8nZWWoFuWOBF22NWNDT8TdqIt1FN8VCQxvSmWMSw3Qaq86wcASze9
ciai3HUekf8IWKP8uxvJC7/5BlIYQaNd+Bqu9vpveeHdpI8WrPGfIjqdyuinoa+QyORk5d0Qm8wg
oHlb9+sIMcG2qxRzwEyptfzJslbULUl+hxSd5N7Bk4dx8BZAg0BEbfMKbsL6cYfQYMLcfcgjMJ9m
F3SbDgMKHCuyMfC/vPOKmfJ2McB7hpZsjfHulmCSQRdAJlCcfxeMMIuAmmp+JHhcsuILSJ4pQC/P
Y0N5EaQDwqdKoomS//DmGJOZUrMw1er+h01jRM/yg2SxsyQO3OAVEakU/1IqfEYq2QBPq25crFl4
/xm19zTRCPcdt7ihT3EYW/S5auczP1DXGdorhqmM9YQyHFNOUSDcFbp0jLal5AMdh5zvR3ANWf8B
1G/JIra26utq3W4N4Tiyh6TGEb8OV2uIBkNYrUZIwHkqR6dc704sIIY+nsPEcxSMcotHORU5gyhl
jXb4vZum3bXdRaWHhO8Il7PQuQsAQTg8vdT7SnUmxr1Fcjpl9N6sJ56KJbykjeSee4msZnOwA9sU
0M18VDy5N1Z+r2V+JQEgleaqNOxFKIpITxhRe59B9DGzT4LG49ZObLcgKnOSyZBEhDSLGy1MRe/5
ViIS6GhtcKFElw4FVVqQML7l/nRIY3ZAG2u/9wP2z8xoUat53qpkinpU2aymeFI0Udm07WLrzpIo
xDDvwYqX9gTgMSsu5+F3c1X/JpxTudu/szszAscDLOeTsjswCnlCvQrbTRbAOJNR0noMH8cJqPe5
N5ZO1nFRAROIr5amLeS5mA2WuQYIxYm5bYOFiTqICUoaAcUZ7DLSw9H6COK6JdBmJFNpApFeytTc
ug5GaYV7ZhhH3Izj6INqRqZis6aYjDZkYvcBXlkBW7J3mQMe9cEDv14n9raeYzbKeFG3JUIqWz+3
ufNu/J97zYw7081wKBio0HkWoNCoa9HeUwVxPyri1J17NeW8g+WC+jhhbtmt93Y8FgHxQKx2HuqV
BnWzl/ObBEO1dQDnnXLCb0RlNBLjkivwgXxqQxphPv2QysBIQh/QbxHmu1lM9kcVVh5gr3xXokXk
gxSNQSEZJ58vFCFf+xiPi+ZS6O1QxXUv/Kbo5uyVCnos9c9CcqIWLiBdwotljuSVDayhjJcrzlwV
kjVvQrfjZYToX9GbyDMUu6VCnu9LeGw2tQ3xaobV9jyGEi+kYWFg9QiyA18R5dd2aavkRzRtbgvD
+5y9EYYC9DLhzG64Pj+rFfdAipgCdqIywIwMlpTKtePsZ0e3FkbO34QJhIuo/xYqlLbaX5hbmG2A
CnUFtPGD+pwsOTIMjf2o9PyEfeIG44fYHZnuTbrukSYlEa/Bt1IwH/Dq8XETfjErUOWFj5EyW1sr
TOusvfQwh3yUzt5PNyZtVIUDpncUZdjY1Xy3MRKsWcgwwU4hjQDxtKpR3iPB5ji9gbwzisQWwlJj
m+kBtbwJwHqc5NyVN/xVpzh6gGQcbxbGHculUfkeTlxZVTc3Cw3Co6E3TxGY43/44NZvZXEpNqVG
NYk2V3HYfQe1BdKIHFypY0IOXlMEeWC77xVN6Yl7A1t9+Vfi2DpemoEUPCW+bgIeapz+OLq/D9Ff
+AO3DrjzhAEHh1R1zCxls7o6oxb00y04OJVlZM1ZbvwLSWVov7XnKzJ7VXiR005raJB3gxnpbTll
BP6IWj8Sd1s99DA6fcZt2+MUg6pVnIvs+0HLECpjprdMc7psCNf4SjFwSAzBhoRNHwPPuBGMqlLD
fwGmlyIbIZcItAdptOtSJAb8mNABrTS5nDFJrRZccJzeWfAOUw7cUtpcA4PPO9YvXvoMQpQD4cr/
3BzibG/T6DfLttHXZ9LyQb0Ylukh1E496AIyILAc0DgaLsX9JhM0deyFCSmbR8+J/BvG9vuj3OUT
Ixi1yM5Tmhju2XBg3LVEzpOqVtkfGE5RAYeSUitZSnDoztFgxoiGoQq4wZ/cnUy/MS7SMrSSX+yf
KWiz0Ytn88Rgq2534XFe+77BwhJsDc5E9dHvER+YyBechp2KvTfdHLCN2z10JG4iEG2Mi0huXOt3
wsrqAaK4jdeLx1bFvFdzkybFq1jZk6lJHff2eoBBTTiA5CdyoLGCDCyvNl4irAyqPJGvG8dCXF9y
AeZDjAygblx8Rxr/ZUrhOQpjYHj1oOzSw70u8KuTpqCD189sZtcSPlI9vwFOPWgAtmh088mT94xq
XKhJsdTLGa+JWrIpzzRU25gnuvUaxBNZzWfAhQFdkETZtM7yOiYaSinAiYgOZuBbRLu3lEz+UPCH
8AjWoccRLkWug+pluK8Bo/jnzFhM+sRqWPKyvcWiaF4Rz8V+o0gXAGmwZS7vTtSUDiQI0ZqZMcVT
8v9GrbZHXIaUvEuvET/FgBkcpIGEMEJINhsg+ayi6iMjRCbom/QrnmsT1Ht8pyOIOrE7dFUkk4qy
Mz1+eLxdrjCSxExiLxnlWcp4jg0R04BeWm12mVtmx9IgNpVf/Vc/hL/UuVN+sfrzuMk//3Hllz6o
/pJFl26IPZJza9PiQCoWxu8IgJpqQiQtsTs6MNDvff4Wu15JDJnI6HEZnm3sSvlM/kaDTptsEAzf
XydxTX4NDvm+llIZrcJqEvvc5eWfLrlWOtcSYwa3DYI43GjmVnRKMeIUdFyJTzOJ923uSBINQUZW
iDtA+tSeoUHTRB8nxh73qO1249KEnQ7fVH7+ScEroXUqfqTn4+ZxwIifxl0GwjAorgNXiKHLRmoo
Sdn/nbHUqfIOyg727FwDzGKkDmjDiRv4jIorQKNxStyMyX84Heztk4BYsVThcuJytaJIlrMPXAeQ
HVjF6dCEcx5Kw3tecMV+AIXhNmw9Lxf+IatKcAnTrXFn8Rb4A3ykhK3mLajkc6MbKvwxI33p0gQO
ZXROY103BAv1tg1ypmi38SmbVL2dooWf0AwadApmGJFkyi7Sd8EVlF38Msl/fAAkvCO3YbQOC+R1
UokKX4Klclg52wDvpnEgDmIlTbYrpEqxflrdTDQ0ccuxKHMyX7Y5CnAo5vPyU0vMrqLsWJDA7uQ6
Eizv55fw1z5jYXvp4hV/ilFTke3mAVB28+zFcgod2ePPv2qhKkv9UC/QCULOd1xU3YSqGtamJaTg
D9E5dNesVJOE+CsaykcvxFhrb2fNVlc9Rh9nTGkeO4sNZ0ObDw+xJiMdedXm619xn2EADu1G9ucO
2cXsdyMkISZW6sCN8bBOqRDl5dLcOTHcju7sCcjU7jdXs5Kkd1HcfYXcu8XA1gqCEE5qEIK2JmzK
n3OPv3QMKbJG50Tn3WKYAaFT8xP2+zNZFBpDfJb9/6fJHcoWTHR76i1lY7myMC00wYtPn34dSwYZ
FscTUf9JdMiNFq9aR42wZxSjXmd4ecdFmwP6DXT1NN7ZUG2ODUiIp3F96IWr83JLH/7vQf2lDyZB
dP6uwGf6QWCPDvGa5Liua3m9MidV2TJnmS6YNEMTPPAJZzNRpX/mBhCvTyX97XMAYfMB2p/n0Etv
jeHo4VY+KzJvu2duGpFn5PH8mCU6gP9VH/lJILrvTQbp6Y7dZoBe3jIFt4JIR9byOCgJXFfGFn+k
gyaqTnhrZ79dAmCIAKKa+rertg+DIWbWmp4hGfhwgX3R3BTSnWpt2HPx3WKQc5D3vFnmG5HXwx6J
MGpjZSCHgz1969fkfrLKoqY3QYnOnYh6jCuDaXSPuGdnJTguuJRe3keBLhusA+WhPmPamXxR1qx3
KHoipC6bXJN8jfe08l/nCd25xdps+DFwgjt35gt0THaXPURmRj5nzgkAvU35Tz+1W2RRPcFUOcky
1NszIkDdtm1q3pcMqWr022wiSAzL6G2mGcaHbNYiK6I64XrxVOIrLXiqEipmqPolJyFb9hgonZCg
rAoBMH5Cbua5jUDn+tcq9D87g3qvdcj0L/gC6EsIr94estTzV6W9XGnNK8tNk7T1s5zHTc4pEnKY
oHmkOr2YbCSaSHNgs4+Uh3hgxaygd1F5dUYHj6w44puRHsS5LMGDkTkRNmp7zkLC9IZ1Ir1jwuWn
VKWgNlq89sH422j2Wz+wrZjWUvtAaphK9NMIljbqAB8nxkgP/TY7ac2RAVz7Vgmo5EWiuvKxqRWA
gujc4nEL6nKv7BevvRIHWe5e5+Fy4x4nF7iZ8E1kI5pxPtckOJKD7pikEQOXfmyYX9gBj88JnGMY
PHk3Nx0gOgZmLZElqz2KgJaoFp1mOwMChI46gMqTGgKKBazabHU64G8MpzPBICtXYmB+68XBZj9t
RaM2w1WXvPTLpcpyS/tTe3o/nJR3dsBtyWEADXRj8KsVgjKPIenPuwEbE6yWnFvVfyxZlOEoXXcD
8+1iHwjXB+MPh/U8gyXz/OrztTMzrmTYeweQq2+1k39Oi3sAage2U5mmttz+0xDn+3E/oKylMTth
J4vy8dga9VITx8EdRKXvdjrSjY+/0FHgZy2Rbfaf/bVEV6jAkoeFiL+lBy71VZ1F88xsENMKmAq4
xOWaSw2vALYfJlMqFbL5WlMNQwLkhkmiTioOa/eqaYBbFIoP5mT7lZY/E6NrLu0uX4XqC0XhtAMM
EiCeFo7uaW0wpG76ZkjqovwJJzf+hmaK7zrdFA32j5RnG93kaAvdeiGrzivhpxBQnPFRoZjHP+7n
3Gpo4oTZt7fjPIY3wa47obd6k6oh8Vkvvabdm6x5Wvn5T/Hc9CECA7psAmlL762crouts4uvPyzF
TsQkerkdD3eZCahGE8Oj4vUGIydqGXB3HVIaOucAD9Om/bTpW72OOv88UTD2C6zXBwihjcNqhtJV
eqmqJ+hPIOHro4elh0zZms3xsooD5xazKYmVr4oGjwItTqdDE4JlTRSnzIhWSAYd+86/C6EsHUNO
wyeNJ5c4rUNUDVLEjZYi2jpYpZAmlh1863KLf8mIee4aXtcVySObH3cnOk2b8HguYxQgGL1zjTsV
1OQRzdYakpde9FyWmsp5k9FknQofznYPD9sNsD1EnRts663fNLGKNbY22O/sEDc99n8wdnaWVHoY
FL43wJeHWEv/PCM7OZPULF2bA29+J5TuHZQ8nFYa44CfVu8sF024dYh4WnVLMpF0A7D6qWNuB17c
EFk9WI7UPuLUEg+EdOrXvxnsHV503DUVY/5UoxE5KbtGq1y4CarUwt8m2O7/F47B4oQZQhGzY9Cd
q1S9jszpzVknlwE9b6S8hY+HGibLX8EI2jApty7Is2l615oyei+YdeKtcF7qjpqgnH1rREdzP5Tj
quHpIaJ7Fpr7L9nj4AnHf9n2OAocDmR4X/h3tvwK8jd64Xlk1L6MrHdMpsqQlOTiH/vuFW1PfBCl
MARg9a4/jJKZD9LZFWu95vb2VEhxwPAeOJEVsotejPF7saIEkrghpAX0YQqwx/YAdmZfpFlb6Yfw
Xs2I+KER9hIq8gW9yPfUwpWTe0ZqlBTJxAQyLgwSqO76K6FB73M1UoFlw1B8S4kGSCio+lMRGf47
7KnK9JNMRG4TUpOvSFoBShX88IJLv628lt0gsy/at72s/vBBaFvZPcndnyQySDEjxP8X4doFM1em
GUoyPYpBacTUgUdNYM6uGuayJlwqHdwlagbsBcBlXDPNzY3ICaUuto9Id6M2vQcimSwo+nnLj+JS
IaHh/qPqJT2mu+0J6Eb2vkscWiLS8Ysx7e+MLEGvfrrvwYqnoZ+OXPrhykQ1lieAW/hXCdJP4bhi
w7FLiQ2hwQ05G9OZ9x6Tn3NSGTmOrpZk/DVNHnd3UueiK7R8S4lKpjCFFtIsHdSU3trPa3uDoYZx
ttsxclmOZltynv9ocaFHCaTgsgapZBVOSm0MOvZXZLwty/R3i3uFQkBNBKbBDaayTKzhBA1q6FeW
N1Pj2P1dNrxPVPPjJPn4iGfEcBEHqEf+L2W+OBDEZEdZf2C/M+wsSppjzeT1dx89MF/9t7SEfPHR
5DIdKyqMmq3Mpz16aHz5eepZYW0DjuahMqqI8kFuxMpU5D/EMRQNV9OgOmS0kU8rw0JEF78N0bd+
cxaAMOhQE+cW1a5XdbLoOuMQI3wnvRdzxRs+gUUwVmceKxcAOO2zG0b5PdnnwN8Wuehk0ho4e15e
gEu7cWp8LL80J6h5OXf37G8JrSTCXVu2S9jajFe7bvd0V4fzNHA8dr8rkNuHPAzrPDNxCF97Lti2
OLWpMSQ4/yyrUUhPMyaUxCV+HcCKPB7rgUjRJ9ibeFsR2HCvZlxeOBV+y0rAIMZ72u0cGz33tuDV
90Bx40kzv/F3G4JNgYyMXTF8SW73ta2p/SghTDaG0wl5KnXgiMzVG3IULA6p0SaUzq+JxgD6M5Vq
oJnMIsEPTkH7yTQ3hrJiqe9Md3aYmBOrHPAq//GRJcthd506+uA0Ggjy9sBbN8wOBTU1j67g65RU
qDpskZANxWOFUy6UgwH1Jv4E7VrKD2tmm3ah5/mb3Um2hb6ehQVaq3hKNUl3je7tMB9OYPdolqis
HkluUqOO3Jpr6fKP3usVrRUhjW0e1SLmQ9oz1vdJsXSiud7cZoTtm7wENmqTRyCD6cUPoFkOAOMx
aGaceToG8rZHpK7JxRBxH/02/ckDeLpIv/AdaX2F43YSCd40vHG1/lYt5rjNg8I4O3B8CYVLsxO0
H40bc3HtyntSnaOPJVjOaRTJFei7fu627QoWOTjdri/1ioCufYHGcqDJleqEMFPq22DC1aMzBxKq
uxS2hEkKc+Sbf/9L7/9BQts3NyVnqCE1qALjamQ2wF1bSapqaMpf7VHy7KGpCQn6nGkiJPoNrsi4
z2jYsNP12HzUPB6OZr7D3rR2ZKLtmAm0l7zPHGC8XIQLoDJg4rROL8WwsAqSDz8L7norJbSU6YBM
4v4/nEonh8fNtSrAVd2RhusUhErpA+olXTY49vSZEgjYsPawNjZpOUqYHzuUwvwMsCfPjWIhLwrU
WpYn71edVoQyi8dDrnVRLu7rLGlGTNdoIZoxe4oqGvbU1Er2TbcOyLqIOiuAkYyk4QlGsLL3Ox88
OMQV0LR1M/nWDOdAEVY+9cax4qkNsXcEZCC09De9eozWgpv++HzKSERqUhX3Zh3Hf4t8c4sKu5ol
hKqQz+N4OTtNngtoony9aYp3JEkhQldtnnOIIIpP0Te5BFmWcLCN4lIIZcdOOQbhJV/5Fyd5PzAe
vdtnQX7Qw+IFQdrcLC5i3t3dMSyIyWP9Fbio6a8Xr5SIoYkjMXQB+zpuOQey7uu5Y5+VcfL2kvC/
gUA9YRtvfDHnhsUlqv2inzHpMa/Z2kI2+nP3QEXnzcqg2syGGhoeZtVBqZJTGdp1n4MIhvjW2ll6
QM72l3uqSZkz9GqC9Zs33HkRvC+hG1udqSn6ZCsHFfQItVqmDWl18bj5WHA/kmxgHrW6QgRZmwXP
LU/jTsXpbvc5BFCHYaleJ3l0EsO0T2zZxBTqBO/SsX4YStkBnziweL6kbjatbwqfAOVMP1lqjIrn
sT3NP2f6RpbXxZr68Wrw2dd0X4xh0F0z2d/iU6BcEj5S7LOE/COAul3oSz1MI/y82wicpMtNEst+
xjESf9Z+WVihNynZZoFyb/pi0fmo2TfNMxX9TUyGoV0iHWD4X1ooD+l8OdrOsmV0X86JOmaPYYOM
/SGLEjShOPEEKa+zk/Fq6qDbCeAA5X+SGBjygSQNKAQyLXZ0klAFic2KYlqojY3xTWC7TXLTtshn
zAQOObgQeZNTWlFVyWJ/hdI0IfT42ZRlVi/DNKaCfkCjcJXYXsElqNukxWHhh9HPTyPYQq82uinS
7Ig6CFKcg0J/uJ6TtiCcAJoo7sbRM/wbcg1OHGcPgeiEYTwV88pg4FK5tkt/kTmZoIDn/mrbc4Nk
Codyn+zYxRLJqq7oE4A6JiYkDMugBrvvHIUdrjI9qV2WK6jwjOHhDtP3/Uygi4q5s/SgeuEcrif4
jgHrJ+EqhLuiIXMnd49SowXunrZKZrgG1t9Phq8onT/xfI8sUAylxhm5e7ZkdTrftvNkRtP6bomd
vgN1vueSc+2Xd2pIT8zmGb3qNtR7Xfd/8Kik6laUYwXRNxfTxx2qgtFOT5+h/peugq0r3oWQOM6d
HaJhl1Uq5R1y7iNJz2A5p2FrhO6yOnkv6Avi35IUk4kgH1m2Ak6SWG+heEELmV4AQVPFj0CvAWGy
pR07QlMM2RlkweSN6vuZNf2Bpk4Fto7sWzkljrzRr8estsrSziMxb/B8oWlTAjgJULYFAQeihfSh
jtUqGA2cmXhXp6OEPikW/9Tb528PwTNWg0tzA68XHnVgCmZWCOtaUQSwC5vek3n511C1j2EpED6f
AonHPHld+tCJq4bU6fsrrR/2wIEmZD5uUvBF+ilzhszMmCKEBxFrA2ssXIBtQCjuK3CfhCxhDR1+
9RG8RpQ9Rku3PCK1RjHNoRP77Re0txG7y+QZVYSvo0y5aTAeFp4VFSFwmiKdp9QIej5QJzmHq8e/
nuSxKUj1w/x+nWERMnTmmIfB+DsYsqrmj5ErjaE+uEXrQ/VgASist4GQMXPz0eS7DDsEjM78LPDO
ztMsl/r/dvQTupS03o1Q2Utkoxr3jsufs1wVO47Un7VEwPa4nI+IvFhP8W4kx8QoUztDfQ0oeMS7
E75/99mXzjEZ/bRrUZNHiSUFmlEATeH21WKQMIaVLWcMTQfmT2/ssRjmaI2c/UB0vrNHXyoObpXA
M67jYy3FBJbEZjVY8O1OkKsD+FPGvrhJVIPqC5Xgt8tx0Q5wgAseuXHLrrigf2NBs1BjB7iUDvag
ZgjM83aXJU4+OG48wazkiFwV4GF7jN8dwDIyuTzJWK04k1diuh5CygmR1BnERSLe80ROgo2xM6rm
DB+XoNMOW7DY9j7JGNWd5w4/QohQKIdHCoRc6wnbD2MHW0CClKwyz1mzRuXXswLx68BpaRRFBSSs
XI04RCmVNFHyvV6OlvdX3dC5FQudVeQcqgzcA7OJzumwothodoVL3RRxNEM9KsQc/l05RAFl37El
eaMBBvKtq8cc0BpuV6S1Cz8SF1ekZMB0ou3f9ebqZb+8zwX8EYVO05uhtxE/+Za0TJwNVNAXme6V
k5aDyNaesHjHb+yv2rFHog8dkrzig0SYeE2MrO6GWhy/WfV5XIhmuaX4iCw0OaHloQ1MnaIcsbUp
hWsb/zy1Tp23Rei6PGmNBfHEFNn1uuTdf4+xokPReM9DUhnTOeESrfqmgMokPbfDLG2AhbFda0E2
8u1yBF3L3j/Mxs5rcx1YrlobmpIOyNayGNoTE6HlJwXtmJ6t+7aVufb6KBym/x2jXDdx2EogCfkB
EFYkOliF+i4mBsQnhSMP0pzEl6JGYfDbPxGx6xQAd0+xwAA0LlSbhjlx+Uxu7fq0rpNlRDv1mHgk
eBvqdG54dn30/SreNvRY7Znnflb2zHlUwf0N4M1pctf9VL1bL5GlcICbSk389bJhafZsk4ker4Gh
zlKGyW19XkJAM7UweMmh9XCHy4ZMwdBCfZat//KF8Y84wZcLjwPAD/ggawPNHyjkwN7DU/eLeL6X
cy5b2xk5WQmVC/4zSpFPW6VL+e9qJtD6gnu9QgQUHwpH9Cen9NPfP+oDSIgfCD3uSuJ6wAy20YJ1
0xYVrhbOxe0SsB3e/eACi6j/1b13t+4m4mMbwaLQncNerBZTzMCH1/dN5+Q82I/BZYLaX38qicCM
nYVXv+9AftUoSBO9NhgXAXnOlbc4sDF1IrX9OiqmHXE/nmhAeJ/wbP8HRbWeqQHhsPwfau1P+Zc1
iYfvWPtGocBvON+o/0uDJ3pFmTCDK1OvJvbXAAEg/jxE465qvqRVWfZaO1s5oUbYpJaHHxaDy7HK
0RmV4gpoz6kFrvNoNozzzeJbFy650W4XG8UKIW7oBYoE+BWMZ9gXT0ybaNwuY0OOths/AQFByIO/
FGryS8/t5gvzpZ4Kl6a3fsqK2nMm8QDhhMBZPGntGlP85UO9YFmS/dUIVdrbN4mxujN3xgEZ1km+
ehJWUdyev+BtFMRmEe2ENJ2LqaDnEYmmy5BFSTRE6UYV98lHsr6QoJZyCZTwsEffZ2YGf6c7yaZF
kzmPNDndIY7SeSJvB2ylK63W78VPtNtwW4t5FPLONCfE5MQ0mO7iCLvpVzWNyzi0EMFsJUImw8uY
oWAze/yRrxrRq0ETzouCJJ0roHL6yN+wKHOJC1ytxIcNSRs8gDKg6W0722vB/rZG72t629DVJnC5
NcYPc+5MVDIR337fIw80/TiqAdsz38gkxNKwg+pWwhF3S1VkanHMpKkp/6AW/lK972Qwx+d3DeQP
/26MGZ8pqJ71aoZOda87l+wCVs2IuNIXdrNR+xFze6Xqn0C2ZjCN/dJaFoHXCMhITB6r5B6unrIh
TwLBX7VV+dtu8lWwvLANMrTqnyhSftfQarBkH44d0lQRPllrYyBPIPuBzfHHUkuJDmlJjVI56Cc/
im0aVDXwt1GpH8Jji2i+bgzOC8y699qeWM/kdmJoWNHQwZiNGyBFD1uL6In8afXvvlHgtkldVLjw
duzDHsVmA4c3/4XTiKKu7mcsLjtlCMB9gtfpHjkPQKOt7J4BNaLtTk5cfssCmg0LXnvCvNTnEzWR
PDCp95nogpuItcV5jDUJ5HI+N0RmzheMQOUyt/gJfELR+y+neD331MQsx3QjSAR0W+o1g1d8yj1z
jR26t/vFTjtFEhPl/7eqvdOMSy+KGRSZDpM77bhvNnfJdLmdKhOCf9iORe/SFE2mJprRcAhut/LF
OZubpreMPORgSRZ6X/hCeSDD67d3IFjSfnXxrJZJZQMw7AxrLjY0JbAsyNnJ+7vkgznMAixbbSuQ
i6zJTTrpOTBQ9t2bJVpe3W4sD8Qsws8ITJ/5MRC6ycuIHw6L7LydTIQcMxeWoaveR5ID8fqjR5HO
a0ylUvgdkds1BtG5KV6TZ+tfLByEf4OwWDEKpOATtbj2U/bd4Z1vOWCdg5CbsS4gX2ieV9G9zuvD
5vRhmWiNM3wXNVN48AqvEuoFjMNzi/S4pbCyBCrLELARhIN+OZSJKXk3X6QRRZrRyCqVMtC04T7k
FEAwPXRmaI/mJWwdLfBiZcYDqKaNGu39pR4tJqPl2dQJCBZ9XWWva9m0FzOpZwXMurmzM8dgG8Vn
u2B0i5FA/DmbnPgEnmzb1SXBieLpdxJCWRaAx4VAvGGkqhfwAK9FIynpz2N/OlrDvgIkT8AvwmmJ
uesFo51alNshDKywfMCafgFOsJQk4kPPnCLNFtrHKXUenfiwVfaMOfzSGI7LYANViUqRE80siKd2
zgZe9mT6WvUNOg0XGqnotyV/Q9SL0PRYKu3D1gJkdUCmnGRzQNo8vnPJsJsnQmR1KqMBMIE8PFUm
DFwUxxAASNUURvjyYVX/SEBUemE+A9w1AHWleGxaDY4RGmmW//a3nQcybAa5g5ADt0/pTODUOch6
BxaqAG8BbJGVWBfbFRpDxGApATYVROfkP7tWhc3UJAmbJthIfltdTGVsnjrFHeYPTM8y/phJ7ZZV
z0fcwcRjkD/iLTIuHpJg6/f+CFp+w9oW8Ix/2RdeQr0fETeSyzgBOj7uGY8Qt0mJmFKSs/jLq1cf
IqCIR6zDPhWp1CEKg7Dl3wHe9hsJCxhg+CkOE/WsUexbApJfw6nCAYikmH4i5OPeXHgil63Y241l
w4E0svFWf82s7ZGR/K5lRZ1PsI4m+oAwsQmcB1kIkJrJzz+0riZZeeH2ZwbKnQFtWq8yRucswO8q
SSHapto0OfEaylfJVO/aGatk91xclI/x2rbCx4vJ/wiVPOi2NJTOcOvNLJq9kMgbZzEiiHjmSLV9
IeTgithCkg+466+p8LvOnRuw/TdYgQcgIlxgOtEgoTS2vquEmRiXq5Pm7OfX3qcXI0PFXKo+wZvD
xnpVXkcZmEc+mQ1ygRkEq8w4qnFx+qwktWrSArIIazl4du6zuLwMlMQMcjaVRfqxTt/gEhzYd/+x
6Gxozyp4cJxeLleG+cfkSivuxqkyzyQt42NtK7hyVDy6XTruyP/gLmKcqvtU8/Lsks20yRUhEEjY
s0HNInWx0/olM3cgwVtaIIWXc19abZsiUm3lM8L04+JYj3DVSD/g4c6xmVb/sop89vbJgXWyhDHb
n5d4Ach7mXb4Bysfb+ZhbdrymzkQ9f+U9BJr1qLnkzM6Q8xiSZffWVNv/Fsi8XMshNiLoufnDqtT
cOqDdA+DrjiUS8xYbnhDCq8bCzf1Sf9tKZ0ybIyiqeASTQfz5RtlYwdbC6CpQ9a7435MYwDr8IyY
s2Cb8up5Zlc582zeO/f6GWQTYzXdD27WBWipLRdzDtq5OLamEiQapFne8/JVbgVq6VmsjLMaOxo1
xWpCoMRMxChWvMy1hQ+m5K3R5niWb/hW0sPLmDNvFybkVHsN7vHN6wy7CR23Mc+/eQfkwnTTRXGZ
Ozo90h1FZXxipNABEJbpYneX1vi07boZ9iMmRj5OD9J6OTodIOk7TrIQ5od2hg6m7CTPwAW0KWVQ
h3sv7Ii89rEJ5Dt7ZiWaSUGRGtMDiiQXduMB5d541+KtQtZsoYicF1K2qD4PqCzo08tmoBEF4bYO
cmSnm8s0spodhlaeANgaGJpERh6MZUz+p3TOmLaXkKl2XEg8OukzIzxChu7sLofCGAbup3oihfUe
GQvAmoPODW5TrtG0xUW/jfgYgpoiK5eujCb5gYeo7ebzw+eRvRWvUEoYUFWGFui4L+bp0hKCG7ps
58uFhn6b8DrpNB8bwBd8Fr1r+yJ7pU6MVb8xqsmqi/I9ikmmK76GyJaZWuYs9CfSjJbRhSUEP/27
c/TKDQq5sYRpjSu1IFDC7rQ8tlCGXG6KEv/7L3Vjds13tOE4X+x0vV22JRo3I9v57TmPDddj1GaV
a4raCtqTNGRHF8sFpiE1aHcTQuURDjbWzS8WBfpa5wRHZ+tNrHgh0PhNCkmZPJmZAoli7gCXGLTK
3VaUmyLpTYTLCDcJwl9+oiTjTNGYADZS78rAEwmUz7V8IZEOgA5KRJbQz5vBvMuEVtFMNoYjhlvE
6LgWXJBPMUjzXu+nAkbSBkapgIiB6thL7TLxudHp4umyqqFJBVI1tqQm7bMCgEpBcYoSiBI5yOM8
m4l7ysQhTtEZ2fYn4QNmNcDYyXTRKjrSNxsdnLuuAvm8a7Vfb7ZSCT78wfxjTNMIhQc56JF7kinS
SlfU673ag6RdjEFBQ0o8QSpwjXbh4JN42kyHbaRjnQAD3nT18f0olCNyuYO+yVhTrQp3MKYN3FHE
1SN2BU6D65CqB4yTg61E/pLJiBVx3OlGJzkaJ+/UFtH4a/nk6L0ROLtCQbQyoLPGxAGX1rGO4MBH
rClEo5M6tIx3moUmTPF8maP9gai/Zf9DJ7EWvC92duHurh4i5oHGp6zX8o8sY8P11+Elw9dbOjis
1QEGy5oFye0ZaJTfdMG0V5p5SGnEIfIX31cHrNNkAo0WOtdUHP74yqyAc84QcGbdGxdsutEQEnbY
y/3xKP7HXRAxhpbrPVKbxTBqU9O6C7Yttk4lMdFh+6eOxlA1cy3BDwiyGH1DJgUFRKeQhR6quXdE
dOh313Acd338Cro7hL1CCcQOSwGmRKucNkTnvaNhcuzArsrgUHs9fSsZUmqUso4PRh1hUveS7aHZ
JsAufkPkAfphLH3S7BhgalORLbuxTKEDRfJdZI+DyeF/656l4IQwnT1k4CGFB2xd8Q+KajXMzMyd
H3FqeXaOxzuwo62oVA4MgcgGlGbLZqxd4d3TCy9YgnqQxIgbr4G0WQJJUbqIr6kL9DsBY5ifgl3p
RpTw1FNknoQr8OfXT17qIT1eVee7ON/wPKWddMWg9QuwcicUJgYWQJCptSBp6N9h97iunoSleE1s
ZCZ0brMgNnSRJEBLXcYmuiwz6QsYl6Rt26p27ZwYB3FSXc0rjTlwh0XcDIZ/bwlpSUvlD+nhn1sS
LJEu3mINnu1VEPSCKGEcItxYrcn/eiX1Yb+VOTbeFwcOVug6DEF/jh8luLhHAGKh8PCIVuFYvL5U
lsTxX2SIT1DiVWzuJPUgljybCHyTDboNkhbcrqKB0vMiov7eyqQ2eY8JG0z5cny0TRqHHnUycOmZ
ITVz0ExmWJCKTgAehVJOEc/ms1VP1sXWO9wCYKxcjR51JbIMnZyacCvETVfvwrVxv5Z4HyG66KQO
oo2rMIILQZwePyZNwdfXQKj9K95YjokoPUKYQ3uScrU760rW79NPWKlECJlbWUJt2SK9O3tmOkI9
OuSr0w6J2nPWJ9LFxj6vcxhhZNYI7g4KlIE8Vr/V6xYDZr+XTVynKzAOQnETfB5KsR50Uk0tXdsl
On9/+W/hj7MnWz7pCb5obVFlrybdBxX1t5eukPf2xKl27n5vpkAHrNUNTl/C4OzM8Ek3+/I4mAv/
/hcauE5/ou7/2bVU6943NklmCJQiC+OLxyWrsajCsRCqVynqwi1BF4L60HZ56GSZr1Wf8R+rIPBz
KM78qfVu9yDF4LJ9DdZHGuYlvpb9989A2v5HYGS4UdHCaXjT0vs0gvPubEUoHw3YRXcu4xSXpr2O
+OZWstW2fF9bFtnfgPFBZ+tJosASd0/dukrDOBotJaSOfKbYxSfcfvkCImVBnCmi+Gf2Uxl1X8nz
PHlQJCWq/wHOU4pcHeBRjvOG9lVT6PRN1r+qVLjt2zOGd3ZvxssOt8lKDHHUV3lhkRBbn+reehjf
Xx5t9QkUahm6HM4WpvJ+iJIiJ4OFBySbfzywpglBbxJgGt9C6m6JKQ6Yt8utVHfAMJ2C8nTkpiaO
id7ljzJyBemDTGSN6WzjWsTVCkNWFXvOyLVrHVqYFLVFBbUFrti/PwOpj/c7wUksHCyjzO5FB/y4
4j4FS2viyI5prEWFwWM8GEqaPeZBoMpv93qLKNAHxtUZI52N4pr6OYfQ5OID06JVPxbrCYbmv66w
moLH5EhEG/h60Xb/eNmXB6UNjcr7sNNlbY/Wb0jwIg/lpNn+m6mN9+lq4u6nEPprGrhzPBEZGOaj
DBuu9qVhhTzECmEE/pb0wVVEkwt/jieRRBSKaUxcB3AbVHSHYHCtshALOYiAArntKAozb6jV0Hac
AVeQT19tMm6L6zDMKPFOzPVjrOhnK0wB1iht/Aq8fcloi5NvUZ+5/wiNgPg4jsHM9UrnowNKhEag
+gtpfF9Y/XqsHI/TD9iJ/tHOcmIFKLJtYPjIBKc7mjBWXD/1wxh9iCVX/zZCw80aAN5ko/Fh7TgX
g1906lLsL/u8oE2dTUGWMJuQMzfvImsIumq2uxbCw2LfYeVCfJLDNsNp8JZONsEqaW2XsBWp2R4y
UpPIoKVpbSGz7eJ9hu+l3UmwOoIp8NqOf6IeCDqQW391GWnCRqMnRiu5YiiqVPdS9ubwjtQrsboy
LAs0NDyh8jjMysVuNNGMWDpViJujM6s940trDKvyNVlroiCXsUk6aDN7TC+5fTgpj9m1H75AB0n3
I2c9EHT8amPVxwQMKh83VyK06wHWdqBb502Zg2HnJOXFtQ7fSOpCqsy9DJcY16S9YqQ2pYakaJPR
Hn8JWkuDZ/3OEGiOM0A35LR4dspD3ofPQWAM2GG1V/d4RJWRmr5bSb1f8VvQUkobawqA0d8Q/p0V
K7R2p86+UeR4UGRkmpO/5lCY4DoK/3YtC3acqH6YONVLSsQZPTsXG7hMfyPHSSONCRcwW5CWKq3t
KfMK/CjEIlhXXOWpXr0bJRn+Qg0bhqNuNYcuR54dFLK9evLQK3ERggOAaGYd46JU9/dG0axYdPv/
hp5viGeP5YRgyKZ0FCkyY788K2UEbKBpls0dVuK0LREQWEnIh/Q4NEEMhaT41+qWdafMSYGzg7n6
6q8PcE8SFFSJeRIHs+OgAKns1dzfEEYzyMbwFCsj+VtpwMuslwn2k9b1CF6/BQZ/+XHualgIpOsz
jVVSfxLohw8EMt8rnkcn90gXSe8U5PjMMwduz1r0IKpwQzWnVx6JwrxVRhc2BXIq+20S7DBrLRBu
6KNKu5AQepTeUGyY4F6CT1Phk4uMBvuKZ2zDH/EQdxIrX07oEjZsUywjHDPNDEbJE5yTkHGd7KTL
lHOVm0lk1oX691QxJzIyMhHU1N/W1LUEchswodyx8x4FmZAtRuMSG4m1HFL5yNDhO64SMYFTmCs5
texkx78JpopnkNJ6LlcsZS8G7tmFNOBurq7Rs0aAXw5JA2bi5ZD/Sw3vfEzL2QLnR3tx6pF5NVQ3
Ezux1VYDfsYTh3SkB13pQlN9+Qy/z9dVTwJcGbJYUiHZk49yPV7GRaZ/8ubIj5YLNFM0rXSOebyN
wreC2+eVQXbYTXslGf43Yg/nUM3dH/5oxRT4Oz0W07AtvkYffAccTo/2m5ouAdx7bEZQYOt44uT+
rLH+GE5YgbE7bHj1tLOgz/uDBnV3eaLP0A0qAEZ0yJ5L9dtc9O5gqHxRZo4CgoUv1tQQpxQW3sGd
aTK2ev/soiSv+3t8UKd5Ijn3xmrNwV9yCnt8m0PO4fDUCkbFwD1u/+i6zVSR5mivqSx0NnEZGosw
NH9GlDiaIWCvjlpR5mp1/v1Fi2mm9N505SqelIFNCxMrgDDVf17DTFlygnGBsY9I65eeZ2dnEkUR
y/kvqR6QHMABQBIx5VPDf+qN3IBhzXLrQP/G/ibXfWAhfrc3c8T1jrpcTbP+uDOwtZjldSfJVU7x
NW/++33Swfvfr8jogoHEuM0dFWzS46dOEbrjqFGweNakyDelekpGZ7ua54Be8chC09+ZeKdmhJkg
O3zll+J8EGIJN4lRrb6uCENLzyypV0nZ6/XjGDGYolBdtvSX+CyFxjWITO60bT8HU+giJIPVSmiF
n2MWQFFtZnXmaHLmDQPnZEKd+Ipxw/Kz/AhnFhkMFcxiEAfNy1p5kHHynV45vElXLDUISXJ7zv4h
NE8zInphJEr7h2gx4uFGNQCoab8HerRYUex7pbjfdl7J6pisV0BktQn76dKHsn9PUWlQnS0eDQ+h
Xp/JdoWJmwE/U7zx21XsbGwCsOyhwh7imzVVk/dbT7o0pGqbokrZIOWgjfrsWZJ1+CjDUQQIH95g
pfJ+sSg2fF/+5fE628pl+7K8XMgV0G2bDMfJgI29KXQSXzKwkTeHCzDTmVaEWqwNqSwSJjd4Q4Ie
vaE20jcU24CuQbTf7Hho71OvDma3cS5gdo+Pq4VExzrZrV5Y/OMWnn7QQoaGnxwBmUoyTlOqdDRC
ICudklXma2LwbRdj/68nZ1qIr3ZOeD4H4ZAs//gvXgE9yFInjKcUmIobYFwOQqy4QYcILGix0B5b
P3hhgfpejBgCghEHeNbKnNo6suZ5ZYI+bmQB9OJCGbe6mZ6ORdl/AZTJjzXk+ahqnQuWbjWhxRqb
5SsZENTA4BKbVc8eNnmNEGzqFrinGiiYfRhJ5N4b947rpxYP/CeKaWSHWFzXZevEbeWe8Zfbki+Y
6LWchs90eR5wcChy21naKg2SaWcy7V/Zz4dQ3yf6/1sX1Y2wYLaDURQ704W37lavIil9m3AA36jS
i6V5DfjHemZ97Rln9O1wZSUc2jwADX4lYrOm5IZuVwGAdixWKHewP6RL11ieR+ISoPHd2Ssau6Gj
iPfBHjAUhIebjsdiDQhovUJ1s9W3c/BKZuMQP5/zF5K0jCXN8M0alVFbFjpXJ3MSWAXIblc3Wp1y
pcj63SpImPK9IUj7HsNaGZe48Hc545UInYOFn5e/QOz1ezS6iAcMdLW/Omas+1l71XABJTPAUMDr
55VaPsElbv5t0LLwUu9BrWJJs9KLEJA+ms14nlnGVaaZ2a4UBy7j6stNJS11j9tCzUB4HCXYHNdi
4JprTRk17p3vwWD/YLhAJQNzTCWeCLCTICYgwPwfSAcmHY7mSmszU63KJ6Xu2mZhOWahSSpBvGrz
30VAdPkNGnoYLLVwZQK9zRN6Ju6norPtvBHJeKLH6mlBjaMLCC2RWWs/tEfQRYlIwvi9j5tIUocs
f+WFigCXt6K+G/ORcTbAb4leCdeHpViIHKFfW/i9+pqmz4wEV78f7BiZVI5k5IPLPqLsu8AxG6kp
30Ka7kxCVweeuKc0cRd3mlDqHi6/FUPO4yCGMIVdG8z5SamapepNb/Rjp2We4P8HznSiB97zhQ3r
Lp/Ki3xnqSD6pIKFGJFkKT7Qhauh8u3sWU3VjVNjrpqjnl6gAc3deiY5CuxTke5CU6DIP+owmi+J
42au+n5HyOJIiyX4BKriqI8FR5rVUNjq8wJZxhxl8t/EBqt9aNH8L+JfP2H4+6jqleUW+JA3IWxe
CfqAUuRpbBl5sF9bu0sw+mvKQdRcb6Wn8NzrkkyOAwcAXs+pR6nwYXxQeDq+9kNwXyDfQvdBnpqO
Cmsd3Hc7P50ZkY8MP2G/jAcWfNl1nBB7hoDcaP2mUCIW+OtG4czDtLoShb7ngikOjy+GDAR13QH6
wpyfVUcyDkdZ3EY3tVu6YMy3EZhVZsxEj4IRpXa4xICcvZoXF6TaX+Q7wuzC5wGXYYF1r14S3eiZ
8ap3VFGapHtA54PXl/G0Mfdl1bDA/zsngVr5eIyqiEGsl4w5V4XJhYDeotCncuFr6C5L9qixrOq2
BWybKGtKSyvdD1wbCKk44ulOCSWqOrrx+IzuhJtHqbE134FAUd3cQW1KquVn2ec4J201/jvB3bM9
tdoa1YbMMZepABD4QxH6WVAuG+bp4SL+owNZJOPd8aIxEiW5plWnkLxxoRpTEjn8id8yu2AHBlX1
WvaPmlGgcq1WlYY1AGlkPQw5oy0r7zDoaMzMw79xeulpModXmg+taCH98lH/pDxvlPOyn81wh5Uk
ns8ZH7CbC714pOiav9agqjybv2z6Jba5YpaMTGA1X+GhMsyt1Wxlbi8t3Iln8FnJd4GG1+errkmB
vrSdJyBZhi/xWoIflJkx9t3P1a/XJ4xaBPRZc0hWJ0n4Ju1N3EWfPjPKYVCYKbLEF+/Ey3KqHz3x
DYtgnKrDD/ahipTo77oORqpAlWlc7wTm+Rdc4fbrGrnKvDHxclnuv32kqLsgreLuRDB5aqSZR5nj
dHsBjqd3YMBvzjq76CG6O9OqVz9Vn7iYboORfqaGblwfi4K01xb+7Qy1ipxrhSW0CL9UwsbMuOkY
Qb6bBkpLPV5uTBKnQnLaa9Dtx0qOP1/cLQIE3LeKJEVOA/HDnzdRA3ew9JTpCozE8h0bMojDFnuD
IeKFGyuyWy4IjqgrqOBCbsoRBqTSiNLHkrmNupYzX18v7I8qA9dAWahurgWEYzV8VCrgyD8wSyUw
uI8uaUHduSTu6ai7VME3nH1ZjTJeAX/LIu5KRsb6iy724waksQdXXNlhss9nokdkETH85NvY+OnF
0Q6FgP+t9DUcjOS8ajZ5u7e+Jl1rTqu7XTE/UuaFnvBSOdZwdfsRBfbvebYnFherBPHHV9CaEv68
IFkhG7JtbZm18CGGMirjsrkOkiandXZS1k69TqrBcN78ibUQoLTXHq0g+tBqoiIw6pQGtXU5wrCe
5pmS/mRtHoXWgqsVXYC6uDNzCz4VbyMMjxsagPAq7LjuYS83Cc7VwpY1kf+3wZYT15v5l7uhZmzn
GWX1R/vbOTi38qhqwiDdLuh8+BMcc1d3nnNy2SKdmV5H8BVBjJpGOQzUoDHOYuFFN8xYemriFZ5U
lnxepI4irJkZ9mMT3iMniBi+E7D1zy509WVpMtlNZUmTg+XzlfjI5uHx8ph0oCYV1WUHdKTwzhh0
KcvPq9y7CNjcI8tK3TS7uylNh/4bnLvna5g85PLTaIYpU/vyOdJpp7rkJN+Ugjf9QxmZokBN2XRm
gfH6LO/lkicA6bCgYCdiyH4Zt5xMBFjblf2ziOMBvUAfV2+7S9+Bt1fs2VOZirpAEK9iq1XMfs7s
jDMm99T1eDyVvV2f3E/CQObpeKy9KzyLFn8FP65y7t3IOBTx5tFul+4q4N11B8eWxsWNqqpnqlMY
cjI9TDOOENKyuPI1S+SItm3KemMJkv+S6B6TBuRjTV/bNdGu6oT9dTt/Tpp5Vu+9ZAaecqYMtXmX
DhwHrwYbtDCcx2/2NPyIy4ZUGuhuCkEUkEhn4K/LiY5H4IsieddkEdvlqwYGaX/UTIs4rpX1Q+uL
/CcOuYd3En92e4CNdZGfYl4KGJwL5vskPaXvqQIPr15FieunmrCS84g4dxVKFgeXEjmKCY15ZcmP
BqyFmMajK4GvALujK26jCfeHEhP9kT0V6W0vZfUEha6v1pX4Z9t0FAAFwtqy5xwggmi3IPl4QsJR
3otJGd8BhoywHsng6vYGOcqRa4aoSkLEWNTkno/p7AV0h0/yTaxpNqG8Crsd3VyCB5sTpSTRLy3j
lgaLtCbOpOzsM7SQf5IlzleaHduzPRUDiziHrPpr7w57v0OmO/Lfet104ZJjIs5JEWoSGMCHvfgQ
KnmVOxs+QhJ1wcbAWfVSoXyslWfFbTRWdeBxw9sYdjox9uSxB+Sr1+21s1NwI1Sm4Nt61fQPYgJa
sTeTdxZT7LiNYnmGYXOxv3E/feCVcrImLTaQWNwYNFSJ4djZ4hRivaZfcpDWv3CWupF9wN2yO/jk
+ZGyXnhP6yD5Mv2scXGH4scM6Km5tHZqqKwjqDGBMktbnLedHkW9RjnO0xV2I4Ce+k8F07/9nbXn
A7MlKsk+6wKlQ286WflomMT7+6tNt6N4Tb4JL+mg4jeaAOi4tVGsDmpGslFo14YAbfQAWhJAqm/R
XKxFGf+SOo6cHXw+d8FUWQkfSmoGFioKrrbfXo46866iuGt0rmAmG9NUO/KviPy3tPycVilHbT9L
ihHlBPZHJMnKJ9ZB4evmIsRcLChtc4/d0puTWn5l5zekHjNjnBqK78mqNPnEmJz27R8oJ1yL0CFq
mq2/M0dLS9nkNPh0/ovea/HSzy7pGaJJwAjofl5esQQphXlBOWJVjbG7uCKrXlyya9o7UrkHZWTh
R35Z0XFsJ9k0kCLEQZre4BFugAP9mnRoUl+SEBHeFsgZHHJGlnh4j/xeiEGZyA3rbzhiWIcLMh5J
H0o0CtkX0sIKaLZkTkJOy/3RSrIECLrS9lJTyxl48c/v+24frCixRQuuUs7Bc8U9lCqOP/YGmJt5
SMqStEi81W+P5livcVzDp1AycrqNBGhIPyXcEG8IeBAqlYQX+jP/ReQhGbfrQm5oMK6Rq8qHsNnI
UiFLiaSzKwzoVukVXZKxbg5SLQtWPR5G9YDINb4nv70F2DJSIyCFYDgAGOPYzQoCrnQwp0y0Diyt
0vH1kChAyuwu1fqlnRCMmsuxd7jwHqCSMacDJ5OI5pchzi3GCF3ifmhpROQ63jmIDZjQR7ZJwSrb
EoQkU4gxHF4udPFNVDZV6ZKRzyzkbCi1Cpqa7ehd0BcAgtsZnKGGVs7UpXn5Ufk/9hzB4IowFbTI
d45vSA0UbeN9uI4q00y65k6BssprRGTtlasDaFJ/Q14ojmTEMzWOgTZ8PZ9xS262Hlfy3LMBTExE
C+2v6C+F7lbxhO2oSTLmLSqwiaA27a/6VRq6i9/HgTmBiEwIrZeQ5FWHMuckIBNS/n1KCQDnDEQx
COG3b/8YJdrALVqa7jO2T59aq4jsISzcfZ34z5V/ffJ4KWC8bRSv1+BbXjQTiUVWnfSTiDAvHJTU
F0Y1OGyYuwVA4Pj2iBzITH5sR2c1lhJ767kYUUh1hyulq7Qa5tM+CzDaZSBmwRVtMM8o5f1lcyGz
0IgOw/p/dJjoqW3h8XirNSlBBH6WP3DI6N6x9oegYXmltx321JZRX2JOu85HDRIRNTS0UicEV/X+
NJDked6lscYJDZX0zpk3bYQTsfIeGguby9kiwXUXBO8dN3hqCNp9LZEOFnXHr/aXtXJNXZYxqbtL
60jMx7rev9hSoxGnx/OUEBkCTbZRgHOk2uGKsLHPRoE2kiViUFuJgOt3EisJaYw7tBYkbIcnRdD0
NquIshiNLlCwWwCyxm4y0Oiq/4WocxM18KaG/olT4Rr8noHGsLUeV9pFSzVXI+a7DkyiLsQby/iS
LEit+mwg5tdoLCiGEg9RUNLQ4daKSXSV3fs6ywWchoH/g1iewXE1+qwedQQz4DIlo+bmts9Jv8cA
Eb9GIK6S8iO/3S8yFMqbB9cA4KUMcYArvcscNS06JcmqREtk+Ao07uD5mGqAflsnQpopQrb9ysWS
xIr5uvwZ+VAs2PP8izeK2QnKQf5UUyI9tIzDh8GF7gXp7HXS3qtBMcLdl0BVGcGZfG/Cvhr2rTfv
Ea2S5ZYXM2GUOYcSO+Cutx6bIDhTTP6N0U6U2a/1Prj0QufM5J6YyxiUkpmvpzcEpO7eaxlHSHbf
ZT3BvaJMQf5P+4XrkP57Cz8use994bh1mj5hQaaCSNQsUiM6oiotje650OmayGq8yg2CG4FCGNGi
R8w4+CRAauYdt0+t3B6lTPuELVGx6w28QT1zLQPEZtGLfuXySPwVCTmn+iRcVyMTeBNKiSo+WAqv
elEZPBUrj4miQi2dPq8H1YHyuE1SRZl2BOotrFSwzAOO9uM7PVDactUKh20za/lDQUnVjy5E7M1c
HMQsBIIiyCaP7x4xyj8xu4Awcle7Q9lhAwyG/0rQv2/c3iHd4+IMNeivXHa29Q05qEaFcN5+I18z
XB5xpd/bjr/IuAuDmMJmqS9vRxuND3nkxPzaFzS3aI/KtN2rpHhixBXqrNRSVm87akM9p4LTqV2f
WlvU4W70XZZ7M5Ug+JKkdJdmUGCFetRPn8Wu3c3cv/+5jyJKjrlRP+YTpPr0nCL8gfm46j67maMc
jKkiyCpU/zpGqH04otvd12eY2ZoKEtRv0nzIJp57MAhW2qpZz1EdJCk1TwI7+IvL7hqxHfmjdRqV
ZpwP5rn6hiTsIA8E8jUnl9ek5MTVc741AoWXFmgS1oexhIzTFiKRiJXz7liqEvyZ8XwLJe1e/dws
1T0EJa/qrXZfucTFR+joZMubu6UThg12nitUv8w9RbqZVC6Dgr9F26l/P+EPRihoJ4BftppZJ48z
EuTudaTE+jV8gW9a2pn4Xv0IPqI6qL+hYX95g/prNyrCYu5ujfraj2tA6gy3Osjy/xdp/0JqSFqC
FdONlRKXi7sjlH4BJ6eZURe4/jInjhHzZZtShrU0qnbgXsB8vxVm1bSrCl+3rpM+r/THW6HPKe6D
NgsWXIvtYKp6Ukam0HRTeTqswZxTm/n2MTKIKTxCshaFiGgRk3WmXI9w/+8avHuJbajWADcTwh3s
+d4D7aE6Kxlhbd8W+5XGVM+k1TvtozI+lL/wUMJUAFWrVhc2eCRKbk5/BZXZzGuJ7C1JTZgQ155T
1aac8bZj/qs84hh9v2sd2jgDyH50MAeFi3gwBCiBXbK+fEnS3V90D9OZBTX/B3hWR+Cs73UPZtNu
46K8js4Mv3Rez1OpFCFJjps140QG7gD7KpENggDSMnkjqUZzqoI4tFbSeCVivFcNX0sSFBzNZUee
EDKlQlFbdngG6FhK9u6VAB7u/n890V7geHqBtyC3Nbrn/PiTsASlsvQ9uC41vExvx0ia3jJ4ustg
IA7r5VUV/65O3S037Tdzp6+OauwLDB/LViZtAJ2kzWCcXdeLm47q/00ZJFpp93awCtnMmgN/FYFf
R33lV/0RWNiv62O31X+QKpId/bC8M8/UMb4rHXMy/Rd1Hn7gHef+aZff+Vx272ZWuElQLtt30cft
4o7/+7IGmAJKFdwoIz5MAM1hr7Z7pfNsOASzoRJLwg+BSccfKxQP6WNXVOF7jl3vp2+9ouzUVBqV
v+yMEf3uZpj3otZnjHTSUO/1GJqgjW7aGDqd5AfDFFm6sFHlZTyw3H3eyEAyLo+A/6B5mzbVTEfh
Z58E4QMvhlX88Xwkg7WpVPrCAKP4GRxCGFTa9MVtraFjcG/9JIdzvg8NatOWq62kA4tX22agZ1mZ
Qg3dCogwIQPlWWbVA7OYAH51zZye2VqNrwoT9wUnXW078DXFcKimUlh3hJC8M2hszgAw2/qVPuHK
VdYVSnq8ZUQvVkvskXtzMuvJ5SxTbyp9drI9BGwqiEg7R5q61vaNBmb8ejHted9ZXF/qMQktZGgd
bH08xtOvAJtNa863/kaHEaFeBjpdRT5ZEcfz7/LfPCgZzfuRndqNFZHYmmSWhY/tKXZdihPxF5l8
E9uv26p/kNyl3ECClF1lRkSjcaRVTCo66c7O++MIIbaxvXD+srFN1HvgwMMOx1Hd4U7Y5YjrX6LT
51MQraJR8BQ64yguW7IQQb8ey/Gprwd2fmqIpHQqqKrdF3Uk/zHrppaMBBDjJNNopsxWqgNQs02u
WbxR4beFXxFT9UKrkaCZTJ1qCX3QhQJhif2Cz5KnBYgjHY3JPsZ17Gnj72bTA69DeKWLjXCTVA16
JPQHKOPaGohqx4drMX7lTfBiR+9diRIU6pbIGmk2RaSfOVxfbaCLaJ5P3vewiCNcsCcLa1MZ8PbB
5qU5xH5lCsHrigKg2IT9HHq/51W0jsmMokNjhtEFQusOIpVWXU+8W0tgvA0Hoyta6OctGTroTpcj
8g3rYudGQiB/+jUQddsbxTtx0hja5bC1hu2S7j7OD/WuGPKAJDn7sm4A4vk95e0fWN42cze+7EFb
UcWnKgnyrLOiObV/e3tzWoOvRVZqBTysNNTGv3V10xaFTJmyXUF1XeD8rbInf7U9fl/eFRwqJQwL
x7uSWxzu93fSzAIDifOcIDIBAEc/Fewg1NkL79ayevNBu8Qx863jGsOZh6ez/E6LuvtbOC75m+Qf
SPdIbnbY1T4V+Dd1DggWJ7jVXAJfxvIPBe3Y3PutouxirOoSpqkBSv0SgX4WfelT0L3GtzTaWk+f
sfQeNY3sPa799ssXZnE2K/FJlKCX5t376TldDmdAazc9ndvpKv+nS6YD5Mzy+pUC0sqtMadAb5Hn
LsIRFlie5MX4imJudncYQlUKgMQsuzAFym0gct0BCUEQYP7+akOZX1jmSZL/j8cjVtgQyvbMC/rS
Ibth9NVpEvzKwhY3PMjdHDuWy25KcNFGIKbSQhUwoOBKTyGBPRA9ffMkJEhaxHHJtceQxJktTlyT
qM6+3xvDCd7U4wvOOpo0uli1Y0jnaY6KmwYiwOfPs93VfczJeOdJM6RfGnzDuFxJmUYEr3KrzZiA
LeoJt7miusiUdnGr4uYPx5o7bvt/b8mMLTAI45bqdSRwvxP3SYineeD10wbSu8vzxbFASI89zmC1
UQb2dctQICOqTw2+NjqQ5Xs/ZdT3BuwNCcFTkFlcc3Oh0YA0Ka1Dafs+7dxtrBqM9tNhhVXbyLNp
E+E/ZiD/vndznIsOSr9XFaUuxQ+kuy5L/GtVjycUw9EoYOE3ZgItG9x6mSJqK8I1/s93jkOhimc4
kspRrpMircGyrZpKcvfg2528RhvKCTm/44XyanbHbdMrRYf9a9IX/xCLqN2gZEp/w8XBPBlqf3SC
JbHDN8MdOeoCEKE3ZGJmQFpTuDrw0j/i6C5QwhgZU4pECIo/8RhjUiCgSXykta4Vo1Jme6tZefZ2
Ctwc4w1+NDmCnzLwz0lPnVvH9teBElSe1Q3sQZR1Fh8+e2zSW5pL5FAeNg5gS+l0i5GH1Ynv0wql
vV0i6oG4vZs6bdDtu3BJ8sFmDrlT4KdbpOR9+YPzq5K0kVFvyfTCaP/B1ZOtp6cRO5EyzpiJ+2aA
UQBVsI7PK/lAVhhN/bU3LGI+LiYYvqbyfJrUsp4kPcTaYS09qUlkkPJCkz/wxjcwCFCFJNWAt00o
prKS12zei+/XgmdV3oRwyjSXjbcciXMoTZqAT2FhS/tk1XFmyKFbd/Z7iF/kRLEYJdY23K4dGexq
JvJKFVXDXgAWf2xmM9s6HpKtyV8XXKn0yKPoZJp2toZuPJW+SJGf7fwoKWt9SL7sL4ofMGD6lcb6
XCb5sjC86lNkEXQyYhTLenWwKt2SZVwhtpVFmFEIZkxQeLiU1fsDSKwV7gU76+LO2GCzi5z+uCr0
u8NgmrhaHIVpZD3hosDmc0g48TJ8vj9k0Dm69x19k+7TxCNHSuCpO3ARdgdGJNOM8XgRYfUAAHFy
eG+uzQIjVoimrIqaOM9Yy4jJ5Td7USFO4GhNkHw6vJkJ+3WjjQJDV+HrZAaE9BaOFCbQSf1V4FC+
k5mMvwq33Tx9cgtX23arL0HjIlFJmMl3nf5P2N4kMstuwdy1aBg02cuXNvFSe9qCkHsmYMHfQHIy
au0lIJqOo6EC+8SdXinbTyQ2QjcTt3nVo4kXZm+K5LmJ4wvBmUynHd4O8VXAW4zeZwC+z6f5opm+
DYlFfhg2SkKDk0q5fNSi3K4BHXryu3+dKFIadC+gfLCZtt3OI3Wdx+bnX4Pf5/VdsjefbSE9Vw0l
o6+eFajQnoUG3+YzAh5YuRA73SN/miqjtGx8HS8a41dQ5Ftc2qFuQ66k/P5jrmjWduTHzRDyQmnw
ESchwQcMSBj+7uh9OGJKTc9BM412tS4PFoahCWo2xkHg4ATUhrnHc+5QNbGj/EoycsmIDAgh80f7
Op8faJp+2fF8T12eE8mpa8Dsb7IucOr1U+i0qSm2NNsIzLsme1iHOImd1GkzIWSQDhLHa0zuG43u
WpP1RjQ7/Ia7tuWNclgAZYrCZzuA5B9o2RxedzChqN5kr1Y/BCWvVCMbb55Y4am1PCzc31zTvTyv
WFlhZDoRQSVuPBSyUyN6LsBqPRWL/k/nZA1OS+QR7y+55A771QiSlkF3p+tfthuhR3JRtr89gC8g
k9VycUD19Z7D7ajDPGeAV7Ueqcfc4M5cke4jGz6lGEkAsibg913sD7fABuD/GQH7nyD6C2NWXjM9
fd9ct9RvJQq9E3V3DXFvkMUnjSDtcjyYDzUp8kCb0L39xZ+EE5/qX45eTh0fdYq0OJezUVZ0ffic
yuFXXMFiMr1maNv1SvsHZfI8lnl5p71XkgvatdE3zzC2MfHRmaC0Ly1RBGMdybl9o1TkE9UQHGCg
Jp9uZ74dLsLpkUYMlpcqbww03aWKBN4yna8/EpBrlG6a4G3+37e0OIfzbGnVXRoEPVSYBBqHzxh8
Y/qmLz21g5vpVvg76puq4t2DHRkvgyzN9YyUqV1UOlDhuhAoNr7lh0YRLwmon35Cx06kCMGOcQi2
UVj35fZsL97HR6w0bpA7g03gMZyEjtDY6cq1Dfhze7PScnsuap1k0ikYa98BFsvphNuHGS7/5pZ+
od6ZPnLN3sY0DwSeIYWWwYcK/HeA1YiBQFq62Ggt2zFG+19UONagGgtCwgic97UhMBz+7isrI7rY
ONgRt/6e8Uroi4KPNOmel5s1AwjgtHI5cBG2b3aUtFB6CeJoTdYYPSfKQM/sIIKAoLq95HzTjmg+
HerRs2K2FSLwYd9NgnmmOVc7LeZtqiL5uy0r/Qk/3lyvD8YDdup9qvVk0Pagzr+UWm1Hb/sSI106
adc5w302Vij6R3WPs3Ct/Du3s1KLDIk7WMu5384pyAww352APa3ZTE6Vb7cxknDGBIAMo5FOBx/9
tlBYFTalqjlMQ5o0SYdm0vnQ5OL8DucYuBeWlcdFOA53T1f0WjNIleaWRjnUeXz9qb2wrFUmEeUV
VEtf3q93d//7oqRYR6Zqis/w2vmYRrxMKLa9MhVpHzAxYQipqOucZo0dQidC+oHyAYDLDtaxuNgm
Z8SpxkBHbxYV5OGXkY0c39YOZEAQ1m+mmycqHGG9xWJAGOhatgHbs/wU4b435uSlrz8Wp4X6s9KN
znU/rzw0G/xEtjvOsQHZEAzdOpM+oK3p+fhTGtkOdE0M+WjccUesVwRl4y8F1sjaOb8yFEGMFJRu
QAW9JWh/UcsFOIzn/WQQKqxZLH1VR6mDRvFCqQ5Kyg1gE6vzaLI/ZOnnpXd/9jaHKPLNQwmiMKYJ
Q81u26wtCgsN3t8AtebUawNiG8HBi+/GzHeUiT4t+w5FM5TPRMKi1iACYJwwnJnXVFqnd3pH8+CG
9pSLYFvb2lYxPTDw834r4iOlka/bHlZUmAilYDRy6pJMRdBc+x0GpI0KDUjn7BGpVaxRHcgUYKnS
ijZ00DBsEP46AO6DAfaG26V1rRugIQCOBJZaXQiykFkwHn0FCavUu5HwSMu9RPo9cW31GUy0dc8d
ozGMPXnQ7bRLViEE42S99QkLjCD+YkrE2azHi/1PhksQjr9XsWrnotYaFevWUC0IGZs6qjwJOtvh
2p4nfmm2X+hvjbj2U+fPEjrZChkElznLQTSYaEnvCF/eiUzTZONnHdKRflUT1T2FECIWZMoQPiF4
35Wj/ywcy5ZWLXStbsE885vM/ZLJcI4WZxaW05CXUM8vtCDYCZqpyzdINY8BZ//vjYA7CfrBHqW0
223+P7GJkkk+uWE3smZ1QT3o1KIZfUBdfAFYWp+u3TrXV0OnJLrDDqK9i1zSm2a44irw/228RX8Z
Oyqcgq1G0XH7tsd3FyHn4V/ZTLiGNPcznm3ot0jpA+zaOKcMZstRAjZ95RllUWAYScZzqtQerr/e
wUs6Lk3EVEMAGtp1/STvf0ssaadYZaNNU14bH5rxju/Mf2FJjWuMWFbBBeIgsD5ayGadyERamB/+
jqa1QRyQsbzEfmIUjypOLS1BgcH4K3va2AxvOI/b0oUn+NCE7MK8wEFzOSvDKLGuTBO6xNgd6hc7
GQbEg2mkfxpB8WtRGzUcKqp+mJgfiQpc3exBGAD1KkL7syPnrN5Gm37vtpitTTVEV/XNBqnyZj/W
z6bGVnXLiTcDwnkKU7YZSnFFc/cFbZmBtmJrvl0xTGmoJTgWohRvqnpFSgUtg34tYgmLTfrgFm66
BgM0aC/5cNQ0GzpzS3UgvjSuTpoX20YfBUnwbDAeyM0Dp45ikxTpeMOD3CtaALdIhOJm9lI6QroX
h33hqY2wqxOztBoLwDGr1hwzEhMmJDjulhWpUSadCR6N83CCxTv3c8xqvp4hoiTradbHbw2CAC70
VGUT561dRVIyd0IPrQL8DE7X+Tvs5CQRgD34aDmnTiFKAEPipHpST58Md/BFU9/gHLAB1ziV+btZ
JXwz+05IKLtXnXaNKAymt4zPrY1c0WbogVgrB9979+/qRzacAhaLcCBtFvtM3jPDLLf6Jdn340tK
XrFNnjqm+uUTJAinulY9RU+GbqB0j8j49wm9wCax4HIoHngGlapU6EG7+iWyfEy+mmRHiOw5axgx
rEYzrbikVNSB2VEUmByhgkjkyeUIGH5JKmYG5yb7FOx+98Hh1QBCseG48na9IFvbEcQV9hnjYZyU
ArL3K2pKuw+3XwY7+DQ0G505H4RLeAcgA4jN7pCvkM508N8jSufgJsABcKm75naBYZGReSVxcFwr
wJXQfSAqjeSiBRlYLWTMpiiQ7W58BraFVpHaXWeww9o8bvuMMdoMU9GnSv3u3Cmsb0Ke1mAGMk/I
hgWMvhgYEDx2sKJGmTwy0A7Q+w4Dl7WXsGFy0G3FNNcXD12RJQZvTfPsRU5qC0Eox/sIvcBIT88j
i9Or0O4PrTMX6IRQagebeSue+BEoA8RLsX1Df9ox618V5HBr1SR08RDpOOHvgCKo85EK83nVyPKp
lzvFIrQfFlQjDaJyJNIexHE0zR10Er5ilVPoHnRmr+AkNZ+1sAKgziIjzkwsQQDKNcMTU8HxmeNO
nhi4evciWzfRFmh2Y0Pg3+kO0OQZvEYFpac4undP9eC1C8olETICScIUkVjlCTXHwUAJ6Ze3gPHh
tMYG7PzAHNAisO8bkUiAZiPwIH29Vf72YvFisQqZJZtF2ceVsaBu+joPRpCvh41Y47hOx4lylbgr
2c8zxe2IZZ4sBlnL+aCx48/API48XtuDlbdLY6GODryMsnu6IajT+ga6g2k9AtaNrfHXefCglTsB
dQ4lNR7QnAhzqeWde4vtwy1Xq7l9dmNxzY+DA4Sok+D0xTI+8X1D2B7/ZSQmQYUjwkRyj2xof/RG
/DNZ6VqZjseLcCkf/EicGUiHJdo1hGWQUEMM2E5NQKDvuU81dfC4ah37HFes253zSa18eD0PZXHm
7wwdIbsKyP+k24yfDO6NA0YRRnX6pqi3O/8doDbBApzAPhX5knCCf6zza+64I3Cv3tOfSY1qKL9y
umW7TnAT5mWLI6kLWxFhwzYKx1EgxUDEa3kOYFhnXqXc+SnCvRGuav4SJtU9LOTsuNdy8xpj9ZBi
aIh9S6QT2FDl97xjQbzuh36Jqhv2NMLvzo2pcjPpRz/cnR2seD1qOu18txspZ/oncMY/bTu2wezq
IXyRQyD3zfTdfP9sYfRZ5VF1TgRbOzAF9+E7Da/JZ9UCK2g1QoNxzbrgA1EjD4n9ISUJDxI6MoHg
DZeLf5VjZ8xlwXTHhCdxmQ/ieAEXl1bIJc1tRa+G4o6vfjqqLoeL3/SG5AkHuOnCKWsiq05nApoO
wrYylpi9TDAsLexiP+m0HNePH/dciZI5C0BhFX04moyIXmt8z9nsHwmOkbK18RLoWuOzw09xDyrX
y1t98xBfVMLshhrdV40CP5Mo39lHW0UXWgnHjDqj80YINDHCDVP+G7V88D158fuy3+9HuwlJ5ODe
0TpjlWbVTtnpMnHIL0iYJFKOnQidSZok2kFbkwnkfWFmO7GyrVH9jeezM5sVQgymNAmFppQBmVIA
5JqYGBHgGwgaho8eviZ2Rdk0x+hp1clM42sypN7DYsnSC09aoenesQ4peM61bN7BweZIbgm7TnFb
oXXSP5r5mgUT/ted5UwqFNOxdXOLkulHWJZEHYuCegDbBtuikV8cp1BgH7wcuITdLd1fg9tDQboP
MyTncsk65JMVFxySzIRFtJ5fdcP330Gb6shSGFxFmPy1O7SwxRpcrmdMQ0EsbOduO1kFLJEOPJxw
wdbWi0UNbU3DZ4U8rRCOk3tA1jgFAnv1oS+y4vpCRyu6u6vW8r97jvaesCSrZjT9XcZONntobZ5x
OmON7Q8dDGwTcgaif6uVYK/h3YxlUDsF3wDRcYasLFohgk6yVy26Jtvse8+CPZIKtgzQV3cdDmjq
q918ugmlONkNTMjEqbqfliay1DLJdJn9iuOKDdkPP5aN2x96fGvySMbRm9pe5/Xkk/PgJ1hC1FKs
hDZVT1LFfNI+6QL1QA5fQeYRAckVcD5CU6YW6aG/QnEcet11ceUqLzcFe/c71+FeYL+FLrz5IZ1O
+KJqj7isSH16A3+RVFbs0wVN4KoGf9UrP+TDRSU4/DRptpyHp4+n4EE6ikaa8ag8Ft1XDbVVoDs8
jZAf04q1/I4H+5TMTNSfzIDIDGHynzZHL+EBMH372j7mpZOKUCkYkSRj+lotkdwVLW3XZqzig+aP
2WZeZyHYr4Ql9aDiIIx12pYbLhf0ID45UeHPflP1fk5eCU3DwyKlJyzHg9yzFh8CXqMt+ASR+rYH
rptgqqF82BYqT4Lt+EI7pNTKlXWEGhWNpjrDPWEriGjiobNrb6CfA/0DnuHUgbMM5ByRZT0Ef28d
NM2x+3eapqMSt0XL0nkYaUJAecyb5c3/oeR2O8Y54r9xPEpZoZ49WiuOy7oq/vHdnAa+r/om+oO9
rOk9Cgy9K0flmdQ3edz86g+bS/5Eo54Cfc0ijJKdQOcaQn6/uqv+a8foU7QqXA2tvVtROrJVFTdG
CiXVJs24F6NygmEnbqosU8ThbVtHEIzlthg9q6iosw5HMP61g6GOokUNVmLwqQ6eeccP7PE/dgeI
K6dOAP45M78VqtI/S5ZR/lILu8j1Yt82CrO6P07vBKDNCXtxZYd07y7+iUUyvoodLi6mCAlI4s5+
HoRZoDo86zRO/Fl6aYWj8uvkdhZ1F1G9jqeYVz/BXW8YMPVGAn8uJ16MirsMz4A6Cy5XyG9P9Lwe
Ltbay8De2V5jf1h5rtqagCiEkc50NxokViT7KlXALpFhjOPCv2gS2uZA5UCWhKhvfEyYaZogfodA
h7MPEFwQxjXADSmYVFTLWoFRyA/QXYpq9XBsDn696U8X+9F0Qls5LkfAZKdnZFGM724Uv17KFxjh
5XMO/rV7px3jUQAmwTTgrI+fLl8+37sJZSYKy4XiRwhfiZz+96NT/c/zfsu6GHiVmlkeqXKgrnLD
rysGAMXxVOSxX5+5AIu70SKelR3WxstWE77rJM1aYUCqa3nURYeYVPr8Up4TyqsN8gUN8uYy1puu
tvlStCG4YSR/WtWRTppPsWmu0IQADNJKas8IS9WkKNDMW2IYmUhYEsZ2PVh8V6qTvtvWSyzMNiOk
yswRvPituBGKUs9QaypqvvWUaPhQy15uAk3gtIiCQtgrYMzP0ZhpkojE6rgV7RXZfFU3IrmEdRe9
mL9lr704G0m5IlxnWd1v8eJ4Yqr65GaVxAtSAyQVoVvelYqXdovK1KWE4sT4okgfYUuOQimJdZqs
V7IHKkfJ73AFb3wv96/H6soYpj5nLvbghFH2JCSr+YDtzJWgzg2QaM75R0QBf5ToffhRloNesbGm
S1/mXqGvvZi4dU02FgxGtIG3AWDF09PJyhPwqYQR8c43doUZ72jYKwXX+VJONIX5Ld20cw3g1QHl
bIO/v07P6mfMiTnG8pJqVJ/usUUqAmunq18AsWTc3Y3WrjfXYvjhJ5hUMbJAnPxrH6NkaTT4ANUH
qniMd11CWFmcDK2LqeLPebPfIuH/9pHhrYREAM8ulllC8w3+fyqq610CMS34vqeWWKhZ1xsgmbAN
dTO1SIn6imB2afVp+jp3+dcBp7uFjvEjz43y4J4qhIz7ZBqXPvrCfrPMuozFdJC1tekm1SfWIRvR
GmX+ijdxLo7dtbP0GiGL1Y2cjmetH0/3qVHaVVoJ9mt0wLLlKt7AV8lOXpessd/aMcYBaKxtPadO
WQk6nxIYnW4qAVavqs8YZ5J+a1vfgCNHWEZPbWj1ccAN103p8ZzjG6qLeCYvMNHtY3l6GvBSvMpp
o5JBr3RrArH/T7qsFVBRO7DYb7orxXPBVtgUUIB1Kr0QSnz/UZho7iqaErlsRIoBuM5aO0/CxO1M
vcINZVVyFa/uXzAf/BLSCSEUDBg/HUi+Ulo3Rf42WUnGtCZwGjXvjqu1ohXxv1O1HXblBDOd4V8I
mCGE4LHl6GNmOQJMDqlr+rAgC7YeRWDHsFy8c8BvQ2TUcH4iXi6XVTYLUB36jo1pxdnPejszrE0y
ZcN5Zxcfw7BYytD+QnMXgXKXD9bepkYMleJJQNhl6Hyh74GubaciINbF7ApOp7H0Css1iIov39xc
pinwuixc7GziyS0aMq0ceOphTqog+WYCN6a8c9ouhuFPLfZCymO3EAPxW8g8Tt/vShyuVulTdNUe
96TgtHcxo0/N64HDrwqswUfzNs829HRhmhb/JfQzyu48cHpcUGftSqzfVqk3USQJo4mbfNoAkzGE
nsgJqHoHGJoTWGfAXS7Hezh4NtbB+iu7t23Cn0aUmuSPsqsgg1uJV+tlguiV6w1aqsA+ZOsdcEUp
7hLfPRlmU1DylWek7djfeAm4hOJPcudZukXC6hIsvdrw2r5VlFN9o3teX/qJk6qyb9TKbfVkSJIT
vSLAb6QWcJzksArtLju1fsSGIoz86QYfCTkU1xeAvqgotUx28Xw8r9eJ3HQZW5+AnbDMVuUEmauU
o+3uhTNRRCmxB4BC4YaTyOjV8IHRLm43LHgq41D/ch6PrV17vdMqp4PZYBA7zEkr94Vpc2RWy8Bh
xjnP10fWANEZC47gXQ1MdmdIy5hWIh0PMXBMz50fSN6kItZ36qpqwRA3JqAbAkY0/DLmfWpBjlLv
64GVP2bf+SKwfpE+u4CaUa02yUSLz9m3WD4zN1q2mGpTaesTY9vV9xLxnOUe2G+OWumKk6x8vwN6
QK223bxje0B89N9tFzOJz08Dzq8cL/akqWMH6/nuwU2rgQPkAF32Rntem1WdKosyUrGRLw2S8TU+
dXm60p/zyPqD3Dc/7acYv2bPqYte0lAbK6Qp6kAhMz4X5mlx1u1csm6vxD+bvG+AhgPPIFmxBYAX
lTDV7a/OBa9MPWjBHresFC7WBFWb3hmN3VVmTNJnI/SAu/BXJuh2DtsoWJyDyuK+JBJRi04UPloK
47slSjwF5aTCZcSjdwMTUYlXjPqbNanr8XKymhp/ZhsbdUpyyf/lA/BxmhyU0FaUq/Zjm5m8QixY
L+dr9oyloTOxEDMKbDDyx/OAKvz38R7SccGXgA+wz5fAIDjHo/+iS1/eA9UlbLYzgYdIY0XXeHn7
tkFy7tocE+z5rvO3VRM0hYvvi64BlGCU0PW2o1oYw2XCyzgZDcs0NiY+zUdlGHpzd/VuI97aYzLM
G2L+KlDXh90tdxZQXGv/C95o7AEkiEbEK9SEsSOrLI7OrmT+TTeWq1ePu4Q5JuXAAbQow2cHxGzq
HS2sTGZsNBsAy1cWtfSpveVAhl33MvF4LZhxUBXqVq06Xgq5Ym2GEDW80U2Q4ydT6L+bR6sT7JSX
aD5qoUOnDeon0ilSnWdZBfi9lkFKuqYyww80L9F8BzW9ZI+YJlw9VqVKa1gLmiz+SBwT1xUhUo2t
HHDc0gO9WrsnfVSZF30Kyt6vzhyU/J1xhTiuyc19s05rkKa5Jsa5CkFedQYdifBvw+vWzWaTM1WM
eGLddG/q238S8ajCzJSqyvQGnOo/ImjYBa7XgRabfax9MJypDgcabB60v/xN51kgHc/NMd00dLCm
rDT39mlNwoBnq4AAloUI0jnP/kQH8BtdlDYvqik91j2FB4KgudU2rrFbI+ILZfmrUdEr4tP9sOxp
dp71VCXunRvhOGi3nbdr8qVtnBJ0oRGHYOeLlYZqk24WOQxfIszt917XEEE9uAiv3h/7Zgf5yauB
KiAt++FFD47PIwk2mFqIfjMG3TPuPWR6WLjmMA9o9xiFGKMsslBQWvhve+ex3mJT+3d4WvedtjBT
K4wnoJymb3tFSUkuFZsj/pV1xEqrAW6aOy2BPrhS4EFDOTCk/zC3g7vo5/q9AbzhxtJevGwn75Fz
zR8T2cqqBoccEjvkSIK0/8OIkg/iT6mVLpjvTz0jaYnwkKWy1qbk2vDo1flAz4BWTDGUV8IzHqlu
BDJXEwMLpWaShZgLjoQDyYcLx0/uxlp03YGYZeHj0+3r0WzdHtHfaSs5Kz5KFyDdPtTqwMdmbV6G
9G1rvFhKNtcYEdeLrpVZ+ni4AirsvEjzvUGJ8HI5149/qe8T/o45IaPIMYz4Hdg9WaPw66Lhr82D
GoaoNez53Z4vtigRSv81hlnsyOSPPYffJd5nF16Bf9gHXZUxJedl2G0rX80kr7PLoxhpIKck4Fop
8KeYibL4dwKbOK2ZfrwhUJiltanG9vKnZAUKBflhOmRC4xmQiHLCW5cBynJLBNhyNdtzPGGEMnA6
99yaKhuDjRZtWmPe3HDnI3QTY6xL1cxlhg728/p2T3wwo1k1vbBAXg1UGCrUD+Wp5DjaEwYJVZTR
P/HKBk2io31jFrH/QT7eUG1QW6N/6VhJPS0U+lUywLEGoQLdmyFT27VTFNN4tNCooYPqYBKrH5rB
4XdH6vrTyjawZowRIZr5Amad3AogKq15pEIwJf0dgyJeR5+MPis0a1WVD+mTb1NMZbUTGl5R9QI4
e7ncAwhqLgMipFn6Pam1D4o0CJukj+XqlNR3HpLs88WTox5DbOGZsSoonL6EvDzudg7eazpeJwHJ
HihhkDaCEagVM04JWpMmzifnZ0CQWO1tYRAl4VVUQlKc2boZW6ZtKnz+p6jyL925xgqgddHASowU
IgEOai2VWm10yLOlzQIIkn08BayMCaIo7w6sFa3ycI4RNve5ad12ftOh6LHwzNDD0zjsaT3hiLUf
GU3DxIQgrYl97euPvDsfDtMkVxW/Yqs+o0ZH+J2wxjUy+4XA8HyJxAazswl+BFKx9zWW42HojPyF
sgr7+pxDnGR7SQhfv5/KY0FYTsEp72c9hO6a5dH8Q7NxIrM+zcfPj9Cswpx8GCCJ+o/TW3zN5A/e
nvLQVfvKXwMAR8DzGLN/xX2JFxervqbsUbxcJLdYOoO8YF25PUYy8kZk8y52wIfqSNzArFHyy5pI
9sTdkGa3fQ+V/CbssZTz2ksBNuTx+SYn+P++HZv6iT8VG8PhRynfx8CYwVcuvt6fwc2xI231zRWV
QUz+QLDmvtFaOw4V4t94u8TfzE/XfMJHkWDJSZrhsFrID5SCFbPcvo3q34Kx6uF47xEKKQ5YTcXs
wsf2jiseHjFkFZl5maxPWOQKWkRzZgb+2xzOW4V8M4lbCdFxIZvR50oYkGfY3ChCTCWlIbKkt/Fy
mzn81myX1WSehGD/L/2S/bHGH37dkVr7bOW5eogwpPMnjjDHCLnWA1St453fzMp9J7uNsdTjvLmR
aNYYq+b9mq/prykMJg3KjJb+nflr1KPModTX3Kt6xTgd04DBzHm/wi3T6BZDjckxDCmK0iQ//zLz
mRao5Y21Q1NkK5r0bGSF38EFbByRWQBNCwd9sUerqe+RB3672xOtcoiZGfxFsYaVU/54ypp1VjE4
cL/R2Yj6Jv/Ibo8c3DskaITdfx0dHFYPJIp7aXWmuhPjx+xETgJpReVdo8L9DWIMFGpj6/KWH+ZX
wt8ybevUkdbQx7BOSkQf5KL7uxo1/twoQexXjuiz1VwR6Vg36bQiL4Ee8Q6nVRL8eDLwVd0Q/5Z7
JmgPFx/nQoKRl3oY9blTK0aJbayQM8g9Kb6VcQYvOTexbmK6OKIj2LhTek2kEWE4EkuPS43h3Wsd
Ht2xrvXIHVC2iFf0ukEt0pp5gdST1oNk1Ba56wAW2NpwibA1MXuDwCfBnQcQ7z4Jw86qwNz1qQ4D
NrP+Wu+z8v8Z3oV+coaATsjEP8kkPXWZ0OTSQdsLmsLdfGLAx0VCc4bsYJLguER/l4EnR3+vfutF
DiuhZ3piTCHNr6KPo6T+B9/oEd/MtLc78PRxCLTYmDrVjnFQxbl+CZcn3xX0F5rcbVXU4bY0DpUn
f8qwA3FtkrDZzyD073bywqhjSiuQoKNxj2QnAvWCxh0HnAVUCRKTjeNTViTXAoqRIbzsWrRt0p8B
zMJdxD0Z2LawIcptg7GbxQdQTroCj2Hy9uM9hYBk6wGrewXKpiHUUxlTpuY3mMEj7b61q+N92WT3
WoQ6eL0ookcY/HoKeGbmqBGn/5pPHLvSRT4xe8/qA30NH5DepxeqImhFYH+812CXI58gbsUwhqio
j/wFon+0d7omRMuT62lKgWylvgW3fsdskeUp63as0jjg+9AQVIrwrYcbxXiN2ng/KBGJbcmDGWxw
Sa5ZtW0x+DrqZEAI2SxKOQ0bmKFD+wyRRn9q9ZiBfOcrFkW6Ye1hb9fUyAjxR0xjGrXmmsXdDaW1
PLX9O3CJ8Z5gvF/vri41jzKSTdxV+Vvba/Nl3jOncGxMatCbYYb8VzaJ/buKccDiQaKGFmL+yBoX
S/s74+42mszFdhKlbj0xurTSLWUWk69ufDAzVwTa7eMgak3RlB9YWmf85hCUV5W19yFfcRSPSZ/a
Ce9N2xVhOCBcSdmof1IJrkslLF37cGgC1gkvGrVFxtyQkqgi0UscapDPkKHcerosuV9IKvx35Gsc
uuDiIFW3S4RSsAZJJPBRRHaem51JXEzcOZ+dglT+pZvzk0pu0WT2D1ZsWf1KMzsccDyp5MGvFAXw
blG0C3r4HCBtxBI1b/ycpadJRsVO+NBrj4Go+sEKJruDQMKzM1rjpyrDmqTMnqedryceeT7xODmc
cekhtYNdsN6XFJcWT8YcUO6F/9nQSt+60qLcNhx22aj2mjTl4WfhrEGLNpGRmy6Gjme23umkRyZy
A7oY7znSYXPvoCRGZC55WwN01dYW+YBJ0fBP1K8h41GQr2sY1XtgLIFTDK88rLVwI3HkYcLe4GR6
x4Z588ye4G/hvHKjjjrDPE7x0nFjt/6Zzhc2dMKe3YQZEJWZJmZhemGPKObOpCMHFEOe9DrQrHdD
vcTHV6Yei+OSC7VFZKovkkA1MdtEZMm1HNmFST6cDqWiLkT54ZVU53h1Jiidz6NgOkNy2gQ88FGN
ZV26am3wyKZuyootm8vPSwwbdOTJywxQm+KdKhElqxa26gLI5BcYk5wiGPg01tl5mH6WeR66ZE5y
kQ28TNXfZHD68vbhZG3BY6XNPRjK67yH+YB8acw041USnal1UVhwYfzZo+8AJdXC7tuwQFGv7d9e
rr03CZpmgtTufK0s3vRk4Z1PBTFn19hVAiuwIqnzyR8xuNalqKDpJw+XwGiyih8iFWwBoM7xt9x0
pq920fIMBkAG1U5V9gm2PmWaaislMreVtuAJs/fCrVqHcnhVBRbHbQVIgR2xV7nDvFyjSXL8K/CR
e0j6C1TtmAFtP2ksCjpcLb/e6TEYCrBTix2+F6XOhzlQaIRvxefCRV7/79ENsk3rb4Yc/0IF84na
ou/RjWLF6dOsSJSXHoCfj4OzzfmstPRyJzWpafvHHLWIE9R1iVl/U7oph8OLc4UpFuow6aUZ8r8N
ePyNNfgthO/Pje8FnGz+Dt/UbzcX4vwRPCm5bkCJBgYsvQ9/fnL9zZ9Bslv2Jt/2xZMgaiWAfPlO
kYJ7qygZJznhlHAvUEgVJi5SwixrnQdoZovhFdtV4dZCOZ1AFSOUY8GG0Ab6VhT7IvR0dH3+k5tF
uZaIkiy5JAxvAUQHvECyQdmNpy84O3I65a0AUrnXn00gE8nrV92dP5jlWAfw0ZmsFLnQJIloD4jz
rcGPWMAtQv9JIeo5oerw32WiMqYbJh8LS8VPUDFRMmHqU8rflLzVNKOzufs1IUga10J6QKpNGWhF
1SZyXtTl6UUN2r0qOBte2LcITChKGn4aEM9ptxV3Gj2tCO2QJL0nlz6qeR2oQkNoYoO1/PUZowbP
UvO0ntLMGdJ+3OA9RhGbmAzJ7LKXu7cQiBbE8UOJ7y8KY3nYG7WU9oM+CzByTTh+bf0W+mTxL6Cn
uHIVu0V+RorLSdM7d58Mdy7X7yVmlGz6MHqr1Fs3YCuBIm7weBTjjC/8fi6H8ZPVstrf21U6NYy3
oIVyQcGmFKQ5LhOq7FQ5VLK0rjGj2MRt8KFxktsWl6Wh9LrxWWpocTSJiJSV6CESmeZz0JRG28H+
kOFqyJKF37T/SvbNuGJ5pGP5k6bKgks/hQEsm7D9tzzA1RqoMk/nRSFPlP9r4lokAszWrboWNhRA
IyszwEW7ZR8aJs4Y/2ONdf59OgWTcXZz1z90JpBetoRrEqZohlFuog9LO04G4yV4ft1LwA3QOVFz
4cv5Wn8bMEnM1uM299EGGem6X6t7O5I7WBa2OQc2Ng2ImNh5BYEiaJ3XJ4QMQDvk63BQWw0Mgub+
vI+STZJXKCjrRKNzibTq94FifvrkOiWpm/0li2iQt5kfkYm9r28g1j0RbMCWdfwiDcTS/g8+EGaB
+j5hmAR+OF8ijgFk8CUB0F9EjM2+unHJPVq5N7mbx+0pW5l1qp/mG6qJeSY6jJYjzZhiA6xfphoN
GTbxJMGSI9WVldcofcKR+Inajx1fbVJAbV/13c6FXYtmydjIJnON/beOZF6w5LphSIQNPfEL/eo4
fhLN0wWR0femymbCT3WEjzyeCNP1fHTzWJcQIVZb0ux9KBZmcGEj4AG4fGA2j5fWEKVjhAQ3nYID
Mbv1HATAYDVtFgwC6u0MfZUY8nu5tf0O6WNd8SJtCiVnRL7ZXYlcIFEDahujV1UMok60tb7ysD4d
Pd1fSYQXMrPyYfKCK0zexzn4qAtKqQc9EO2ub3wsX4J7XQAtxHYMb7ZnJI8KNCu0GjDvvUPvHpBQ
yYtbDZi6j/qJ/hDyUYbUB/lA6vHJGzv/C3cHShs8TnvRkHO7A6ZY/XZmns7Iu1gNou5UMv9uhSIb
IMVhnBaXwzmoB78j8A0V8qu/PFGPd9+MdzPc4uvkfB1Qtd1j1xHGd//cZdOiSM6XYKRea6Z+pSRQ
CP5Wev/zUKJNit5kn7iV7u+NiDrYRXyRqA38oRY0jmY8s/2561To6rpH14qBW/LnZkiTMIBtbyMM
jhONNwzxcyNBG/HZnuOOnAIJsi+5W6cTYXqVsq71heIUaeILAHXbefHzf8o2gAvAld1m/oppKc1o
Sh0kUE7seGkWblo2JOxtAyOZ2j4Tkb36BBbDHK1+7OqzOinYRPiYsX0E6XdqjG2xLqJFHkdmlkx5
c2bBRMSBluRDa+jy4cRbSl90w9tsYzaAkQtqvk8X9cmpsqXxh5jEjSx4i+V81Ii6kp4hV7F+Isl7
DTHHB0u+OKmhOISsJNo8gus+WNHyjgPhLKcn0X6PIa8VYgu2daQEBb7nMaeBDWEDmE8hGB/Bg0tX
1lleuca+cA+39xp88/RGGAGOrPSuk/AtjukCeYAaLRuNzOZuFfZYJYLwaGH9d+0gvziIYZxFinGB
GF6ivD+Mf96WRwC9nFpe2wJf2ZihzkKELyKK/BM+86rEI0OsRUTn6dO9n+6lKJ6sI3onwzej7Eqf
308329rm/0niOLyULYv6VexFT06kTZlcWy1DKGbGas72NZCtw6imMvpyU6rQElhHeUFRNR1M6P+A
3YKbhgaGR4sMRe08uYDVetMDi8H7sMGvVfDmvU9daT2OAx48AbN732kU5xY0OJVbhTl2a2lGMkFu
qjPeY+s8tk9vVydMGkOfRjETeppUtViopM04IjDqKeefFTQNZFY7UxinnKQNzeL2BIwH+uF4a2HT
ugmMdPOT/KtrDG38KNr9YIEZDO/rVk+plptIOm+WqjyVBH05g93HapnuRL3R5YygBu+Zsv1HizOQ
asBifhklAHzmbhfqiXKULN35Fw4lrHs66Gd8i6kMWSbzzN7b7mt0gXAZqqllsnSQ+rFR9aytK1LG
QKYMkrqWVZKBCr2c3y1HsIuaP3qtYPWy7Igfn95bCP2L9Q6lC5vu/GM9lri7rrB8bw+YX9jXh4kp
Ryaf1Ru8qe0Cl8iSjN92BMo88EJqZczHjE3lYiq7/NyjamSJ9gN8TSZmONecJy9a0m1XwuOrOaiG
dEoJeUUXeCRyz+RJN1sBT+Wl43KBbdk2njBAP6tb3x/q/1fW/lkN4m2rJ1Tu6z1wVq9zv4g694j/
wJ13GaTK3mrZAVle/8CXOIZDuIM8TZjY+M4pTX/4n+rXYqfCYuWhWhTO+NG1yRHvUmWEDxo4X/ga
MBaLINZL71WzoTIqlZKsO1Z++cJDQBRDI2jT/k60yd0K1M0t5rgNPMCi8NyyTIIEx71Olc7spksu
JjgbbJd8lfiolZVTSW4yxxB3B+893+c7OHAGA4mZq1JNUflqMViGF5aUac1QcBqea+VyUpx59GEp
Wmx5OrexVxk7d0BstE391vBBjaw/R6p6w9s0Z1caNslpwx5WyBuJL9wcjcm1s59BuF46w57xtWtc
PjiXgOokFQk6vw7gxJKcKUxJqHZ4nGsZd7+wd57R85yyECrxoIRNNfFHZ7taQ14unFeu8J90dt/j
QfEgYC3dWwFWn4XGt7mhjQxYMAjaZAn36nhI2D4TjgPZxPDz8mWd26Xl4hkrUthuav9CqOAN09EA
jMNYb9cc4429Qf5r8Zhxn6P/2L2RuASO9Jxz8xp5/FsgeLhUuXnU5/CyVvE095yPFuQqJcAUUZuL
GZoKSgRUVoyi2qqL/C428t6uPM9a6FeYdRSEh/VW+6OpusNLh5yWOPTvMIP5K9OGQw1jtkcV8azs
EG2pNhlihmQ6OlSOplTwqdUYkK/G9hTudv2bJKJCB6mfyPStOgFS2e9OCJHIIj6o+8Njq5lQkzdr
UL50+0Fskp6vUO2O+1tyQbk5zkngocTaTCGOCUKOhB21BX7xFK3+rCsz/uRNJSYYhYulXPs5i+Si
xr1Kz8kqpG3C8uhHhgssJcr1g1NyBD0H1j0NVLMvO374xSgioBfNPhborIY8QwgUIbgFd/yaxSOK
6DrY7Vi0MM/R4IsUG3da01VYs9G+5EqeyjcKnVSdfoyTf7GfnsjE0IeFV4Mp+oPcCxUYolcnYTBY
KoOY3olKF6WSpweTLVbvDste3ZEpehxE3BLVLeCSaDx/+XWL5Mb+P+V7PdPJu3BK/A+kdqKFyrSH
H2klCJI/o1vQEpICZmHLDtRQdZuROBVD+A5KXqEiYy0rtN7ou5Oroi7JLrDdQnVhXSFsz+6PVUw3
3GvFVAbkg1/8XkVWqUofsEastIhT2i78HMt2fWePaegzBUh37ds7ijHmpkQXqAecG1H8Ft1F0BZR
hw+bvuINpxZSXdWUJKK3O2Si9lrdHEmPjjVHoA6XEd4pHYybOUgUJ8n3N265s9W8PVjzR9e0DqeT
JmWR9+QOABPGfz6/Em8oGsHJSEWdW9mBxr4F0F5m6dvWZlsUWSEzPNn29hW7oozw2jTpTzoqGsjh
FVFQcVG1GmTn9KQrKjBupi3IzDWWkW1TQEhNGzNHMLWKDXW+gnjmMu3HjB5bJ67Nu5MdUqi/xr1N
2A0TYkdVsZtLoRcD7GUtjWf+z28ek4fGRgefKE0eG6atETHeBv/nWiCATAv6HqcY+UnYFfN3MXW0
7tWicfNkogejvNhL5z2MkpyrBMOEGQO3Tmy5o96NDnxdnCPNe7/T26WqFoIsYJY5jSLxDtjJZOkM
CYbyaClHg1s6yZKuitTcCUuFkAm8mqD/N9Pw2LzqcxUk83aj7rEIn9cRikn3BQihgQzyLsbQoOFE
8LcvjpKA3MxnebXwalj7QLcu/u82xVVAn2qqrqLu+WKAkVr1TIldmUEEVvq8FPcTcKwWzNs7LePe
nEp1bKLqerAdb9tTuB9Eu58p2SnmVDyjYkIvU+urWQDDRBHIdYVVZ1Kyg7eTgqsjhN2WZAYzRO2w
L/bb9MpMex1kaVQUTOGhsX/Hbu+jnPKba7U0qs7ldqeumcyf7D6sh2BnkqK7AHyJ/ZzjK8QO4eX8
O//Q17FLe7hwezFrBGM8hzDM2F00zHHU7CaowyEx3cp4Aq5kV3aYCX9w1sk32B5oAZKs7gvtP09q
M6n3/2TEJPxqY1Hr8ovjnfQsbhko2fs1v5gc8EpBXRRFKDvsHtwgjhEIhMIOMnfvbzljZXjceC2m
46m4qoqZ7k27SjLlMqDQcFdaOEWEfNm8/YMYAHBy2QvgmrsF1kxuZg9r0+uDqEzr2RyhJzj8g7pq
Ud92f9q4lUhpkAUjQslWPCzL9Nv04yAiGkt8LoaPouPeg0jM6zl4lJanBK0l3CbmHql2ar+lXd3k
FU0j5N56QY0HhUeh4mAF4zz8WEvUs3CB7zXCNkuE27wtqaoSRky4kdIXJOeOp8RWm5Nmquv5qR1J
70uMBDs53BFKY+4sJfAh7voONerMeK0E2IqIrnrurb1F6+PPuODHhNPC9OKuDI3x4D3SL8e35Q3R
evO3JcYcj48FV2vYXZ0RUaEQTm0Y7CrPDQzKCmfGkVZ/WSq7oG8lK+Da20R+QIqiWPVqDlsHByHE
4ReYUY7oxaHyM1y4nGf9o0ja5PPap+jJJEhmOvRLEYF1nwW11UbcSxgKWtzFfkfzV/r/cluXN2Y4
Vknf4QC+HG1QV3iM9owbErGiBtqQLvlu1UcRQ4x3MqknAXFuxlUCBs7MDqYa7uaoPxIJFtuCYyla
avu1m8ddtY8HXFYdpyCw4hfCV3hwgvBgxR2zhEnWeZHVlRaZe7day9cMrsooPZgN43hEG49Q28h/
v34DmCEK8WGDXtgVYjceht4msHq4Xxd0i2Jn60u4LWkxI1DJMGkj2Yp0byLe+qHoctc/J8fA0M1d
jZV9pUPbrqZTI/xbSj9NYYxoDoHPyIeOJZMaN61jZ4ogPTBB0Yx5WKufTiq7uwep5Rxks545/9bx
OVBgBqfwiK+FUHRmXlokkRReyhpVXEQE81Y2xu1N+tL1kZcpIDwTVODLdm1FnaOj0cCfPSrOBQH6
yHiqK5oTKX3q4DmcZ6Cd7fOqCbN0R8rammRV5iWQFpPRtvoUP+g7dXJv4jsSKJofIwT2QQi25SXp
/X3hOGsS7lqU3cWF5CrEU0XvSlWMnwmvtF11hsh8AgydE1NHvt2zMAR9v+xQOu+FPl7Bo0DZR1CH
1rh0RzCi128P4sBRjAg25ZotLx94bqkFhjjGkNi75sb+08xV5ivG5Er7UA5LfQ1lpu++A7T33SyF
nwcm8JTVLeK7vIgZJrMTKoqMAJPkG9EX6JZABh5VBf5mMK/geHghw8d0Gxp068fNH1XIQ+M9sbD7
fzEZOEV1Y7FE/ZP+qQcZPdFP1aG++Ar8vIPdp23iQyT4H28fHFlSJOlv9hQUjCaXN1U6IWqA9yEV
QHaRL1gU5toyzAElXLDfGZ+eHZ0NhSF1AozVpNWeCyYsM+lvyADPGZ0TUA2cqTOgteNkqiWeTh6H
BN1Zfa6br1A3prHHZTcfsZ/N2HzHdjEwDL28pxeZFK0b5GJbolajQEZ2vCDPk8BKSWemo02Vr+xC
fCMAfWnBh/cNXPlanuZj2tLUyGGbj4qqRHoOKMuQzYgLcdKJha7FbgkNcL8FSQzQWztoZrCr0+UV
oBHw4cQj/55W2aT0Zb07lhbPzkqTrAo3NL4sJC3V78Mw3iqEITP6gNsyg/wJ1nz8l+W334Y6wmSg
oT+YApdi3v6qORi2f/lRhXzwt0BIGUrEsJOPT5K08h1cAElxErM/NHP+1MYJiQMuIFI6HYG6gy3z
v29aKIKCi3We289je+uZP8qhcj68q/BnXtU0LlsBXseX3G0Ig2GrRpGVBntKbboPn5gVIB5ZhIdP
P3UmFqNL7OCB7uyX4nnaGlbzZCytuwUAk6zLGKyA2bVy2NcnIj1Tfl/aP2MHRtWbzB7tvV0QM+qx
Oel3yWFj31jv0iGQU8zVouE0T6d0S5EtZmarWO2A6caDH3tvi5VTS49Ad/3bu/PzPI/x2949l3I2
mfdPHMDZ76TUvdbZ728q52uNspb2LldOQ+FJlnxdRmv3NFOJJ6x+QqhfPr4RecQgI/FqFPUJwsg5
UkVfJO82CsgvPzEAwfJ+kbOAfbl9MfQNa6uP4rLbevi3oPyqHZwnEWVRUoAsma6nNq0GcLTboUJH
ADfOpFH8RSBEBhLtcVQd+OIq6m3YF0KzqU7jyC+zqWPVNXXYrx0uZwRyvTKCUl1R0n1mm8Z2Mw4O
D52aHQtybnvWKwCqt0x1ks8vPMkdaYUpVwYU4AijlUrwAfOUDnlSgG4bgih+h7sfuyXQgToM6K6E
nT6//qcV7ObvdInmlGr0hsJSLw6EGF4JyBv6jVbh1NGuIZVdopL7NB6tWLoUJQSwG7X6akMs1EjW
13fAZDijx3fREwhhEhi44XW5vErdsY4lgwlVAkuU8SF9fkN64PWL6X4BEtQQLi3nqAXcRgKV20qF
1SuVioaSd61ATtY3DrjKDnBhRCuTobRQoZdsmcAEA0jB6ovF11pd3WQbEjFA1pzt8OFIht9SMEps
tvk9HzKXFb5tkYdEDa2qUZsbh+y0fC98zBmcgD7dXwoJJOumg3/VhkUXphqXS70YeZf9yuoVLTC8
ZG0MJyLdw6Bw8BXIhyDx6fa12B+1o9FGktdFSyNVAG02MRQbjhqjqDaRbHCMgV/0F/rGEaDCMtz7
1fC8nOcnGAGCdxHpDgHfBQ3eNlxjfzWZ4do26FQk7QAuNO5YOV8YdvrhrjAU+jkqJhAxb/nJsKFc
8hfosHTlD9t2FxDmIQYxh0TTOyO1K7TBleC0JCoLg7jGkbRp81rHwwYwIGKOaj84drTGSvGxjzQN
Bv5hrZmwiOOL2lpB4Pg//UJJ3S0GUzLMrP/0m5XczNFF9K1oFcYqEZfdIm1EN52zIQY+kly6gg+s
mFkOIPVyUd6eQA/pS49TbOk5MthvcswqCWCuhwZyV5zAQLYJqFrgd4XI9f6YcRyoR9QNi0k10NW7
xRMdoSjKn9AeQ6v74wF3jwfYYOJfOUrrPmDOk5zjfML+JWnUkt9fufc1OF9Fc4xpImmT8LFk6Ss4
YCz6DYUsSlAH5D+0RAQRxijIw8VhhnOML4PPPvJgXXnxiALFgGGFDVrIQiiKNhr2dVuyOL66Wl3B
XhNEQSUmgabEhuXmAN+5CpTGNnfykGloyuBkY1cH8L+Pfx+Ayonj2QkV3j/8r83C5NggjgRnx3WF
7SxRgXk3HD3XbogToDl04RJWOxzcYYlmyUcP1T75ibptCIGh24nQx53Lsm5YuxZZAdBMa8kplpPp
HXiklEUy3fINlw/4C1Rgt8FzacGgEr3AgovwR1YatMGfybD01ESKAgCty//xv3wTby0Qx/Z/5Z3j
rEoS4i+LOU5qhZElO8Ba67qKmkncCeCNjSUTwkT1XqygOd2QRVP3+PR4OwSJes+b/69hcGZ97hOe
0COktSD1w7Q5/4alSxE31MDo7Tobd2Kygwlv6cDIMOb8nnLRLn91oBv8RQk0Iy8ouBj/1wAfq97+
JwE7s8b/ETF4qNkTKHm1zWcuBMmGHVukwP55Qu2Jw8JusfSTKPCDvLv0ZNugHOnFR/P55vd1G5Ru
quMjzKDxa8ROz/LVf/rAd4N47iqZz0fcP8riqTnS8U0DCNxzwWzP+WH48btdkoPy+Jdu5JSbc2Pb
fWS54aMNj8YXTCdubXkp37Tz5aSPFsUBEzVpzBGCPBL02/lHxvXtySbDhj0eJebTOICgYg1oaaxJ
jKUErlkm588eBRzK66zux+iZ3OM4YzlNlCbYIyqnyxHQkEPExe+i9jvJn9i+NXTTYALd+zvfG1ru
SvgpmtAVbNyrUAlIfF49F8jexZ/hLk/iKwZk7MF0UlFyVeTdAYXFlCcB7o7dmrfRTWxMHFCirTet
rj9LlIvcf2YzxisTEunz3hD2nDh0XaYELfT9EZwuCSgC1kuw3JxfqwXhLwDErL/jcQDx55HUbFiy
JUybQgXV3g5pv2axYQKBzJxSZjLEjAcfKFwdPA1ddeHbKGSKwHIMlNGUyiAE2s6UdSJ33HFa9uwk
sG32pIs3d78W8+EkSRA4Ko7FuQBJeKyzVzPDFi9rx5AaAywWtHSEhlu7dAYDcZvydKJXBvfcHtxw
Ypee1ed4YjCu1yjyeogYokrRs93qX/Vb8g1/IlJlajS0QnPnthvkiMd+2uq7HsNFE0gisgp1Ie6h
89sCzE6TJYJg2mEfbF8BV0Y8nDhYwkTe7Ka7QzMNy0bSA3APF2Yfw907qCJVx0zoYPUCBvaJkeHA
FsD3XG7rV2exyGmYC9fVzzHOlW5/ZaMtUooL1pTjKm2jPitwoLQ1DnMqQSz7c9u2vGY9pNEtHO76
Od4uAti02CDbSCimzFZvH/RDqPANISPh98Fxt2lZoqs4pM31WEr0aeCaqkEuWHKZD1Zh4FiR5d+J
QnS4aEXwLahJpYxAA+XYFo3XZ1CQhogcyQx1Q5tRZ7TrqhLTgNIRUWZ5mCUOl8u1vpCgs5ORt+0+
3uo8+eHZhfyxvu5k+FB/M716jKzUnES6YHhGbMzM3hhKqBGbN0E58X6AdXuMYX1D9WwOpvNNhpdL
qCq04U8QW8VDbHbDsi0m1jmz1baYSNQ4+VTl8AQiR2sC31nZ270jPwYCvAAQ32l60l+SWdrM6ZQ1
oaCNJLVPppIBb8kZfKeGNlVA1HjCMTDPdMutOELBUS3BM+NjGwkLhgsWcfvmtrzBuC5OFDCyqYRv
ovzYv3GRnFQEgF62sPI7vEVcFuKVqHl4qAvWhI+KwiAzipsgLLfZFxRfsgxnZKgTgjRh2tjOG8iW
A8WyxND9zWdrWmIl7vem8UkFUXwx6vlk8+/VPkCQfzLuygpJwAg+h8ubZ/MSR4D8BOsQs9JzSUkd
vxc4LXrL8RkT/J8WLPlHrt/dlnKjsoKAVOJ0hydJv9jEztAJCqOhxO/7ntwwf215Ry4YzUU99hR3
u07quBneUfLf/tuJtDA4LFFdD2Lxw3gkSeHddyRcW+OWm1PIbWyLFS1Tpn9xSKs53N5Kq7z1JrKW
77gu/5xHVppFY0w/TiifzwXQ7D8MHohanBObeGHLr79cvOg6Okgr5gTt37pF3143Dj87hocu3RKw
Huoxw4TrVH0S0ZmEBCmTSP8EJOo+ILpxkfaIZwx4QFbYB+5L9Z6w9F0SRGGl17xGL9Geyl2VHxwS
c6TvXmHP6w4o90d7DdxCGuUA8m/gHZONEXdC8tIpmN2V8sUmHI3HuULJVTJXO9zEW/683qze9asw
m4Z1g6QTxR1IDKfytEJoCev1qRI819PR4R8p0HaKvypvbA3uSmesXzQLVEm8DgEHmX4PzZDinmLW
DS7CHJ6sjkaCBWtCJ0vm2hW7EDVYSrB8+ceFXoFkoRkcxSANbdzQtD5zKydqVzXP5JjY/K+Tv9bI
4i7RHL+XK9fmCsmYwAophdUABWKQFOGb+iHXPD605jQIFSMhYB2NyeO0JcZI2r0fycDJw0vCkv4y
eiMz2/3lSFRyyklX7/EqQTJ2tXdlTFVL56PmGejgGpy12Et8WUYImE6oPTubfmrB0NSueSyWz1MM
ITHcVNpv7E05YuuATGRW4XUJYHJZc0QAnoT154rNFHvDIiK0jngZvXrvKTufGuu6KSXipWqqdPqI
AN/TLXRODqTs00kHtaspy9jLRMSjq2Ps01YqfsVe3jpkOW63d9MY+aeBW3H5aEvzUu4FQeg9coCZ
KKXBT5m2OdBiY1MrMw0/uo5VRF6vVszJrDNERJ0rWbTnlIil9qWEYPaIDtjXjVgW4jB+65V2+Lv9
hYlVj6oQdnj5BwgAEavY8Zch+fKle0lB93BIJR4zr2ufzy8sXVz3xY4upxngAGXvXtRCEeQ7ZR14
R2hPFwsUV/2X5aWA8TpnFD2y5DRFq1IL/mUUh0QidThe5/YP3LE3KfycvIfOxxBcrdB4S3aQBtLo
eTtdCqU7d3vvNSNTWSmBp3J0HrZbk7beQGP2kovPK0BX0ipRmk88VVRVVhVy+jemmlAIOc/32HjK
wvfVXOv6fGA77NOUBtdU1SUlJjFbgNaybi/S3NtyFY5HX6a1nrpEJlnr6tXKWvt7ZggGawjnlqCk
y9abADcSOK7hqisxhcCIsvPPSTUhNKBJflhX48FIi6v9cfnAsGdOHAvey2v8Wh22ZMAEn8t+0gjP
D9DNFaHsb6CMl5I3E48HakNPB+L0PiWeIw4FVF1P3SFA3JYlXLui7Wv9p/vCtdTzLJOjXuO8WQ5F
tBtVMLhFr7s07cw8D4WFNXE8vUmm3Y8xa+Zrg+aUZOIhkP+ltNCnN1SF0uJbXJiuqcL1t2TmjuaB
m3tVss+JdA8YwPF074DCL+NHXEO2YAaUYvEVThIQPJKJ1duXhrVwHw3yoIRq8XKUceuyfIbFSmUj
Wzd0NCk4/wR4WUVpW2aqAXNsZGYAwGzAOkyRewryg23kyF01+DS2/TzOd2mBeW25+6NT2Kiup5sZ
smRIRyg4FR/gBGWpFQ2sYRQDPIaqQnvQOVwqx04Gft+fweno+Ir7RwhjySrP4lkjvGE/VyAsmrbp
9Tsh3IAhNeFIe3z3t3fXCLw34zdhkyHtSU/AGtTIPaT7NpKlTKz9H9cILKF/ZI5VEJc9zHf1gW+Q
9wiilFRjA24THO4N0PxVNBq9wuVb+Mgsl2FNhHd8C9cbSIZqsbLbrSA4DY12x4TXKRwItDS1eYOT
cR+dGiU2xftBy+CLbIxvrbebWpHM8bD9+e5tzEHysfgyoranrN4DN3newfA9BRXAzhW6KrN70Spz
mF8tqZc3Y14PjW81LjPeWvGyqArJbP+Nk+hjSybE3FaXrWEJkw05Vdv7Q4mIxUy9D37RYmf7gMeG
U+u6S87cvcOqB/eSIQF5pyYun9pQFEqnmEuOIbXtzBDbMnYaA0YoQ4ZxDnFJTD3lVc4CHSysG2XQ
myQnOcthO5qOaRDMWW2CP/7lNVhf9THM2MKSmXzg0cK8NtgruwoFOJjLEyFM8ddRrpkE7EepuSbZ
p2UwwkbBSCsplWrb5w4CwHh8segz+KW4xNrgoqvzI18s6iXRtzxppdadGUhq29v5KxG7SoZmhbUz
klr2CKQuwFRs9V7Hj1a4qdGaPuSy7s8Tvbe42j7+UOCS0BHI0jvHFjOZkSbASmtMaQD/7MNUx/nQ
M4os0OrmWa7OfZQXl1B3V01hxSQ0ETNN/ZPnYj52cT9E9rr6hKMRn5m3F0knU+zThFaN0g6SHauM
AbBV4ZjYRFGW3cxZgfnkXIJGgsVYW5mhqVMA1OVxd6iz6ZdlqPRaHYDRb5jYOi6nOPPutJi7KJn+
Xf0VKX56t/nwL81nR+eV0dj1yEsfpbCJ5XZ/IxWw1o7p66OGIMQo3TKGNAn5Jr3DCf22oy4EHnBu
XEv+LtVsd8iCUh9YRyoAbX5XrnZ9UuTWWn+q6CKXvZPpr8nQG+EiKalMW3l7Z2tOsT6I5kBByV5Q
MqVZXfKM5ka19hiy9Tyf+WIN2F2w/kjADzyZOSehGxjKhbD6ClTet6cxOD2lOMzkDeukjocPfVel
Y3zRyRc1HR9qRrANgw6cfW8SKjzqkEBDYMtVm/3ugo6it2IqKlE1xLClxx8Cg9QlOtGFGC4kSIQH
3R2GY2GBVUlZGcEgKvjooZD5Z+W7+Big5EarK/Y0Ttku6G2nURlyGkER1zHcGqRG5dneJqOHd0hx
6cXjEELJu5YTUmp0OgVaPgaPgIiDdtFgf+3aGommrE4u73iLUJRLgGsRSj+1IuCZV/FEGLYoVdMf
ENaUX9s+vGsR56TXezMVbjgaBs/eHn+Mjxd7Ks9aYLAKIX5Oxgmws84crjdOaXlxqiqMEa2sHzzA
4u/mwm61k11DPvEEjA5fgDsfPRy1ZUrnRmJI4eCeSoQIkG4ePcM5h+Yea3pQuPT4WtuZ4yNdon+J
sd6yXNO8yjc+gXTT0Cbc7XId5vZRRQWt46yONJtoLY3Adj34U9NnPlA7Z1r2Jf/Ta3c2My6/5qZF
yc4aywWUXYFDqVKYBqsq5EmgDnV6v8f1T3rS3/OduhLd7zlK01M6hQHnx/rxVfvCPSHRq77CNM/m
PKMz0frh+bB7OqgJNVjrcOs4GC7CW75p239K3PZbs4oBuZFvJv3/CQD5RNnAi/0xTCE2D+ozZZqu
koqxdI9/lb4V/e4sUut+GWAzgDoz7erareFA42LzOZkE66jEZkOMRN9DtXsjgF7zLzyT2/7wf5Wy
Zn/bzCsQjK+VfYM/UXAQPeYTZs0S4bTPk2tUppOMJZiDMqGN8J0R4C4zO1CWCvOAFxOZfpXHFVwm
FwgPRThSUdrgTgxRiEHCQx4tk4GDFYz43QABPRCFH7HGDfOVSFa/16Po5Gdppdq3VDjlmn+/MckI
naQLoUTX9Z4T8uhk91DHUlPO46yh6ZYTaO1avf5vfHombH7kKMVUBBitHcN7+aC6STfTuaH8/Ndr
Cp73+M97vOknyMPFA6rX6Exsdav1XpIxUMPiVAOuhG7Ys8fx87YRgknq9PiPVTl1IW5Yqg83BY8L
rDQ/AQqszplGr1iCSsLUMPGPM9BxKGDPXPe0mSgbQnklzkmOEbvTZ8FNMxflu6zq6jNEoFr89tnb
cS6/ydTH/XGHrgnK+XJfMJF29mv3gm8nE4iaA9dOvOPXWxRAav902pmWSi7OWo5DLQ3JjGaWqose
r5g79t7aqmhcMmvGRwxiSn3bRtZQvtHLBy/8wkSNj9itqvdEwj+RePTMmSoP7aoJNOznXM4Iw7Ww
uKwGIb2qESD4zjzlqwWa0cWWaCFTqMvkN5tnKZTkMWijS8Gkf29LOKIy+TvbXxg3m9De3/hELImg
WOgDiW+KULsKzDfYQSN3xWRleXJZwgARLcdyjm6U/sRqdbbFPc5VbJvy/NyaHD4qyFlRTglb/hU4
bMiqTtsXmCQybqrme2zZS2xdJklS6zmQb3zehunVPSL59E2AXBh0AuWRH9+IwMbzWln5VeLQShwE
XgHcWC1Hh+LGFFn6V4mgl2sSxmJqmD2gifyrhwPNMJxYdSINKhKVy1gZK13fK+/GA2GIn48z2Fyg
CfyiKC8Ht8qe5Ig4xr8s6jVx6QrWoj64Qe5BxQcdCtco49iq5V5TA6X20xzNyUD3JXYnFlNzz3Wl
bTRHpPw0AfQgWk0/ot7R03rnlShwRgqGRmZejWeXAF2XIoZ/UWWjsUoOXC+5qUcZy0F4QUlo+/te
I7hCLP1GKYYfJaUm8at6S8w9cDE1iMp0vKHYu9eknUYV5YKWD6ZF9BbcbFl1oBf+Ad5bQnuphD1X
+XSwH24flZ9UutlAO9cSGJqtQNGDN3QEmm4oy1AgDZRcy7M77ZAoS4Vv7j5WHeOKE17tB6TpE6CC
9CoC0Jbn73XR9E37o6CIyk/2DP8JZ///NoRvvm7/j+TsQRTXkkek4c+U7IAUNXEhSXU2FlYMxPTL
vI5jBiGA+5TrNuBPJf1eqrm71SZHOXpSO2De3HRUaPdmmgebKjCAuo55ztcOigcgyRvfPY82aad6
DKLI3Y+Y5JOBDalp2E/LRNxS4xOEUDTr+Kb3G37Wvr8PqJuVM8snluykykI/unAz+Ym09cKHNDCe
0UkvN0Fovy+AL5QqtLgrA6Le76ZoYrJduR7smHVnF17UqatCuqhNF7KTz8TFCEZEHEAsKvxkXMM1
z80WMHgu4yG7DQCrBtTPbab8Ij49NTzDB4l+lmUZV6qauFxuFmt9Fh4GxJ2Lqp4pjIhkw/h0hJz5
B5itykxY+rhB8UINfv5Q+LWe35jrqY6TFrD34nAqes1G5PTpKp07k0Iq+L6J9foc4jWVBf2UwI2b
pn4Th1fQce2sADqgNMWaz7LD9wTFvH4bHFIf5sQ+rZgCz7QB6a1WXhihdhl1kHZWXDXZ+v7wKpQt
TWD54AcXZ+dEzHdiWa/Ec/W6fIdy0yQeu052TcTOCd2gKg5Y74om7alOYvJoMSdRFcOzcgnCBWVr
l2PDQ6rwzcEbVkg8zDitXSxxY8csTrtKAW9jjXGbrFAXe8oT6zzR/bv6xYfZxoj59248Wzzv0ib0
ddiF5KR8GOtOldQqWhzWm3ubRCEWsuV+j/jrHycZ7PTCoRUG9u6MF824gqTcomSNE2lFvMDj7tLj
mQP/vG4djzNs0Q7/42XUiv+3HOiECT5eFuO+qCxlBI3/vP7l/rbPYa54p0xiDGIyvwCvVKh0IEMY
4NW8t3xcS84RAsre+gtqZAG+EC2PV3D9gHADvWeUGMuxH7Ok4wQMQ2yJRmeZ6u23+1KGbQRTQ4yY
sgT3XIK3E5/9z5waGmpgCfijygwyFIxiyVwP4sIctpMUJuiSitN8x/odVgXzFayyOc4SpNQ4mGp7
0VxeQsFr/ixts5/wRyflgDJRrYuUqc4dVnrA/ihOgI7OIsKulJB6EuY/veLJ7DbpCdip1d2SV7VB
4mvAcVBMXl9obIakct3HoQUrDT2OY9HZYOOhjtsONTzzgwiuNl1hihwFlKWJaOGG6Gvy2UI3jCdT
bibVUF4xPFH1es14me90afFzXMn2LGADi6b4U64sJUmtf7V77hpiH14kaUXdU8zfVXdtFO6u3dxR
zqRbgaPsvTQhlgHelzRxvuSVrfF8oFXpetMB89DqZ8EdmLmhfjx2kWDS8me9/KuETtcsONuhoWw0
Kkaah6m1PQVqDqauKFxBUZOreL1c5EOY7zvIG4aLPkB/EmoaKWs51JPJKgQ7z8ZMalEgZvcZ34jW
totq6yqw/3aVU8UATSa7aHY7hogyDCUlHU1HN6VPIt45F56L6GesVN7v6IJw3Ec1/F07/A+xRkZ/
S6ZkC98f3otq3v6Zs8TA+QYk+jh8fafC+tT6TKdBwoE7EGOvgBbj46xFG5I7HfpWfGzMVGd37gRJ
4U1cSpbLsJOeGhrwpmCZn3MXt1fnw8rNKiQuAPIwkFfjrOdu42667c9S5oR2KzFIGWWjHOnfapnk
6eLhP6zeF5PQkdSGWGMRJatFoFtod4aBfsgYBHAtYtqXDQGCPn83s1YhIKfSV1z2B+PLWY/WQyxU
GCTKTmdgGY71wvSB+331sKdNY5moageeeLKmKmrCfIrSLJkMlc3KxjFQkZLXj8Q/vkJPVFbQxaR+
bbugo+7KOgC81KJyBfN823OnXd27EdYFCnovsR3miOcwFw6fzF0rMeFWXmvPDncLkTX40X0bukdH
rZodZ4gckSuqI8khG7JeRDmfOWB+tR5LeGUJ8sXcnTjSlmaHfCxLXzm07hGitGqJD9FxUBFUFqUr
5ryqP1WDmlng8p09MwiKY1ojRfyy81eU3fDUHsRsJyctwV9TQaUnOHBVFA+QMATEf7pdpf/BsX0W
s1dbXHKqMWMFsdUcHs2eb4oQhpTu9g3wds/ZLq5+5frbuwk7jEpOvcfr1v2oNju6DrB5liTsLTs1
2BNn2NHqBQC516xYQ/WdugCbJAA9SA3JAndHv/7Zb5Lup/fIgUafmt6xlViN22GUk16+6Ut9c3L4
sxQarHNTJE307JBPVA0SzfaMRUvgWcekYILTO1FoyWqC4xcqrWlVw9yoth2M7+8qa77zxfPOvRvH
ucdemnScMuRj2gLB6ZgElbZcukFw3FcuZuyhTX71QQO8kBVoyBHEcNd0MMUGPKLO5/nv+gIUYHgy
ZRDbX8t9FfmOuQEYqo/dNjg9eLCu4fSUXxNG/lyKUeBEcayhD39CvXYk17d1zlA947Q9V5jOY5Jy
T70zggC/PmpEw7mHlf6vzlf3iW6LicMWuXJ2k2KSOW+YbZ1yLYIg0xFuriBJnLXJorRosF9B6xpz
75nqm5Itt847+08MwKezTUiVtsbFWDFe5So+t6S4vQl9zHLXCn3wqH4xVSQ+E/DavYbkM/OgaQKa
s7Sz6NzwFw6xLw2+CVpXjOiWwcU1Z6ybcVSHxuMaLdWzb8rBdv6PBGN8Pb5FlMhRgxlO+AwowMMG
tagD0bDhmrN1nXGGoOTTY4Yi+k1cb2i8no9HZlV+9aGaxvGJIOMfNGMJ9Y2xYFIxsK9guTS3cZ2N
vw+TtGKPVxXgTXrUdVSA5tHrXyYQ/l/8rM9XfG/3PrFZS/uJ+TZ5p6VIWhenEyZJdTF7ZUOvUmcA
yHEhrJqKtSDnmS9QNV3MXzq8PVvBH46Hj5iKDZ3MsbYcYk8j+1oUIyCzF/cKi6kW8AdYRMVCKg9C
leiJY2fUUAB6hgS58x0itxHbQ79ZBhhgD4L+bHeLJE/rNh2r11qz2S0egDPlUpRgLS93agC6SuXb
+NZXxZdxEqnoqJg/bMHOyt9JZt8iwFrymEHxSLszRHqjV8cT8DBpa/5KcLbco8yyfxJD7nbc6bjJ
cqODzTvFxVbBErXAk2Ej8Df/ICn4xt7Mv2IzjDzELjh1v9zIBBXJfcQ+kgN4/rMw41tT/drS5c4X
5L3XdWGGjmwjdIeJ/jjMkHIg/3Dy3Y5HlR0Uf+LyVAGvhHCmuSrRLilqGmc8Lak8YMjvQClBKK/S
Aj232Rr4x0EfYgM/IxX1tF16HO9zFMHGFDrBDZoCQ5LpI/Bx9FCTgNKZvr2wWBXJ6D+UCS1syNPv
LKl6FvWL3ZNiTGg130/QP5YdlGbvCxVVOJNexyazj/jXSV0FDKD88k/OkZwhFU1AaCQDVxAC0GAB
yrUZY6omvZUgeUEXJFtTrZBY4OYhd2ee4lQwYdCSkees2gUZzR4zKik5jsJUzDLihE9e88qvdAka
AMSFF3ab4xd/Fr8PdHkMggoiMsecmbA8ZA5yMNexIoOQEcGR9qq+RbI7g1RwFQylXrgSploBL/Mr
1TkVxgt+nJ2zjOgLUyBIppubNHvgnFZpwECI4bbp4sRYHEJfn/UJoyx9YarPWHtLMc4prERylSo8
I/4M52ynJ5CGbN6ykYN36ZWP8Rr/e1rJAQB+pAL+O32F0k2BFLdtuf9Dvt5XPkdh4nJtQgz3mNma
8M5MObWAy049TT/D84AGoASwk+8zSkpwSF+Ld0i3E/LrUWFrHJairV3D51/Avqtew/YiPqt3QiD+
RWsVJw12LTp0kurpFWM4xCOk2dvfCuOAAU5ZlbcOPTaphMgeaPuoiJll8A+adJxIDWY17OXUtKAN
00tmyUug61VKU/yEMQsOm5EuHPLomZfT0U8vrUjnG9YZ5pl6jA439odxySO4cIGQ7OQjWkWJNZ4p
zIT1hW7yckmVvV0rvkdOSAEvGn5JXfso6NG5QJmqX9OYn6IyZvn6tZVCoUcCXv3Uy3TeQm9MwxSK
ppuCFz9vDYVSgnZzTKkodUHk244rAkLvk/dE+YXVF5V43zE4irFKAVWSzVKrutOzVDpAeaxe5E5N
z3o55L5HzOsqeIj7Ry8KmMEMLJnocnC54FuSjXrlAx2tXq6AbSridpgIkTy5pe85WWuRjczjOLB+
p+5B71WqBlFHBcx+ZWZzJooo7YX2wQPiwfmIxD6Q9n/RrRYnqFFqjvbEHn+Eph8ODLMjT6RbuvpR
jZbJ+5of/F3vXr22cbnXTbfRYde6M4dvYIt/Dtloma+Ig2UN2qOAHDWcSQ52fKVHYqhJqqxSp3Yx
6njpa9eslxuFVRLhSEf6kjN95FCthzFNVIebhuLDNfNRTpLUAp78uA0KwetQe2i4932pQzTp+yx8
KiHxaPz4vRaaEdY6LpeTm0Az+BqT9aOcHTj6A6yBCQGxZO0lcwFvirnAP8MJb8ESY0kyMsLAqMR4
Hk/tCJcsei6ABLjzPjl07yrR4VEc5jJPdkdhMV4fndIAzwZn/RdVCa9RaFX7hQmt5iUhThutvbFd
VFt3hZ20NjeB+lm+WJUTUjoZ29/uLkdY07lyXIQvl1hu/B8R1hxGb7IwLf8H4c9GMS1hVgam279Q
+bRW7Tjt3U85nC6AbYIQgEDAe6wyph9UBtYgbzXCWprNEiR+6x3ij7o5rRqiawrW6XixdlS5cTXP
fcfudMkjk4kv3uP2zu/ucALHucvBPB+f1v6VvdJzyLW+VsPRFrFHQ1/qxJjGea+ngac4+u35+Nd5
CB3EXtFk1UuRTzBPLlsNlf77ncMuma6V3KSW0pr0ZKIBehFms4HqUxS6F6SaaYivzO5GjOA6Ap/H
ka7fdhwxYV+JlBO+b74sv38yuhOpl/nd4FeH15gqOQ9lIEYKMl5IgqY1P5QEGrpwnUJIPKSJ6eZC
a9VgqbWHofziXefTnpr7XJHmMmGCOvMeufkVr2f1PulC10JGt+PRNcVyYgzPjYjjVQslDne8G/GE
PrPrVyS8devaM3z75upytmvbOze3iRamrqXhSfwDN+sGZna1Ni6dZfcIQyq2ybHQCxx5Sfh0HjV3
17LckIxhJR5lq+K26Q9+mw3bOamI/xzB/cyzx123pmYT4tORRUC3/IGfP1eR2s+PDJFj7UXB03LN
ohPWvZFyIa2BmO1q3vo+gU4PD6tkPkpiXbTFpBTqBYyuEq3WjAbTQV0DArD7kWzT3kxTKFtcdSb/
Ut/YgWERMbGkq59As7IgpB45OCHu3cxiSlYbjtYY89NNOMNyztAMyFhyD/cMczzxMz4PA/PKlITU
svvKSvgrOgxN48DgNrWC+riE20lMniUpDJu4J/HvoC23vXDzf9ykQf8XLYju5JfOlOhD42P5CWvq
G35tkmdbicaW6ifAHMLC5GpAIylVfX3ZzIbV/rTaPJ4XT39xOPbJj/W2dS1EakHmq/NN19y7AZJj
0rmDSjGa1wyWDP67dzxl4pGnkveYIN0kKLRRT62Rc2RjTsjnkVLqPUJJSMPvYesc9hPmGQgBJH0n
wNxZTQDsbvFnye6u4HP8Yo4wuq201nR9QDR5ewpN5OpbLQ+0ZW5MRHFniah2NXf6UnJ9Zp2XGaW3
KBDbMUFLo7WwfaCyjQOmPdC8kbbQHqEm/SwIJS12Mk2GtkG6jzod0KRrGn/F9NjZ8fM6uv8uCKvE
lMMgwOIxmBI/Q4JXNOtnXChTS8vhqUVZlJIsXVsbZ/lcEZ43wzvzneRCTd6AXnwdm/XpiFRL3zeq
7IhfmBuBUyYaDa/eJPXVxAvXSdzfSryCCvKKVLKrT0ygwKpt9PrpI62wX/NTI9+k78VUCqKIsjva
WAYdsCo3CZzpXU2jjKw4oMKucsLpwEapGiSLoCNreZIxevgri2Gm7AhHrIP4r77RJa9qA8na95l4
Co5om7Ua0ZUsnq7kBhRTGW+rKQG6RzauuaHdjgr5o4jp9vVYzTYmDDPaHJsyODtCzldzYHKt8jPj
pPZ9sHCNQFxMGSzT96SuNtivi1G5/LGKrFnnRMeTVQIlgzK3e4cDA2TxeIrJhCVtydCjraRMoq97
oG1uE+gpCh++5iw2l1pjNLIDL8dGND5WPjYaFWk8Kcv7C4y5l093UNAHL+37z33SkZgIEcDhkKCI
4ZYCH16pFywAjHxHLs34tVKYRJO6PWcvXVcYmrd0WILooPUxqUXlG6zyjj7ssgCYZr+z8OrxCDbK
TAh2AkeGxDbbsWmmi+iqx6lTOzijVkN7QWWporc3UyPdyTZKNGFPIzX2iiLeHJR0Ic0LJQIpc3pW
7NPcv0aclIdMy/Ia/gNfM3c7AGc173hU6sOntuttjo8b4g8KZI12Xmx0qBO0/1Qvq5qVxj6R8YM5
fBablJNrVSicI1kRHbOqAKgbFYm+BhSlfxGCI0KaUJ0MQk6vEsW0sWIkla+ivz2VigBQZkTHT4m/
9aZwiHciltpPAQC1UmoH6ZXFOE7pSnAlOLbivl/JCc52wT+vSQOWV1VKSfHt6gDJ9p+C1wftqMlI
NCHKPXvninnfD9ddpsbhohhY+cZ9JmrEyafY/RuB2cRPOVV8SPr9MTplVQYhjWHCEtTN9Zle66mN
N8SwnVJu5nJRpDdqAEtZ7nALW211RHYNUcvEAOFq73lIiDTs9+x0aNEzfyDKSkfjDb5lKyisPrTY
t39pZejcC6vgr949WsO8hzc/X2sEYmA+XiFXrNFIb8s6wnuVl1gq20RgBNH/Tsm0rsilAlxY295I
v5qsxzZ94dbXytB+SdqZ7gLaaYWUD/XTcHKeFk33VpF6GMmSX54nX1Wd9t0mueOGHN0n3HipisDs
+w3q+FtPJqR/uIk0sIfXvYCIWrs9B3uxTMbJd8DbT86bG9fvDmvbQgn4FI0qXYXMYbD0ZWEPZK4Q
vZ1C9jVPXJeWnwA7bNjKTenRwbqMvjJQRg7x8apK3cmNY4tEfPAUeZlXfTbk+wr5Na2uynPONNNL
UOE/M17j8Zz439Tvqs3g+N9XENvWejXBOwAatqsJlAyhrPIjmEfSumWwtBjbH9muKr8Fe5Y8KFqa
tsad9GhoZjfonLNuA6UlBKnTFgs+X5SI4F4lW5T0iRxlQU4fn0wqqf0887i9/YmS/2IFIkZSqwXw
52pgeON8QYbU6XjackDCH5Pvg2wyMf5tH+otUVpSmmJdPtmcPYurYH3s3/s0duII3S7XZe1oYg/l
/X1De+pz2zHtbgaS30H4jXRteFWpLZ/nCncpkRLwum+WdeWAA/7JWcEGa44TXW8H68FM4TWlM6nB
XRH6+3AHFrBWewiYBhmIGiwg/s2MqwQ1MtJ7LFeJd/rSxKLO0WIHdFmjSgOBrT+0tjquvU2r8Ze/
1bYl+/BdEYE0srayzr/F0veVfz82HMfID264dZ5hD8t4ReIA4sEewi7LDTgcUKvvOI5n+/klwD5s
Tx/vxVII47VvFr4Ad61hRAommbaxDvzkOXNbWyzlmH70NmNqX59GFDSKaAMMyyV5nxSkxgospFFL
wqBMGITjNkAviHhtOGN4o0G7OlEy5CQwLbOmSQDexWkYHX8/7ncnCYAzOKGsPP7yTfGEznDtF6Ve
ruuI4AQ4mt0mBh7ayI8fuu8I9o8VPsG/LsXh0huxlO69YXBUTfywe9LXdnTcNiAaMZUaDXwFhK0Z
iHXs6AfeAW8Be98OyCBL+M+Ge8bdH79UwpjXq95RLHbp6xEffXszs4wNpq74QH2fMy8tGzo+xiJj
WBVn9ji6LvvIVB5XiBx4SmwRjDsbe/mQqgxEJCysMAXqAG+OzsN9ib50q1zMbm7FzvMg3qEQLVhb
W+cXect7STl46g2qYN8z2zQeGZ/Xix7hhJdju03lFKoDWV0D9Fn/BMg5yTEUxcOItEQCFH6ZwSa+
WfR79ClMo6xvQFUVOgaCeaXocEUc0WgP8yRnXhGhsb4nOsBacamP2puLyymq75K1c42ke7h1VacC
ijegzfHPj9o/ik+HAHPWrXglK+Tx7uoW5rDxycH6WPv4xIN/xb76MoiPoir5JzY8gEl9t+tMIcAa
ztwvHdmZk6HevxOiS/AIF/210dplrWyUB1KmZ6z4j3DizGhGpfIhvljX+1WL5SURJpNKG1rFbgx4
2IP/UUC3jYHlgftxAgiv3UCjBhd5EXVAWYINsNInjhFBJ/tACNzbZsQIWFiEXFy8qb0ydhpK9g74
dEkOL7OB4Gx7UD408G3fpk08hp6bD7o8eTFjirZEOBe+N+8ekUHuC8Bw9I/8smRBld+v9qbMaaqh
2ifrr+bjrXt+GdBoQ1a6b9EzYsOskMyGf2ygx87nTj6WxcOiptBU9jPoXsignYW4skVr3PdZDdIv
PRcE4ZZ/qoGWQyjeXfwd2cOLIB5awMLu+MXhfFx2PqHIPt+F92WN7JuI6pOroUxrBhLJahWrzGys
8clYn8es6MVXe9DoJei/zNn12FDQCIq1ZSx8iEaDj2ViGOLme1HZPrCSHDU8Hm3ndm6mT5vxiyBs
sUVtFai6M0TqTsrYWCqAH7bvXZi77E5l2lENCEhSI0Qu1atp9AzGpEyXvamuYR3REKVd+W9w7J3U
rwysrwM3x0cuP1xmz+urrRtQ9+IklORbHAIlOUU9/j25NLWT/F4XYHK3rwlN85cwyEDf0eYrpvmB
Blcmfpk2cOB4x++kGNrdYhaZSh5y/WWP33a+KRVerUMelpirI38GLjanyEorD8LBlLy2sGi0ZsgN
JnbCUibQwNenkfOBLEJ2XXQxlePq35OB9BXKGPCthieGIuq2sCyhCXi/0u9++FxaDOu2i4l6GNQ3
ZG3yp7oBHY6iJKx192qLD3cwDDfW/RnOjzHm/qTiP6gZoJRH4JjvMAhXFyiKsXjGXVnCZnxV1Ppt
JRIYh5tr5h78tz/h87aDsmyroL2tiOmOHvfXEndHz6dOdwLqzY6NLgetutBfahLaJBRbwOnHh0DQ
zjRPuD10TH+Sfk/c4GMEk6v4/eIAFhtWOmFnasRbcal8KePFFYdtIk2vJM8x5LKALuIJK4+3xyO6
9hKyKA1ZmIPxf1yNZK5SgmfhM5OpUr45imLkaSQiA8Tjmfk2Y6+8EY8a0s4vQ8/gN/ZPhEO9aMtk
flcNEpFQyZEz3pcUnBqtNg+cVyGb3J9h7LhxgJ9gHHoKc1R1MSF/6TBZnv0zARD4dv2vJKYCIekz
zbY8zpSFFeMqFJi91j0EhSusIVmkcq+vwdxgEKHQ+q/2nrMRtX5eO7Kx2Yvdf4dmhdYtxY9iL0JD
x3XJJBBOJPtHhCfmPbpghH6W0Lg5e7tgzmEZPh7c9uu/Gr2mofhZBI2eB0H2JvEyokqh8pLpbD92
gvVLIkR4PSzMlN/x+2MfHOLtjribRIbh9K4edJ5Lcgdyl6iksFjq7fY/yv3evyRsfmccG+Ai8EpQ
cwW7Bm1z4g/pHnkcj9zR02BSodHfgD3sexMLYQVMtcvb+ekcZI+IwIYWvuM9mTlffjGRekdDNtRl
HYNl+09AK7ctdWXkxREjerx1UxfeSPnqpBQTBpyPm1883GRczd1t81PYJOcOfkXHp9RXWlYNlyQB
2KgczoHM6/PUZIHOowVMU7zSCk/bmbtwwLfpK4CSWDLyUoVaPGOmvBAhr2ZVVEWl6rNvIHVe29tv
Vke5SN3x0S4Y8OQtC2Ghgcaok9SYVUnHG1ceHNM9jrcxBbQHR+IESPbLqwsz7tXt+hF2a5exPMy+
E0082d9SebDqL1abxFoDYaGFTuAHTIKOBRRliA0HmT2YW0d3Yy54TDZTuTLRmmripyXcNzyU1MaV
lHP8/nSr491alRlKU2N7klpYcTb2aPY1BLAE1HiNRbIMHtwygeIAWPoicvUI4jVdWCbO4NDha6jh
rwbCnmQLhCBtra0NEPwXZnXrZMgb1GUkRTxs3kvTFNUT2V2jGuF1nVYgRnaeJTQarorTfYFUHfI+
mumCkdrAHztNWSNhTT7zt8xt4xhmT9uQGubKsTvT+to+7DOBxfUTSNyZGYJPo/a/wyYDYcNeU3P+
AbYDJOKnfnqS2I468iY8LSoJyCU1/z5aeNYwFm7L2qU2hUQh4Y1Fft9ON9rlO64stHRSZiVtv1Gc
/W3KX/26/A9rtjVwqWxriCPqDiLx8RMHlQMSK2yn5CbGDNnyH/JoMxy0yLWS2AZkT1Olxjiu6F9L
26j37U1e9xsqKOLdl6QubGVV7dJSKku4PIWfbvoMnjfsi7vGqaCt8GzOKybKqghKDtiqVjWieZ41
rw3jCtzFBbVc9FFZk56x4t69WW9Pa8qasvJv8AhlYQenxF+d2kLU9p3gJPkmt82znOfl3Vz+zcYC
PkNtm2x0AlvB41jspDZYvou2Y4t8017535l0MgvzgW3Uz0Hu38sIexmIY6T7NCxmuY4Z+BKJMIMW
6BYPEFHSWemDhqPZO+V8j3ubtzZ0S4cfHUMd5/6GZem32HAR6CbrHOHyAChkATvoJmI9gcm8ka9u
Ai+FEgknPdv+nlt7eortNACJmmF6zedzC5YqkzOmLuaxaMnTfNnhT4jPQEmj/Kbo8NECJuyQA2El
9iWwPZAPuqdf0sRWVX9Wr+CsxLDEeS7xE4EOv4CBvlacdOBr/o856yJC2qRTJKjU5mHO+ZVzly7A
dLZHxPAaHdQ4yjpxY8MAMfMlJd5LV6KDRuQ0vehgx9qsMS+zeQPZ1XDw4pc6nZwVKj4agWyCxfo2
6FMkvyLP+Xqppe3FeNz9r8TRzCh2RvPeON3Y/upO929PbN+SpWqw4SxHfMVfXCIcQlXpycdPtCGm
6foQSrLj3cx4i35kd95EGDcW5Ujrk9AC1MXwJwBK7xc6XzXxZuucdqtK7unRt/uwC2fWeQwUoJ2p
Fy7jhF6lvsT54JFDlKYuwh+YRfzM4YE4Y9zOtPg7o82fPl9tmmuetF+hf+nZPS5n2mC5gvm5H0Y0
3y/5WLRLWeefxsg/RiLoSUK29138N/mQVYcUSKbP7HzvF8CL46CkQy97Pk3941wv+TTBickHyj2+
5L8tuk1Ez4u85d9x4UBIf+0ojIfZh0KDe0bue0mVPAw+B98C/hQ2LaXs/yRCzmRMDA2B1BjWaNav
5DVPpGAU8MGhl3WFtr58ATUsqLsd6ti9xm6sY7bN6rR5NwsWWO5jrBw3li6CIYu6ck50ZjcRUKuL
AGm7rOH9TCwl4TcOn2djwM/X2vCnlKf/kajLBojLSMBK3f2ZKs0dFSF0+TQ7aP9qZ4NbYy389dqD
uP8b0kyECHPTgD4biA1qAtFx+2Y8KrQBe+kSHQ6ZQZjvIdC7vlniYtUPZDw9EJlSoXhRuGNitMgv
rPYucnLuPQE03PeCv138KYWEFTr/7AeX7wcmOQpILcvB/i1LSH7ZItNwkj3A5vpEx6Fq8zAg0JnM
jSo2U/f/cbT/WGNeNPOzbo0cVYJytq1fz0OWe0gjd6drkB1J9c3h8+5uLHZdfjew7Af+Y358BrgC
umhMr7Jg5nO9hYvj8Nrh6+djgjs3GliYQBiFvlm1y5SpACG0t9UAeGCu0ZLmvT7w0ma5fhSCbK+J
Hby2fZQxxdiLhXChKhmxYEaDSxumGFTbmjDGVKdoArBrb/adjOJzzxrOs241/cyKYz6vLQ+gL980
Vq28pSQkPNYErlDj/K8swniG22r2lMSvMq1z5d1Ee76BZdPR0Sen4a2Sya5GCk4T/8jWYXLSRAN8
MhBqebqs+gwH6hcFsMfy4n3wWCu2JK8I7I4fLbt8M/OKfkytIJYCC4nLgH6rRt6jQtTn8W3cqCou
HD2maM6fTOyUddf4bBBmAEDrkbCZqlEoH4ln3RcH5vaJFMbPRqgv0boY8hl8lOTThtHkRss7zWaP
0LAeKNg13qRoNSV+8nvxRCvjcX1QmTU54PrDiJape7o9oIZsmFNsXqpAnKVpTwNwJeVBTsyPYMlh
1Gc+w0wQD8Wms35IVyxi82x+lv2XDsi7OxU9as4rSAQyTZnxmSY4LomSQrgiSxk4PBJl/3U6+Ak4
kMiDxXs2/gCJUB+0dqjQvXU7VIB9kDStrTRfHD9ql04ES140QU4l2HBZRI4bULrQRHLS9rxkmlR8
z9Zj0T1gl0BNwgY8ckEwzbN9w/CwcmEhbMbjq1F0T1DG513kABk8/w6WfT/7eJADoynJHxJ7uOsI
Set5aNwK6dcuW/TdwWpViZFFSinknx/dsYwKjrn9Ysn1ayMGw0/ojCt8U9PyedX5+sBw7eNYBLjT
GFx/cvhvoel1v6wJjDMUA4pmQGItuhQ+OdGtkMITCwprMR4VXXAwi/v+0zi3yhwHyI3bccYhMJji
wHccPpb0dtRlsUC8QakpwOgj6WChxXlVTfnam55YI++2HjLu1ATJsK1GjMlHV/SyZdQ6miJgboSR
tRHgCvdclqbkFq8JK6s4bXm75MZrJWFgiNDpX576ADiQYXmJ+QlfW+ZsBgl7tjRiTKF/k3Qm3fIT
mkwyJqHZk9QvxH8c/w7KerN4zgoRVDOi/YOWIOI3yw1Rul7qZ70PsUqbbu9bgjW77wUdMwtjuwyQ
rlZwuFb4Y7U8wAt5SQUcuBCk87Ek7ODecsel+FMOUR0u7vMIG6zCxNOMizs0+0SSFmb1kPhtKkn3
Q0eAIhsbXuLZFLFOoarNKNRNpUKYcV4cZwi1laXClyTiKnIRESJanxZbJjjZXsbFOLpawSC14a8d
NbOIE4j9a8wbgSJJWO5tNMVNVqaoME9ZaXMecsQ1isx/zlGRASHEgoJwgzyY2ubEQhIM+1Vr6dFq
+sVR+h47k0gvZWA3Ddh5s7iHm0/vWmuFUoolJlzSCiGiItiF0+8vCFeb9xobT7baFQn6HjpcZM+s
Vl7b3IUGekHqxVcsempMp/wuZE2SWVsIqXl/f8YJ1ifl1EOBRfxoO0DNdZZQxbcdb11vROa+PtH/
p0QEOqVImfRaXqhmGwaWNBNYGbv0sTU9PABnstsnzqUFJFmDl7sl26BVY2yId7zWm9nZk7Pd4goL
Dg05WPCpK7oAxRNtjBpkHxlC3p05QvceY/WPnC+xdU58KZU2bVd7A+TWDd2FG1Dl9qvVeA1hRtxZ
1AD2CN9gZg2IXbsnw86YL0OFJHqkaVvy26LVcmGPg2jcoap3EoKJpVYEa527HWj7/H3VyCxAsSsm
pusdHahUOyr9Zt5ZSjaZKA5WRe0KchNk54KDcYXkptB50IWr6i6bNIpEe8Kx1ksGIVHRHa4feE2n
cyIcqWn6mgaJbrNVYibjBoNmpDzlPnUsLdm9NGetAc3XbxYnVroBV69B7yP4WS0r6G2fTaOyj89t
0g5/eKBUPcw+wdujyGWXOeHBS+21WUaI+/YdMoeBJ+ZYNROXTXHxcTIDkjKpjwjNTQ7DFDnGvrMh
VueHLFWuTNIvS4FUaW3YK3WiiGJHDB4ETCu89nUL72SkpBQ2HUAjb9wBIDajM4CmWaYabfc4rxsd
OCSOFgt6GpW8IDLjXrqsvfR2ykhQLURONPWAgGtjiRZ8TrCfkrJQXllasC6Y5hLa8stUDU5/6FUq
N0REeyTU4SXdvloEq0zcgXmQa5+WNNyP0VnkzmMeYAkGnRkIzqlkhhZL3fgtUVXGpYmozdJRfMUl
S2vqEFNd811b1ss0K/YPZujRzBKl1UNhdLEXq1EGVvjy9+rm2pkvBoBhzo3iqVhuSDT6Z9QYYvLR
uOnneYpjU9DSnOZgmWDYdlRO0dUxgrTvsQsqU1SWGt5NnQBomcY/oJV8xRB5s/CZuqaCds1zRvdB
ggCFDwnqi5OXPvmc4ENkcnajYioaCsaoqZ7vqadKApp85lZJdarFppy4PEW5pZUzq+B02j1nt46y
Pn0KZ90YQVd5O+Mut7X+ljbxCQD9hfFEim5W5XuX+Pp6f4WBe/xTtFDJyoKmN4KMnpMhhQ7ibhOg
n4bJ8GoVvyZAGGXNUH1/ZGm9UjZQcb0RmnDs2f0PpvkXHcKIAPkfo9Jfg8CSzJ6JCBGHMA/y2nMA
tmcC9yBzWT3nHkPserAoltsQvcHzBI3BB5N5ozzXXjaN2rfG8yQhozuoe5Z0qmx/o82eX1Y0dMul
NG6uqt7OvGQD+RvoLncAqr9r6XRGni8YOv8pOIwLZPTbewnqoSkOh5pXoGcQDGYlyHxQyPk54BVL
Ybq45JEpLXva8u/zelwUwIEv9vztsgbRJ5t8sHU8GJF0VJSOF+KgEmQXz+Dek0xV0P6JnSRlGfvo
Qx6sxAszY+2ciZc922lqoDHThY9S/RcaaU5X5Yfw55o8jb4/MkdsLC8rH6jqlcMrdzogegJX3RYC
gpQ3TRGtqnQuSq6GEaWfX9j3jg01ALjmM9KVPzweDER2BK4N818hmiykZ5OCP4CMNEnNcCQbMw+8
L3BfVqszGGyPrtiKU0RWBl0xO85eZVGeumgbwHeo1swczCopsFx6qfaHNF9f+ihBROX/zn09Hs4z
fUJTyooySHlhjSBpHvhENx8UHHYFCCAvz7GQg5j+INaNs493KOcx12enSYIo2gDMVWB+4LUvOEtA
4FeCfFi3/8klPzai8fSUSva0E8E0CmgcyUmuClfvP1YXAVZZRn2wCqMgcmfnXwDEEhG7Bqdgq4Zy
fIhKV57JtJkIKUnXEw5yhzpTvWl8I/3L/t0GmAIWq6zl61g+Qh400+lGZq+7xyxSvqQWDtDL5mfV
3UUrapF+MK7dgfgNE+bLprWwPFABwYnB/FsWPuufwmPiz1uoZOhNOJNbwI12e1cIhX+KX1rmgueJ
RucGTD2sWU2nkB9c33ev+8sW+nZDcjutKJknHanIqkS8KLREo1WsbTgZFNrg/Dh9mY/32088Rt9s
xp2nM0Uu5WqA3Z8z8I61spV5mrD870Q03zD0l5ytAj9tDjjnH5DI6nyWYgwsYz6hnkclR0nlwBkA
MalFOfttBvuoehxUe64vrNJ3GkPG5s1Z0NM/EoHUndrOOXSgl3BtqFjN8g4kHDLThmp79sbnHAMA
siN/i0t7AfsoWsTY0agHkzzuc7rjK8/uCXuFxI2JoODMhO+759v+D90uIQTqyaHkMUzpw/TtGxUF
FhHFxLC27RhC6T0voxQIRZvELJke2UG7K8N6ZaSB9sBx4dVrw0xrRebu+ZFVX2YXWPeMbFTFyg31
kAxY1OueB+mAKqLA2FWcdCgEI8FE1/ZTeefAIZ+uEdhrRg9BAtWoPmv4VEnje9b56DbVXWm8qJB8
bpFzucqX3gtbKdwyK1EvmHeSB4+c7U8jvWVCVgnAJa6ValSu2yVouxteT0IyNa02lbKlJLaEUNIQ
KC1lb0MJgi6C4fWjzvavourgrBxHWQBNJqBfloXMud02A7g8AF73efGkjKtbwndwoJZlTIHGEu8o
GX+HeMBJm4pQYmQ3uvDPIoQ4aeG74tZSnz/XmSBl/F+PG1z3GvcjPdS0EG3njdMgkVIED3lC3Y7Q
GA/1W/06VepKVcn9+pUR0SBrcc7csQyX/wdouakGzmYUHRB52PvCbrbtfqY+VmPk/oInbXFhrXWn
l8EKe/SJa7RFpMaLE0LGe8zbXbT/hNO0NxKOsxOBnXG4r0CF0GglDQllAWKSJ5gj5jBgFuzX/8bi
iH9LCHyIoydQKBlfvcrbeo6uBZIbwIR2+qYPY13x/g54vNYGMYU5PTDd0QhnkI42hSv0/eu3oUai
CQ8JiXlaa+Y1dItrupgsZ0S7vARJI4pVI6EDHRK27lHuiJBI6WSVuHi0uE195tDx5+9xr9PikbzQ
HhozKdCzxO1jEj2q+a+xCoQq54bOMLmpHxkLKY4PCyUFHIcBRd6eNPWgXL+/6LOvEG/fzlPsPJ5L
11RJMrB6JC2Myq8iwxVRCiC8DNibNmePZp2cbMemhdZpBBJqkKm47lHO8CfRkTyvbWK9zjJG/8Tl
B7g2xjrq8S2Od7V/f1wyQwpX5edoG6zEhPgGOp9A+drvt25h4VXRBoDnlPRpU14FpN02LAF0tG2x
UXE8UQ9+NZfFZj3kpA0OBKL7Ty1S0aChAKhy54jkkAHodb73nezxaCTkPOG3Q86+pPhKplbQRojr
PkPKa60enlvyj+VUAvLRAkbUhXixJV3nnkIpdWwFVNwGsxlj2BoVmqnX0mW3CAC4u5FBGLMbsKEP
U5pq3b2/BK8yYYxpzXn5/HJpcfuYkmRwI2HEWX6VLmAOWaDjf2c+pDb52YD7HFAYPRbPuFnRXBvo
gXWAG0NRq+7ule5tYkkrz9o35rYc7wBrvEzp+UhioF8lvsKBGKnew5Ikdre16gBNeUZs7dYCnVxF
Es2i308710BJ8AOytkxCis/y6HZHQHqKCJxK/3+lw9zEEybdn9/RpswnDXzdq0lzl7clPJ6iAS3f
Gzg3ZtSTl53rYlVeeeHPGKNxQ0aMJh3NxxKrVNECjhZGTqoa0l7FYRvQSiTZNfvJYm7botpuilYK
zGbvUso49x55EOrEvB7QzNZCcpQlJUHs/LLSLN0cvI+e7UH/ncdfpXMhYsbnnG5AbbWrTnMSNuyv
SseINLikqtC6MYCkXp+4oql46MrZ2GdlPPkBaE3UG8XKKQS1duFMRnmKDln1Cg1wZfp4dL8ViyNV
SSx7mxRy5q1WWXKeK2HznUJZ/fDCotDJ2cobLKcmEz4Wm77m0R75QZGovyv21bd7hwcfGsEcljxU
rZ7fMHQrXrEwm1Jfp5yawel4zsbWMo/iybygAP3U7irLziHTsE0b6kRb/6Sc03eHmnb1rOEvgTdR
1h77E5OBHraER2VT0fz2OdZ7sMwaS1Pf2tlm4Zy4dsz39LiA0iMImbxJMGwHno/HIZmIL4u4pTCJ
acXLrRum0//3a4I5XWpQtfhXelctT18eLjd8Dp6bbRFjUwq9f+9KO615qg/43WeOUitLNRrBqYVI
0T4b4tdeVKrSfFuUFU9l4kg2hqQjugzZebDM+q2Jcf6nVjrwPWvnCoEFkxCNlCCO4aao7s5fXNvj
/6lW9MaOkbwipWBT5eFgHr5N2WhI7W5/jk4El1IgdYu1GkKQZWnY34+8lw1x0sjcSUed8pHxHpBu
pmQK/Htggv0SHvwrRxFQNw8wgG7G5dSI/qzZC2/eH22bmkRw9pH7iOSIAmPk2GTBaXyVwJ0QVGaB
rTL3SBMUvg4bOCrSU6T2mFVCY7he6RpW7jx/a8ANxX3F9OVf44Qf5awFfUGBLAfbEnKdhir+p3ws
zfCAMyJdyNtPY75l8kanwJ/wAgf2+s+16HzGo05Q15jsQ/XEpoBdSQF2hyXZLvMaF8g9/pFttLrW
IsQPTfd1eVuXidE/V7NKKegl3iOKVXDGouh0+bWQbo+NiMKJQ8153PRA2aMkC5DvMrOHgR+1pgP4
1zImnWoZQOJqELoHYuTiH1rZAuyuOVXJzQzicsbwrtLOdH0gAqK33oFr2859Suh4zcxm78t2yluS
gBJofeqYQkItvQ80Gbk8Fo6xJ4GEY4I7TT2bXlNTtubDrF7TfgnOBwJxO4KLeNN2JchnXRD4MmdI
25gfYv8OhtbQz2Ws08M9ybmT+gGdWbmHiwMxVnmwOkLJc+N4YJuDP3QK8Cj/xLJiqmx6/VE7ykKd
NAjpLVRMLjw8quUtX+7H2TaeitKkyzYiZa/u5JcRbHSzoJP4WUFvhw9cVn+WKxeEea5xB47pq2e0
he44N21aqC3Vhh1QR8V+l3kBeMv+f9zkOnnzepkNNh2wMb5hCX2FueB5vJR1qSoIDC6fusufg82a
FbN0iC88HgGT6EyV3CIri+JMfT9RsSS9vSXe9FhplmjKkYidlH8qc2tsIm676Mci9JcNcIe0NgSL
MJ/q/rAVY5gLxcftZ9qnCrb3p870Ve8QEAagA8f1RveiSdfi5KQTi1fnDBVegp+CXAy0i7wZtJAC
Svy4x5ZhMPcordG8YcP2gIXzVZJswK+LgJO8fiouoekJvuTWvNbJTzjeLUkPU0I9khzzTVwvji/L
yVmm2fKP1Oz4rr65o5A3nkWwXvXMcM27TWvEwsaEjjZkx1Vfdnnvbem3NfGWK7WmObv+3zabrZgl
PI8XjfF9zH+jh5OxTxbW43lyiMoybnJ0RgKZE/qSpuBtqCmp+HAvaALC8ynUgO//NChyFk6ifAFy
8rKwhePJ2F/lFi8D/Ep0TBQsfaVtCMGY+a786QGuCvttW/RXlOiITiZQzq18sCuidcIKjfZUQb1/
Mu6rjorD3ZnyoJpFUpG1moRjJmIGSC+3QziHyUBPZRBIuj9msS8aO1uIMDJRYRm1eOJMxlFtiWCP
o0XXWZzYL2rTZCPwzXStEoZqg6PhUFBesnTsDWxmKc4cXp4QFXngBgEk3xZ5VgDcTtGBSIts43dB
5auR0RRAQ8/cnS5nbqYseqI/TqGTflLrrEbvYCG8bFXVO1G5lQ8IjvPTwN02bfhdQYGKm9YpgaD0
7zuRzCbcfwjcWS+O/8WR0H3DLk7g+kTCQkYWOKf6i0QqymLzW05IMkJHAGF+QgZX210RnBfA3olv
bp5H1txXhrMQowWu/4TADXARpK9jhox9tDSAdBPoufdznrLlIudpIT5ArRVKaGVPmgcWdxHPJPUi
jQCpg8373pOPzpkEgeuncehRTrPLCgxtqsyeztVD+sf4XtqGzBMPAxQ6rfOnU5xI8r8OT8tUxiRv
pjthWR7pFMMoSA6BmZRzw2rWyB1uBXpz32By4tLdEpNfQhPwb8vht6eysAY1NWCI6YDs58g6dW3T
YdJaURYisX5ETqS8jpFVH/E3JUa0ziAg4t5uRRzlo9Pbjw2w867QqqoJekjRWkxKKqLWkeWhUHGc
rc/B+araaiErd+A/4YIZxNZ9Ow6LAnaEIh9Sf+MyHwwQtnawZHsRpvufBFCSYXFoyU7b8A7WTs5+
JiRG7BbWqhYMVnQ/u22VHDn2HzCWn+24fUx+yyefLHRG23J3fMpaUpsTWNowvC3wY+fBuXfP01vt
cd0PyD1XMBBSgzjE+mGj36qQoNF3nCbpe1u48CJvZuHTZBbBdVNgPCbMS7CQWUa93mgQVckUKkxA
PCg0gWWjSjd48fHHwh5eWM8lK0nmZw7bO3Mv8hiQ9l6arAffuOwx+HKjcQeROAXwNSGJTGI5+dN6
CGOAhDHwDQ6cs6a8kHlXoaWO/mQCG8V+X5s08zMfl/Xzief9ZyiW9irF0aawYhAja4f4oSNIKXZq
lulesXXjBWdiwcW3aYvEj837a89qGm9NfOT4NWGx1bLheK5NqxWBBWCLKq58IAhqwSKW5V/hYR4O
yVXx2CSvK/3nOuo4TuD8p2Q2osIAkJ0IOZ3a2/LovUlpse2ZrSTs/0wekYKMtyMdnIkjBn36n78+
p16mHW0DCrYCmffHHCrooWQT2HOM333D2gYCXQ9P/fjrFnykAhmfd36AD3d1yI4605oly8ifQ1Xf
4qxNIF5HpiW7OLuOX4hsvJxLXGiyf8Rykh75UyXLx5KxiuzAff4638FU7Vgx5Xgu7hYkBYoG5+og
1FH+nEN5J/YVvf0ruozOz8zfeb9qoVQosiFbkXHlx4O8zyCfC/AMB+5p8UtUwQZG96p6FAHdndkW
+wiXsvMPjoILy00R4BawxkVzszDBuaoLQoSzEQR+hPgSg6AzwbbfaH+IDVbVl82JbNoooEPYlQob
FPBbzmvjY7wGOZtF8bIcPRkmfoPW0nzlRk+IjuERtLFOxeRaSTKAJQOHW/iTmYQcH2eFRkQCHbso
rFWYA204NyKfTBlJPSCIJe9q39yyQXKus+pkz5/9ptHJs60gaLuWVI1R8BChSeuyEDj8v/FBWZys
N1mPyqjMyq9Cka+vDrE+eQRz0uRcSgwA0NsifyDIwjxr28QBg8vfFYi4IchQvXthuBV2xNGdyJss
2kgQnrJGsAGVqoud/Ro4VV2JBZeMJFkoqNxC29HZnhceKzdILZnB3CBM4/927VNN7v92zfQkpvUv
NdlQ+MuPGYIYn2WsrKcN1Ni8sP1H0HQoJZJ7hGcj2nt4Cse6Gh6krtGrX94IFXmfxq5vrM0L8hIw
8lw3oYPFM/UtBQJdXUPPtdePeOot7f7nqwwsO6stfVqtB/tm7GuDtHiVimYbuWg1OS9yeblJKpga
V3230vswOR4imvxPCNAbor3Ob66zJyDWsRptJTHqpFCE0WD0bMrKgBfqguWPHKTj/UOkaZ34OAKy
297n/l+pNNBClEhzEcMKI9FPE3aKDHtCXh81YfWfnNX/D0Xtc7cmznP42TesNdg9MoJoNQSiazC0
NPwOrN6RtgWE53H3F2Y0DsVolswruj25BKRi9Wqg5x519XquKtQXOcywjZ1FePi9WDBw+X6SJS9B
Cczvknae9fBsWGsxlUShRkKoGt9NuMukbZp99s745Od9d6A/2BPomJyTxKCkFyRjLhGGRoKKpIXM
swWB1HiYLT51GEi8LjaPNol3oY9GjN/ugL0nAUtAT9c/LEFKKJyb3MHSfMrst2UuNj8mIRog0s1v
5whXRcPGyiCSSD4fgLSKuZxcvCbAzPZ5063smNw2xKnpJP1GzM2PQk3Dux07ILvzvQHAHf4tbqHw
lsHcv/wAxulg+9hGfO5r1iRsgQU2sy+pVkpbogX27ORnBdwFkFGr9EPwrkU6h87b1nsccUGyqRdo
gHsyHLlFRVKRZEO8/Z6LWl9AH0Ab6OXRT1bIk/1+7fx2eLVxLLZxyZGRjlmyAdizqr56dEaUJpGa
URKCJb8R5a9OLwNFxp8ApkDMbnWKKbJnL3+uK1uBNFsOmt0t15Ad96WogZRR6XpBbDddWD4yW2rW
e4u7GeJu/hUXzATiM/g9hY+q2NYVsscW4bv5CEWZLDjzrYNas/eF0DTQYrXZnDdvhZSzqaFhsC79
4T278RefeWmHpEADvLWguwnLEypMGHnFzEPhWUWl4urijhpJCGrXPeEqlN8MdSF4LjUhtVqNw8Wq
MNdntTqLURQdq4t0JNF7ufZPpP6b/8sTcN1UrmEIXmvslEJVRXJ8Cvp9L8pEjn7PfY6MJqgqDZYy
WLHky/lH8kfXYj08Xa8BArJH/tWrtzx1hV3Hi2VWe4vU0gCh2JfWOgFPo8Yq2EYXfVxGaMR69WxE
agcwVQtwWBOBa1wJ2EceeB+lN0sVhzwzapKWjoIvoUGLibekyUzNgPZaLrdg/ROBA6xSTqBvDKfg
hzQ1BKLi946B2j1Q7iTEzUO4ZuoCXOeJJVVqXJZpDJxamoLDZ4DmVSsaOwH5xGceT86yMkm3oMaV
Eu9VFFrhEbPs7plrl4yaZBxkhAdYJFAHGO2gR13dYv/6TmD7Y5c/rBIgi7en2AlE4Y4EzDzZ4OfY
TL+Qj8PKZuNN6ma8NgBe6Wk/sKFBA+xQSbbW1+UlCC29l3vr84hNTkirPbi4QA6182xJYHCXz2dF
ZXTQIe+ICoiz3CZedd5dkMxAuyxyza03kjpIxm5Lw0f6fs8VlZi4xNOmhexVIGtp3TNk40nbH8L8
X2aEXFTlP2Fz8jOXSW8kz95ttA8+Ed6Ynpd/aRrN9lA0hBOhyCi5iOY4eNyhZ809YP/3N9JDHXPT
yThWfWn8lGCS9glWhzmSk2j0nkB65CnP9HKJ0q28FPPQ7q6iUsw3Dfp8k/fpO/SqwOHaLJkCL7UW
9Wmds7jqGN7FTCycgYdnztA5jD/nXCOyoaZMeLq8zL8oP2NusPFINhqV3q4BAUN7lAILLd6gj6//
TV8B2hRiyqE7REy6ssTpL6cgbHbO8cgyXH6Q3J7WzE48Tzs6AYKrlIWwtWb5hejSTW12+0CrmA9q
hy5T73UFAS/FXjbvybQeMrUNeDpmHxjG10yffkUUXNL/GRoE5R2uIzfoAekEksU3inUyrFN4qV9M
OneE3CD4/bpU820DPWIOZ7Wa+TvYPVleh6AlWKCh21SIEZXXbuKIWqTpXiCffQVOSClVjAZSFQrg
vkI+F2KamY4cnMz31aMQiwI3sn1VhQLnehBXDY9XAzX2ZcChi2MTBCpLQGYUOcCqDgxkaYXBTpOf
q5iaH/VuNxah8u1uia7OoTIJEH5xixZneXPVhRtV1OUlMyIRnyf+qxlS4ecfGMP6dRUwjMpU1mke
iWuVO2fUJt+7tVH6kcbugBb1VTwuDnSxdaLo+1BMinilP4m92BZihRc5ZW7I2GpJYvN/EvsT1JuL
2usd8SpZmlVqLnzJybNj9DgxhCMMHC0I4zUnnxIdKI3u4VQurKrGNSrpQ3G3INK0ecUzomQXglap
zIirHsuEH/Sv4i1Mux1kIUdFKXyh5ISfQNs4zILgvF0lQ2xZ2AVG+XM9matS3zhFDkjuE+VcHc+t
JnHFbvZ4mnShSaXasF2VA4fgWQSUJW5AnmHAplsvpNYUJpm/EFFn1jUoL/84xFGxuuUI2PoCeX0G
Uc8p3Dm8kgsXGH8gP55kIv5cvnMHiq0crVTKUoW5ZwCRiRLJfPUfNovt2HgfW+RrkLajan26rBKH
XdLIihOlBo02R40Fmby6bsHKM/i///c+3yO3ChChkHbjTBISWSHJeGWyI8hfQWpWpbhnocef/L6H
VVhLxLgWb2MziBNOGB7csqkiumbC8fOi/ySLEHr2/QF8MfTSnDocf6PxhHW+SHDVoR/c03W3jjgR
B/3/gWNAm/OzIpgQLHptH4zgCCWqSTFUTBL3Py7TDEmskwfHSYG8GnanIknT0qWGIryFzkU11PPJ
67V9JmmpWgjhfxVOvTAFzE3HJY5nDJ5qfWgyKcCoDK/tCqLKKOtcRKH9cMmZZQKJOrX+58TELNm7
W9mRG76s4xryIG3E0x9jofJ6Jvnc/5NpvRWMAQ4DMBSPABTbBfqW6/DfJ6M8EnD7gHKgoxrFjHCD
k+ZE82h5nTdloVKA3V9XFYSOGHkOdf+LFTYHwZcpDhnNoCLvVfZCjfyQbSHxSOQPZYCtKp7yZ2Tg
rghWsO57g+CT7L2sJXauvf+7dSSpSolEY9susoV7MqKYbRls6E353DSCdwdJmgGLvoS9sMXqKnFW
cOV5aPUEBaI2WQYK/6BexqAQEAAM5vv0QD/+bBVZM0Iq0kepJZhHUF/TE/LIoBZ+1nAuUikdsQdY
Fcezu8zwshq51T8FWOAMbfgXahRkvWJpYpIp/bY/j+cssFNtgeeIk9x2ihI7hZBPji475VvQvXTy
VwlMB/UxK8eHG5Y4V90BNIDbd6MBOfCdCBl0uJnQlnsYZySkgjHMy5aefLgsRgkLz+me5Z6EzS6z
v07loakeVDyo53c6CaWPvV/LqosWBgPXqmV+YLPO+r+hcYgU2YhwEOlDpJQ6r7iW7mSIMH0rIirW
ryTrvvjD0AJjch5c/8XGxVl5h39RTWuL7pW3aU6Cs7k1Ji3iwxab++jE32uByzBC7MxSZuCFoZIr
1zmYOKOh/MVxTiacpmpTfUmuOUk7hHO0KckK6TB6ESmP7srECdrhJx5dx6RGuk4O4Rc5Le11LEKk
XFxLTydGey3pdmPpVpId/BAVzKfqaEr++k0SDc1H42CCfKieb92oCB6XudVqagUhPz/8ZKLm9Bsi
LRJqlV5nhNxBOGvMwMH6vImq6o70ror8x2VlJGEw+GEVIAHfz+jXt+MkV0qH14/37Nv7m5EdwfCG
vun0TDBqJit/sEKb963IbNqE5clupts7RhIQwWL3EkGljJvGmI0vdVaVezRbblDaDuJL5/cP9YkA
sYrI9qu4eDUp8Br5WO6gWK5c3kgXsp5/llWyoIB49aqNhj2kTHXFJk+6fi9XQlk6v9YxFA3DxsOO
51Lbi2JOCajBkcOnAY0Pgq+7eOTttopTJzCr3vHu93O8ryktdYlhd9+xm0wmVBfbw/dyanZ8TvZw
iMg0eYemOtzrxV4L0N+NOdJEt5w1vvu7Os7klYm68s8HFz/RXYeAHfr/r7q9hJvOt1eM8OWAMS8o
MstiE6crx+R2CRlXOv7sTYocLEM3UZXpzf8Qe/stnCZEj2kRin5pzMxBtPuBp/5mzVkhPkEdu80R
SreVA3WCjpnCrwkoD1SU8hVVU33FFhT+AR+ARSokNk4GKmpMPWrdQbY6B2J9X1jNyEyVT0nBesEE
oxPpnZCv7EOOw74oJOErzaCPaK6/k3aML6tDe/pSzOKRgwqz9/FNdCZnhsQS0n3RIGo9nJUCGYxj
zJzi4/ysnawBW7oPlt335fn/SLU3v5KX8I5J65ul8uWMJAig0NrZ652LFUpdsHw5fcdcU9Urcsbx
+mzF/LbzZCB7kIQCU1ev884BTygVbx26Vno39GRRw9cXRXU4UyBXikfsUsd0gdM9cYk1hOWjaZAi
QwI+RiCARuIUmAJV3/0vE1BHSJFXGBGniLKdkYDQaeNhRCtrzrTikqmNV8nG5i/O6elIThdEIXPn
9rPaNKyPBHxuKNlclyy+SxMkRBmrUyD8yRMBkFJR2stD2E9g19a2BB8im2DJA7CKAGjnMAmbs1k1
abMd1dKv//y/3HNqJ2cZTKH45p+932CUYq3Fx4tuoA8A9THq0RCpPGzFVBbuqlGUejSfky3c2dDF
jWGFPWxgEdhFADUKro0SOYZyvGDQTRBbcsoNRPwaGXfoBQdYjC3497EVRigqxaOwHg0kHlwN8/Uo
oMjj4Vb03V96ER1++0y67PClAoUbTlW7SMdOk23tzWyuK3NgoeyOgOMlPRpMPKjUxMUa65KQs1C/
OzNrwG1UWGp6Aldj4gB8xXGg7Aa+LvK4gHUmNeClvgsyt62facSYBlACH6VpswQyCcsbB+Ox/g2V
bC6b8cIW+tT61IYtmoAfuLcZ6CZguQNVVkLFjhcJQCFJWMjWZXNwIvNmmZhlZ6sHini+K8amN2eK
xWgpbaH22vQo+ExNDF77EIl1UuvnHqEwL7l7jrCI8IstLfqcJGjbriMiS+Dag07Y2Abthy4xaMP7
3c96kzLpndrLjRLJ6cuqVUm1g7JsezsTNvqGTJZlUDpmLeTpNT54S5VFC1R0iRwa8F/EegPdSCbW
+s/M8Onq+QVo1DSgquQ+7fe9Mqdq5zX9G+3uHHxjVTrdBCGPqDybuqr+bEu9N7INw0JuWKUBli8z
uPNb6yTBQh7/Npp5cXCuPdU3LcGNBpAhqKE54voZFad8vsLhAIkAsigPNijHcZEOT7hYpiNDtpT0
YebhM1Z7ar5ymYrxV9Q6kaMLL/f3ffR3ubvmoYv4zWjzQMuEkW9Yza8kUhOnxILOys4/kLKnoCXx
P+azHlkLcgPbCH4ohNPL7ZHztAD5tn7xEkQqkF923X9SOO3RBhOM5pTRQAYevt1qZw1nkImFTuDy
NHACEG+uEnb3OIZvFAWSx2VO3D0iRYfV2abwO44B2mNCVkuqhp3wylZB2rzi3jy4+BFZrXDB33q/
xzm8bk1xXHA74yMSB+FXXsWNjCjf0JdkPmx8Vpf7tHsD2Iwy+6ua3Ccq/kmkPkymjudk4hGB2V8o
jk15P+gue4px7iT0dlw4Qpi0IZErEbh6nXmS9ugvbZchLNPkTqYXyb+XKRr9jO99OSPSTKDEum8a
QUqvl/Xc8LsL480u+Um9EgecPo99Frjah7IDHeeTislhpZLvnStPOq9pw76lj5NjLM5G82qk3ZS6
S1LKEXc57bNtvnUjEuBTUzKheF24aLvwpAakyw4C4Hm8ldVpPsyf06n6Aq4DGgvx9KpwqR1KdeWn
GnRnvkKIvku61k5Rem3nXvcLrB4Jj6++3W/U+mg6s1iHgN+eepSk0oBGVmmR/0k/cA497VpHEA5q
lWvFB2iHvuUpGaowcmcrcnYWUvAk9rQaSQODFb3/AWaRawg4IOt7/r1uOCNLSYDSoRvWDerIVXpk
9ycOIiK4f4J00noc0/VqlLvP0fP6UApC4EnDl151vN4og4NE3pbxQZ7Ie04KbFJS0USqI8hjQnJp
9nsD76SGszQ90QSBQcvRtBniyB9ZP6WaScs9XchKC0JozqS61/9CAa5mBh9tdFTf1yNcyXLsZUdk
IpkDkvycI2POyUfB5ES/2XRtOuEUfeEjLMczO5tiq73gJKxKYWslESa/keMDyuYMyeoD3+5UvfFN
mBNsgFpjWne4uBDwyV811D3F3Ln2Y7hLmPMoAdWyuzYKcLzxSuwIWXew2AyuetzdQ6fvbrLifbV7
0uah1aBH6yjK0EEJuhcXhK01Y0XrSTfdCcN0maBbx1kO5l4GEElBAxQC+Nl+RvA0A0rreD9zcJEI
B9QyH5oX5o1UF66HF+4aWMhEttX59Fg117dTXD8lTgrpEyUdKKwgjRDgO9KZg5lFtj4t/FNV2/QO
53gBJg65sKP9Y8nVwtfYdxGtQj9t0esZ/dcetOr+yoOsPFw+LrznZx8MUREQR+ARvkju8b+/QHzz
QrTWY1ZywxP7mxP/FtPVh7T0ihfB4WUClPptFe9Y4/A7J7fW03n1CHeGc1OlJWGrTusWeLY2v60g
yY55R47atpz/i33rqb6veik7tyI6pMhfms68lpK2q2KmCDpWx7OE61ZGkA1dy3F/BaLKRtZTHNIQ
/R/YGLdwWwBWV7SCzbLx2Nj7RjsTiXz5BUbt7jWAGue1EASVeGa2+Pxhhuta+tDiwUj2ef+qFWj8
oihpmfjRjwIVDlEAMNYD4rbtphkSULNYX9fathIrCYzjdL2qCtiXptODPZECRk/yscl2MJbkGi9u
lwoS2YJh7/KM3M0AZfp4JYoUTGKB3IAGtc37a5rfsUpL8tBV4FchNrEGO2yymDeF54OP2x8v3ZH+
0+60oRqBm4QgGJrkb3xSF3e74063azD5RY91azs1XLKzIp/2ZicoVOnxhlc41nYKyGUqvwbtftWw
nkHMqqcOx+fT4CPiZEtD9eShafW+tHIJKwOE5/J8qUBsBmrJwgS5xFp2BQboaqa6GwL5ce9bPsik
qxcG+BTVcEjyw82tObPS813i9qtu2dtexji7jEBiiZpAf+zQBGUc8WWzFw9jsu1EWxS6EKPBTbV/
RKUpFG91C9uVb+qOwdKPd3/zWjeAyBBDDqkabJgFWzwJNqfmMX4b2Zn5zeK8ZwKl7W3edfmxADay
udFLOqcZ3v9aXKOFYemrbW+/MSHG071BrHOSdZHb0rlJqseqxwWJ8Oqxg9VNaVp4dq/shG49OttZ
ps8VOSaDog0cUCqaVKvfUOK8ytkUchQiH0CTKJdlNuuoqTLywXE7kuuFIrIgg2+lbDed8FYRyC8v
bI87cCezesecha2wo/TtwuVEwu3dJtpm1+fNVewqsI59XjxiF+XJADFwdEq8uzwmRLe0MShAjyHg
MkQRJKANv8+XOdoJBTTTmzN7Zp805/qgS7+XSGKEk7cChm9E/1Cdrh6uWdl5m9dIq7rTeyEUfswF
l4ydLOMbzybfaKcPMrbzeOWf09Ee6qQsHfaY00rP3NRg08TsI+5bIzHYgSYPzEK7RlEfiQ0cyUTZ
mDwL6G+im+Dvt70d/k1SgWq1hJH861gVoSRxlm/6j9YpCXLn9tiSXeYT+XBlNYikwrsR1D91++7r
9bSLRd6r3NmuiJQxueQ4qh0/IVa8+R4lM6oogTBcqRPfVo5YZfbPpP/2XmaWoGQupus3T+fKd4Qk
C1Rmg/IRSksqVFiiVqjOvYvvYCdWS29cDVoKVXO7RiOdxnBeLkwlNBsZXSxAMbaBgKpri7/fAELp
xuqQuitGGM94G7xS6wi/zgBycu8RycMUjJGSO0FCJ6en4eiTYc9YtQgrAh50mGAznHCrXduLe7V/
YSOpqi7rl9zKOcabZEo19tGUqEm8VtHvi77sN31ICaWaTMTH+XwxLypzmxHbyYMvZUW3SjmsMfaJ
msDZ2ONeNY0g142XKCJM2YGN4X8KMwvwtQ+QOdXhp2Of/CPvfwM4oApTW5nOB5924Agsfy6ByIAb
e8bzubcEhM3wmAB/tGqvh6Usmadjg+1RwwJ1j1pQktdZlHTWR64AgDQwiAa54ua17oAmQUnlBGv3
DDji28JpsRn5/pZWiRboLyTcmLZDD+h3Kk+wJlGnSEqlj583OrxmZ/ZaP1d6gsCmOb5hmihcCwfh
qqC9rQFe//oaplrQ+3mOPHVEnGATE+N7994ULEBFrCWQrXudvp6R6szNyngCOkEAWZdIFVURqBAI
u3KMk0Nniqa0Tr5ayh630w7OVOvwfGxM3uDFmomy/yfzCGo9hq2onFPoovJdfZzafvoyMrU59I6B
jV/LKMYUICDpRMB1wQE4JXUoMLgnxYKJBYdXdU3WnPApjKiFF8lhF8/o9PWICHnB/8IOkjx8ypgR
XqOcjTAQdh0pwYVYnHaIjnsbVhZd4l48pR62leLMZuan3ZDZpH+UVdkkfFoH47Ati/joxQW8Oz3V
oANVa7LcUrRCdlHzo4BJT268i8+Zs/yXc/4hkQEfIacYcmgqTtunlkXMbBedOfZAoTIrCojxL1Ih
HvTHgk1DjrD9+2a0rdYXXfsCsHJ5FeblRRLdIR97stXDfeepCV+QcxhOwNXInV2UsDAkx4oROhjv
5L07pIASc3PmRE5JEdZohTj2dS9mcsRXy5XTJjDriz+VRfS9Aprdlsl2KRb8bsJ9vfCNtOV8/TDE
hl11U+e7KDEizds4U8Go4bKgQNF2VAUK/7bsw3V4pJcddtKJSfrH7P+N+Ll8IgDONpSbPOmXLPGD
+v96w1xHmLBe1367zdlUp4ktwHs5GlCeqpKXa3zakz9YMVXuSB/zXjdmGSo2uCVF8u3XTxPSjEPK
bKgyMvzFzwxlJqKG1gAjGq8oS1WsWC+KPwCYGjqZs8c2ImN5T3IUzLcCjW2WtstSvxKuX3ReVwAW
jGgoQEjb2jCMYdZwzO3rM5w94c3J+2mf797l7xJueDnAMwCaJUIWVyVLU46JzD9mImlrkkbdQ6R9
qVq0G9bnG/Ci1HNCkldOipHqHR5t2RRUZvSmyrxCWJ7Tt2pCAFLmzVCVp1cTwXmhE5rV0Zt2z1zl
kObBt8VGr0GMbX/6G5WKURBYd8bkzcOhMR+Q6zjZ9W+id3HrVjri4HViiBPv474e4amSGi8AbmN6
6KL6VmhcBx1vR9cchXSWX/7cPRva+9PBIcTpZ9hh+FbNFC5oVR7978xD/H+IyiRZPb/TJ8VKU/Jd
yguy07djAXqgukxEnz6Ek00Yj5uvlpg44zoefEsWWSaUHQgZqj0M5cHQuINM9+zOJ+gaYxXv4CpY
Q8YzCGPevkP5AC7GgsSmnApee47iD245xh0qxOgefA1RyW0OfWNjzEGQH7UaUdikAFa1k+BEbhLN
E/BNpVth99lSJT46qw84fbZbGdb2WlKtvw4X5I/H9MWGkpgibVGjDqXufGBsa2KDnBhtN0cVvBdN
HD2JXwAyABwt9yE0wgl2+VYnWw2KnkwSkzypX6wwEUCVi5yioHrrdZ43CQ3SoBi0An+I6NlBfk2J
VigB0vNwB7pK/zst1yNV0QIxeKRNjjfU1JO875NGKCSh9B67xbp5alOTTzjT595V/kwxXJ0V4/C3
IuZmoVi4GeajaLi3RD8GZ1oxzGzgRLcHhgpkaKdmNgFueJkllV0VaG+Ny5eNiidaMMiT5gjlyWAQ
+H8oVC5sSYPwHgxbMroytB53Z/xkXxHdrLAl1XczHWDZumueVQRJMT/R8gJsLvh/dJUxQ+z/OMb6
bax1lCKpTVZU04n0gwfV6wXeJ7sw77xtyUBbAHty15Mm690h/Xs406w/2++jbCSeR+5/7ClWMgfo
p5XSf6Lmu5t3MARdmYnc/hF5r80ktOsb0SiuP1WWalmy/bhLB9BV77vuY8fykFiU6qkm51N7Qo8Q
cugx23LF9BdsdPzDOK4GXKmF7+H3uID2dBfXVXanIQ7i2RmM7eWhD7WsyCFeDHTC2wxnvIO23CKc
bbeWnuDZ/mwWFd103AUbvfNd4IuYttQGcmYas5EgTW9PEu7Ywh9HJazoZLIU0enubvdGxPD4V/Wl
pDZ/rDiWUPTZbkM3FLD/e8n7h0PlR0vyjF3QZvONrtr163VpdDxzlMyc7m0svBgkJ9oFJkYRXlj4
Rg6ZLm6JeKt6Ejvjcjbug9dYEMnGR8W7c4zZIwu+2z96N3OR6AJn6/WvDhhzUt8LoZ5wug8EPCUP
JKELHRaPlW4hGtzXcJ7jgvcgITxBSdWno/QJ9Kbk6B6AcwUsVZ9mKW1nIHUTUI7/apF9mjZmy/G/
7SzeJ1xs9ICXd+XG3yEfmLExgHt8MytMNE8QqVGrJMjUB8lAigbf5qkXRYLlscCMEC7MIGSccAXG
himnXM/OX/1jmcjyA2Z9oYrbL3pzSShZdAN47OFsCl1GulmD4rz02jB9cJiP0/Cixu3YioE5e9ao
ya/hUMntRyrCDQuR/5bTv8JdqgYoe5mG2HLGkwBuc0pOlRqtIjEsnDHOWHj0Fh+DsmzBeG6NuZht
IQrCooLmTtS/+Hh+dQpjnBHYCvBWVb7sd4e7N0cNGFeDo4Vv3i47BDmgm/HPF1rgfX3/YO8+EgvJ
ZTXmG6OdN/N6U5DG3fAgS4frEFa6siDLXdyjeBNykfvsHP06pbrZfOak0CpccARR2YWbIlOybTLP
H1lxYjIm4fFiL5BI9eJZz9mVCv5wh6fxval1X4TqwDUOuUiCoMLjXFjXSD5L8obuiwSKBo9zCm6O
sHCG4bHLYPBTNOiGMNs67HngIBCahRAWJ4W5oHGyLwzynDQCJSjBjyuFK/6wnWDP+hWB7BmJDqzu
VZIl6tuUwlBfgzl6F4DrWe7UmoS6V0uUBZxEz0rI0EtF354nj1MpQIShx5C8IBJr3K5MrDRZ7SQp
LCcefPDa6jGVHle8b82MqavbK/6dmAKBTeJp/necoQHfjNgy4p4buu0VywpBrymnZqVsptM+LnaL
1UnpI79EHwyUKMMaDOStDLRwDBCK2tS/RWt2I9wUqrSHg+evMUOJj/QwBZUWrSzxOa044MsPhfsC
48PEgoRZld6zACohg6fDOydYnxAluR/zY85PDB8331Qb1YXA1RhSR64azbx3z8bHdMWI29gMJB4i
R8MqWDA5jx+zG/Yrm0qKBEKcvPWWZJTcZLCAtgFX/pViyuSpBtUdRLM8RAZF/tyHgpsG9M6BARYv
vZLwEVWFCDKGJxaxz/qFT7AhQsq1Zg80AYpmHX7vWbUmoiV3LLPJTyOcaImry+RhI6uLTAaIuUoe
AfLmvQZulDCgjqe29AYfpTSh4DWL/bZFmGtVB3pyxz62L6JoUqgcnb62PtKzd4N8joUqxGvRCtgy
w8mD61jZGUwcre59bcl8x+AVpTrchEEPt0W9eNzR2Gm8XWWyaon6NFkUp/KLo9f2l/Vd2f+VCYQ+
2qdIUt7tLlpoEPVZtYQJb4ZEOjQXR8gHbGjX328iVK0j+0Q+kxPBuzz54PGk64QlpPrAVgeyB8jQ
yyR5fZqmL/Bl5rl8U/QOkONT2IWKXFxpTY/BTpWhPt+7M45DCrs9oVYO9EWm8M/DgLTqBxK7umav
Vet99kJXunWxR17wD2s2y6CIAABJJ2x/hmTU6biDhhIjq373TF3cscjwTXQb3s+zO2fm1Fjc69nX
xROnVTtxFx/YXZIuxl/43RcvJr9I1FPYlOya4cu2X/12fkYsa4P0a/3qwZfApdKDG628qtG7JcOK
pwBfDyngSq2GgtHd1IGgEh0k7poXhnqHHZHEMvr1gu9eQosGFLnjJ6Fc1ykkI1zuKEcVGnb+VApf
rKztIMovsi4YHlZv8ZoeQwxUQ++RPzdDZ+CN7qNJPl0mDNlWBbfeV/40XakNTXW68XYY5zhielSz
7vXyP45PuLNrS7ebJ3UQvY7HVnGA7nKF8gL3O/lKvew8y0Ku63MbQ9W6/9chyiXwhkCYkdugDsgN
8nXQtoNXda1ei2Ydrt2XgJwcylE5OcSvY8TyvICrqYaDb0pJN0xe3TGNid7IJcCb7L+ZKGgR04ab
14g5FYpvVTfFHk/Cy5HTJnhgUHDPE77JfPS4xk8vHxLqMhLqEkcrtusosG/YddkUPzsmaaBk1xVk
MEJ+Hitjk8PkSJUMUuwh+VrHKcpkngLL369U/6bBOYqZAP2BwFtW2KCSXoaMJ7puNUbDHIO2uzNI
Yh14UCTPGtTvLKpyQBwpyg9HstnWqC5sVVz6kUx+fmC4v3KfjNKVG0pfe49yGFfoAGY8eGrSTXRR
Ulywd2ZY2J0Ph63IgzM+OMhWo422cQUfr0RmL2o6GJVdkR4kLhVkXCcx3le9+w6FmmegBhFFeIcP
6srAhpfIWqDQd/PM7abGoqmth1AzxZG6hGy4X3YdbxR9cDydudVx5KYrjy+6IhRu/UJqRY171fxR
sefFlLIhOCsWFCckzLTZU9Jt5ylm5HLrAm1GRFSzTy+gvCN1+ddYLutkF79ylXdYllMSHGN/aZ88
dxlgRozX6V7FfEuHrss6d41gcqI6zH5DlxNAQf+QF2JGC9LEqi3CBpBq8TzvS25SE3P64mVQS409
FBFxth4pQsrDxH86eqP8oLhf3AdOcwmolEODMYnVIpYnuU31PmtKEfLHO8muasvoyLsigqAivsf6
2i8vWdXucmuTBV22tQrVsEAU7Z4Hw/ZuFnM+QM4UgPiQSGqupo9hDypHqfVv+jZtBIPueU249tD/
nA5bUnncnPKUDYvEtCJ09R1IHVdMWuCnYYAUleGQPtiF8yAXUmGhOUpVivoZHKwdXFVcrHPg/6Gr
lUJVPMERvo7LNWnDLu1DLnvN0qTu6ToRO6NdNu9zKpL51CTGS8cdR9l0zIGHccEJK58j6lu+XcWH
8GBf1FEF4mFj9R2/THT1YDjZu4oFusxl1WGJg8Oq1f0B8Sta0fE2a9DFwvRYcEa0QSx6t7aVnfWN
4cEnixKVLt/wz/M9Grb2sUn9mQ5BegSp3cHB/nZ2l1PBDfNIOv4Za40USmj2hUHMDkR3tFISPtXm
zOU8ZuW7caSo71KEas6IPtjKUDhH4NtPbmXcTUzichpAkJTkCOKkieMRtTOUiq9ZcSFrm40oOspH
UO38sg+BCeb6HONq77QsOmIh34DcQ1fY7kuAgwGy3M7V4XuhnQtHQJ8wx2OkBqQhpnlXyEWd9df6
OuLyzQUEsyYUS/vSeN+kfDnE+5P2C3Kkky7sGZfC4L2eDowfv5pEIa5x1X8DcykgzIMzpDnkgFz7
YMdDttPpBiI6r8hghQ8fG7xsQrx/LTD88h1t7fEJM8tLdIWFoHhD/58h+zHusLOfdqj5ceV89xzu
DDwtO+duYi20kPQZ/qaDC5Oo690R2UKyjhun6QjhhGVt1ONhx2bmzIR/A92FZ2XOqwsEuywjsQ3u
JnXyDj6w6qOHIGPqzGUgHmNtFzwVNG7mpoRmoaGjdNvowXRtVmGF4/JP6fwxJVF2hR+2cuSGqhPQ
+4YmwUr7u7+G8hbjSJWBk/Gc2/qrjEPSeXHtBpYNHrHmXTL7KRjqmKLGUOfGO7UW4DrBJ61vBtJc
R5GrP6V1yDvVRgxjFdHlBlrNrjjwV+tw+JOorSfL37VlFoC5qx4id1gS2wv91haZQE2DZlF+5d2v
/XgY6p3zuwFqw99FxIQ7M5XCbUxt4OQ2uWdrQx3+eRvmPZbaq3rl5zTukkNyreV8+N51POd3cHkK
DhQuQYq02DyZaBx1vu1TGH6LClC1yQVORS2kexpPVlogu6R/AkJB7o1+jm1nvag32Gse9aIvCQgb
bH0Dst4/BSPlKNFfwgk4zpqu2fIWgt3armUgGqpbKAAgHTE3/Joobx7ZMuxHXPxV226qCgC595n6
5cyHwjMr/iB8LaaGOZ7TdxbIfZSdjqc6Dr8Rb1445i5Qwan7LpUXiafdIzOoS7l1ch+IC9ajfqz+
VkLMg1BWjtgOboIzCbu8ydqwO5lTbs8ufmfq8G0Tpl1DKq/Tpvt7GSrsty4wpOj4g+xPzD2vgr2o
kmwdfZLWJP6Frcl4cAf5FCJspcPrBBd4W6KBVGb4x++mA29sIuVdmof4OoJukeuzWFJX70Yppwhy
35XAhtJcFHmk7OvJxpXwjtId4KupuMdfcVVqcnZlPervoKL8L59cmGxq9tY9eo42kyJ0WLrZtV6r
ZApMX+vN8HGlAFPINCHfC6PrdDoFD/6EHkj5wbICWCgMUXl8ygXR9cJXKXbYTWeD9jIrraGXwZbz
7Z63nI1yDCU2viFXI4XlEwA3DVYb87powKiG0tY556l2cmlYFi2nFmo94058IBz6PbV05nRv31Fr
WgtEIlB6EOt9QYPfpSM4/djJ7sYf9H7XRCXmQQxnjWM4J7dZFENa+zrCGFopku/LKo6ex2alsPha
UKFI3wQ04V7wQ7omEn6GGGwocm1RcAoPgTMhbVqG2cVcg/Iqy+sQBnyhvmq5o1ixMb0ROlLmI4lG
8GhVpMMujHN+6D/8i8zCeurAoh6kFDSVOObaiGvgsx9opeYOhMwEP4xbhwaeGQPDeqYoy+U/bBcl
i8tU9Qkz0T0twvbByn5aJGJ73S7ZbuVY3cpLsUTqD7yuu2bt91qW0Oxowt5L+hPTNI9tjE2L2Stw
YDTDGHY+FLnd7l4YT+3kdRtLWKa4MQtZke2fU5bee9Y+mlYVVP2PvvSJRQpK2alC/8H2fol/jfvY
Jr3XC+8VqbDjUtpDLbwagIGxPdZ82q5Mshu3lyzbeqWwkJpmCQWssReiTZuvNEPJV8EI/KokkVl7
AV3W4Wm5eqNcjkVZJC1oYI4JnBuCPDlkm6jvi1wg030mI3jxvlfOMyYymAcVShjGFJ1zM76CC5Lb
YawEt8/VawoArvOec+uBJDyevL+p5OLqu5/L9nqeNriQP04ccVavcf2NsBpwOatYJCNQl11zd1Za
7TjmzriLDJRYtRlGj35KMuJp4Cn2pNv+Ku5FIvZ+FFWE2GGBE4yaqwGgbsiq3O95oiMBOdPCT+OD
jLe9HN65qdz+qHaROP+JjDNEdHka/OQGyeObRBqHjqQjLMKxq0Il+QqmQ47BbjVJRwuyksRfW1L0
BTyBTsDfmowPLj1YhHnjgSc/rN+4IY51MfuDOhmu+aH35cVFl+IuJXsEYKiwf6fQZxXFp/v4rK0g
jZuTKyrGtxDoCxcaHJ4cRnPefzuHcMSTyRFNNEs0U7ACzhG8McJ+G9u4cYD9JB8LXgYquJ/7KwAC
WJ40EYjCpuQVMWohFI25TWIUqwDKwud2ijDNs9P+CFfDPi5fXLJ7AjC5felU9oPulCV9SVxP9gnP
ExCSaxaTledvhos/13EfsKd3tlsBlMxXafY5J66w2L2oXIr/vQOu077enjilEcTCoje/UxHg90NH
PgWi+SQ40NN9Gv0aIxqCfS9+GbHHt3Balogf8uLVaOuBEYFQFViD6zdzOJ1I7JuKPVneANkj2aYk
iIovdWWP9ZiYGkKqU0bDXGnDs7xqZajG2u+/388224vI5p+fXU4zlQ5f5W3m31gztPQ4NAt+dli/
FAXdUNC4u0pEkzNbqeXgQPdaIhGdr4RQ4ejbjtI1FuoeFOoqL9aACwLr25l/4VpPkpmj+N9e+mDV
JrCLDZ7GadUM+fHZeufOdRZduE6ofTfPr1Pm1hCkYit105tojEo8iMSMA/OqWQQ5g0OeI2DruN9V
GqQSMrmi9T4IwIW8/joacKq+y93y6ROurTeMAw3qBctuTD7O1rfqIUEdBMmv8mdAzlARATRzwxRU
L/c8C95t6ckSRYirBoKGajTQFFwgKOrZktZEDJCmF1BhRd+eMhWTs3oIFrfpdEsi9PcxAUZtI/GZ
RbcJWQjT4Im8TLLCuw0EKDXEDB1ueqK4F6sGG2zRcMD/cWUajFq76cs3FUkyRtM7vzciNqKRZ65k
qKn7upWtA862HD1UFI3iWYklagm2iHCpSe5T77WFhfdP47vUk/cTbWsLN3/xac8LSqwClzd5N+jb
bKO9BdtoP0zbjNra3NDP3LmGr8FA779BXNZ2h5KfNSwMvp6H0Vv07xWw4A8pmSuxtiCkaXwE9R04
udQ8gH2Dlu5Y14wklQpGvyjF09ZmaJJivNCmtr9xUhwZYKi/bi5voMrOx9sZbUDPzwx7P37PBfRN
r9+cGMPGaJMyDHXYXiBwPami9FNV55J7MkE7LrfZAbug0VCu9uvPlcey+gkEZ9nwYXdHsJEondH6
/KwmXcj4e/59Oq0j3wsIBExbIsjrJanhrrWDmQ45+Rt36ZXYVmk49xNmD322/V0EXDi37m8l/AuY
SOFrrwA7vm0mJogaQlPJqRtc5Iz3e6xzn8jKcny70w1sPtr9fpqSDLV3a5+3AoxI9WQyJNyRkQJa
6IIwASsS0G5qTNakl0mXH56Fd4Qucj4CJ3duI7RScVB/cmrwDwq9a8806D+zQNKB5UNDkehqpb7T
8ggSDCEhVyqI7pbPM59GJUadb+sd0pDTnCjimq72ANh79BNYO82NZm4XeOF9/KdXFKeqKihZXQ6H
Hr5NWC43ErL60gNBNjNXozZn5RRhgIia6c8ls3mT4xDRh70AVGVyMVn41wGF/VaMUlIWY+Jvzf3i
X0j7+gri/NRU72M+MMF+kRwla/4Pv5MxSmvNqWT7qxetCoBa6T6370HDv9wsNgzWDJw8F2nCODU5
uKq6J4B+8XPWjcEWYYM0R4BQ17jzKHFsnAnavIA0Sb/apa2j0s5bkuAg0dor+SCidI41a/6LOD5k
MCI9a/M4VyH3CqJwW8Z/WldaJJTpI+Hr3FG107kWA2b0ZL7oM8CmcJrG0fFn1ySQYjcVF1nVpGCR
MablSSYkiN16ccfxWFRxKptm0i5/54iGFVqKH0CwFKksGXI5/JGjEIEbC4TTTiUJQmTK6UEMIfzr
jNrnavro17eTCb1cmEyhSV/VAjpuBy63oh8TpIg/7tLjfTEXoxa2PQGa7aQMBBXXcx8ys+Yua4Wm
jT10WezQEpykermJGjwX2rfIYQADz1cyeN1jyGHWD1B3TcxkieJRfkIgY7DRqBtcSOA3hLHo5ir7
iXoXqXU7wctDyVF3dK9WyYN/WdVxkwQRFRgf/4brUZ97ltaQ39St+M+0w9NTlySlhsFNsCIgWBOm
ziuv7TX6tp0qlzwmyIEHGP93fNjYjtanssWrDFR0hUb1Uo6WKYYt4EcrguQpi08UB2p7b6dIStYf
DXrbWf9uUBkZmBaetTprp0FmBfxJpoYG0q47NHIexWiNyYJPuRdsa0qOUkZJlGzqOJOYECaLuOA2
YUZ2esYi+prw6Wk2sU/XD8pu1g91BJdjjd4FRbETBJVrMBRBjvwW7uHwwyVwphTpHkPrAFlhAOth
kyz5/dEWDWc14WvPGM++pogFjV3JM7PK3WKWO2h2ndZLFBt06vhT+1r1dLIAxp+Em2C7qGsTcHMW
a2JbmHxdVhPNMAuiDUwGoNwVTTp7iW19ribbCLPHDMbjrdPjGoye82mq/cIbYP+trDrEPCiOBJs4
v0IsM3yF8Fc+MEOK4IzLeh/3dGbiL/tH23JM2dV/ROSe6FVD7Y6B02wwTEv2t4VV5v36BGltwYZp
84LFEC+I1SPKyW3PIbYcgD/GguvI5oWrTtOvs/pTCZYL6JG4DOHBuAjgIEGi2aalDRVzZ+Cqw0E/
WnZvySfyo8Z6U/bVLiGBw3YPme4SBv27O4OB4G57k1k7BglbQcNhhE21uSUBmNWhSxJe7Tuj2y+z
aJA1CbXtAbSVz8zeXTYMbleq3+EvWIEhjCz7tl46vQAhZUC7dZJaYBLQzFLJMDmCLMCzc38JGRXA
dTrzHunf+XGhasAAzCFsi0+Nwt0CjQjTI6rSaq0+PU6YQtw20M5KWdJCE8/6Lfx18/dxbeQgcSmg
XYbJTUP0BFAlnLM+kAfCnLJqbgGPef/azz5L3DzqPS/hhqf86Y/1pM7/I7MUQSCQ4u1qZqS0VKCv
4E6+jvWZfBqswOCi7Ik2ZE1sgveRJkHikqr881cTimL8n/gekk+kHca1yP3MasjLyl9yFR7h+hPh
kZJJZ2At+wehe1DWnHxR9hfE088m5NwEhWNjZS71ebX8Fm+JgflGZdjotl34PC2Qg43lkKAGgafv
y6L05XJWQZv6M1UgVbrBB0m4piIUA9LgnZN3AwPCV24BZ5D1gnEQFT9iLC+HVH68dVrF78G7zFxH
yn78BLuV4ZtCAXhoy2hyI7LqEHF6TjSV4zzlq4Gn/xZRhD2rRaj3CE31ixA1Ax6TpBApp0y4cMcm
g33LQxAkAZPskID1OP6ay4kr+/WjKUfSGGcuNGr73dYVGEWSTUowGZ28HnJycp8qUpBD8whG+Yrr
0x3quifOMf22Gp5sV/A80GnDIyVvNAx8wrkump+5/OBDzjQXKnzQyzYbibK+yfHK9KLuiPyJzBMi
NbM51y2aXVmztAZPi1cAIuzLqerlExtmrQHsOyAxgAoK2wxihPmOGTt+moksa3Y4yY5Iyv3Cfaga
L0edUmd+AC+Nw5fpgdLaFbgt1KuhmRRWkrmXdAD75p6At//UPgqr0nl77+XiyJC3HP6h2E1DZzeO
9AX/s1/j0SpqhNAAFJc6PnucH+43YpO8mbtI+7f1Q8EJZMGbikZJHob3kIkLNzT6KNyw06C+w3cU
k68YJrm7KHZ6MtdiHLbXwuqKCx0OKSGU1k87BqaiLutgzsfTlLLnKdi4Tg0fVVCKN339Hq/Hrhcg
rXSrkKyz3IuX3fkTN6UUhmgtm7siuvZSKpQ4AbJiq/b42+sevkIcobkDijz3rnYEu/RVvl2Rl4CK
zmLffL3FYeMwewKFkJLP/6ty87jWt0X+ZS9IS53VvnBRFX065n93Bg2fre6BefILKQSWX1hTFVTz
CiepnlGflCSerg3KPWSF2w1UsI6Reo8j9mqn4Rrs+1+1bAB0dyXD12Irls1q9HCPjCUsLofmZRHV
fg4NX972iKWYs9SWGB4e0Qr9MAMf5+KFFzYc8lr/l5/XneRl6zuU4Fzl34vq2kwPXeyRaWeGt1Dw
+6PvL7Icb9iKtYUFEoi/rAyEZdZ/s59RYiLuR0oHayMj0+O/J/79Y+YHAhs85lsFh5f0XzgbWs8j
h601mE6YBCiUdgI1jvQW3yBtPoHBy+hZNUqlHGRklRCuo9DKdsr8xoHvtE+kSFxrVYe3TC2kcJ+n
mX3SpwHswj96K54XyQGX9Vh2pv2ie4yrjR++4QIarZPy0InK85fl7hK+QwOHwtaT9SnAbMvSpMKd
f8FrvC1tNEScdpLqfc+P+jt3jDWiSTCiM3K33X41CU5TWKSrcdtP5pT/Am17FlzV0DxJn2SneMzB
bxn81vAUoyvgyNXcorLx4+1DpU7j3JOZjBbmyRTz7ihKAscy6ERngFJs+MGou0eIL/PB/1oalksN
q6b4ubIv1U5Be4GGORDcvjOJkVhjWpRisiV6tm2wGNgeAiTfg9ECkdnhPhRMI/1NFsAOrk+dvL9c
Djy2zBot+3le2nWkYxHLIZSdFtFPuf0gUIS7Mqf/fco/tSoRjEpyv24bnAw1lyDWwsQkCeavVvhw
621hNzNW7TT8RF6zOSHIaToOVqS3uyPn4O/jXfEocA5H1MI/NzPsP9SoQl4BtCLJ5mLKW/K8anYO
I27tyupcbhimMFTZCcSeMll2+Yt7k+e3YOyxVGZqbcCqG5di7mlbMkrIwgz12QfFcYQF3faDxrZF
0HEbTrgfW1/3lFDOpTWeP47Pm/npzKA7e+M9FKUBXaTdXyXGY662JVlCgfOwmlIh6dwylgFi9ZAl
0+W5KbeTW0U4hmuFwT7XmZOr6Sp53JZJ4cbdG6aJUc7uP1x/GhVovQfWUPeFyTCG2CKs0bebgWNS
RSdQxeqQpOlQwCGYHhm5wBOwu125B4v/hQQAQmcXEE9Se7Fg46fsM2pOOTHHxsszMC22yov30hX8
6kcdblZqFeQAmCCVBwo3Sm7Oy+NFuVexR6sZ+P+uTMSOlFrHOwVvXgYcn6kZVAb4afPwX5DNZny/
kt2IX9wMMyrW7xOL+dTDAY758Mn1HQvU1uBnzVBOv+Nf7q9rYlSZDXDNeaHwxGjUHWMco7VLige5
ggZoYG1tjWfvvhF9RM7M0320nEEcXve65Y11eSlGEGSlOXLMbIHcnvfLEbusCoY0iOISX89te9fo
gBC7YhsJLAZreYIhemlq32E+iWcXe2LpLMIp3y93HFsG0+TLw8BoykyyK2FO7JaSCpabnaYhbogF
ySl6FhekgUiy8Imcvk0xxn5oDQfWbVNhlqfWZM8Kii1MK35fLJyIHz19Nu37z7FciAP/iwyVM6ta
U9VGTg8DIu7gOp3L2DA7BCwVMfRWwhVF4T2d01pyMdlBeMKtXuHiv4GlvMIABvm43GyH8XGwbpNo
GjKEJoPOUEJm19uCjDInfL+q+2cXKS6g2pcvmrfeG+niz6kMnHdig/vaVmnc7VX6OOD/IzYOaNVU
sqn3CJzdZOMehXBothjxHdBVMNMeUPE/SEsSu3BD+9KAQb5hAw93l3tDERq0eiTBJxJEuM4vx/hL
p9krfAcNPl3EEDxmX6j0GzqNIdyShyk0uVZJwFglzavZRUnonDQEc+A3Jeku2JKOwBF8rhSeM+Dr
VToPZV8V6tiVgdDx8G/FZxN8AJ/tzuipmLvCDGk0iAn6qzCzIi80gxZm1P7HFNzwnKdj8uWXBHmw
u9faKAsy7gYgHiE+1oe5pOnbnybLvStbcrg+Yom8cACnyQOAe0ny/DMflxlP2KnHA9TxXVXsO2Aj
hbFeckQzjV62OJVXExIPmmzQmRNK6SxvhObMhnYFmtrteCRhywcqowl+C3PJvq8R+wlxMUTv+kAc
tTyuIsrr69qqFYcf/T3SEDLurITPTVad1qdjZT5AhSvB5Dz5Lp4v1eBtIBb2/zYPsqgWOPO4i6YJ
uPlIBx0xRD2lqXaQBgLu5+xx7MqKrbg4t76qvxTANemwMFIBhC1LiIfqnqP9zGh7KXhkRci19SIl
RWLXcSmt74dSmH6PiI9yRfsAam0yYDrw+P0I7RAKzBIDzUryohCXEEFcdtAldMCdmGkzbaYxyfXg
uf5KGF2eUzgczlRgsur2dfl41Z6sMUCNwO9bvV01Fw3YA7gXiHNjHOmwcvvwhNmKP7fPpgF29R18
Ik+WNihVJPWDsBBNeZC4cKN0qqAzOupaAV4vlxdKKqvfsDZ4CEhPnnINOVkaxdRJF8ScCS7eeHSJ
RcaFMzg6Xbu73S1In+oKXO960FQ6bt7CMLTUP0wEiXIsXEfXlG7tCNm0wDa4smJBkBjMtzTM4fu2
JW1HbGL851Z5t09pyeNz/veIymp0iJls5yDcEQvbGxIyAiEiXT7vLZ7OC47RuDlAn4o1zw7hCEnA
pqjL7uSjrJklavah3CDIrBnx183B0ilqf/ghpLLs18zEpSF/xH5irJa7KqGXWz+pDwmMXCparSyH
X/ez7/dUhSjl4vGca/MsWAMRotLYchkVs4SxVLtpSw9cvea2yucq9OQYUswTWQgvlCjo+r9Ar9t1
3wjOkKaD8r1DJ2GUVM9HcRodhTBcVeZq9YmsKUmCrVnoHiayCC7AnXjyHBJ+50MeXOZu+VIEtYVM
rIZ/XK8vSMDb7ns4PGR4y7SCzCIeNQhMr+EH/bB7JfhBi8v+CRPjyyIbvIP/MkjDHdffWvq8lwOX
T01td6E1Fk6vol6IKvhSxACV7IDIBcHbwsX393Ua0QtrGBt48J1epHz6D1pQ0L1VCrDBhh/yJiy5
5TXgYnw5tAexLRwfIPU057jtdlapE8Sgx44yIACMpstjZcJyzdw6bE11QuReTDYYuV6PaD++lw67
/qv/M4zDZrNPpTibPFFm8buIFFD8BDcQzawSm+J1Y569HszmYbxZK9kjvSy84rKBclv8tJq4VUy1
FGbkIdGryVtL3j2itsagl1Xzrlvy4FrudOKa7g5En/GteXkHHfDxUjEWxoDTpRGmNVV4Io5fih/b
SoRS3fkXYZXl2BxtOe7/oQfWBt7tMe87Ihaho1h0xkuT1TTH+yCqCFK6w0w1qxEcGtMQYULsI0H9
UAodd+ZG9Uih49XZtUtnOU4+tRwSbZN4sb7Mwf8gXb8zXgkg6DZ0cSCugrSlTAQ5+NFj/2rOn531
C+Ecy4Y6mjfVXh0eWE2D+V58jOv19sUzmlQ+i3wZ/lYieIfSzrBn0vNBL4Ym+zo6QyfVnGSrppk6
emCXTPCKCF6R7Vgt4j9gFR1MPViyKx6MawZDbHFXLgFc4zJYKva2+Y+XDb9ntv1gidzWotBCXa3C
ccbJHGKsqteiICQv/23OX6Fvepin8/opUcbMwECkv25AbLo3yBcl8ofWPIoAvR3xuOvnSrCpuMMW
pqnx9L+lykutyzDndbGe3YGr5crd7IxYhU9nCSwLtwuYm0EKCoz+BkxXGTFHYsYquyaHI7eX3epA
swIAhraNdwtWNzYWay9c3MdApSRTM8K/L40vZ8qZ0h3EkRblTVvZHhof91L5ZSGGroohy3wK671/
HXtaW4dVtSJPe8jtNXI+3oCtJGCgMJAeOlazdcX3yoWQSXASKIfcaECM5vGElw1CDOcObtDoNlXn
p+vt79Jy7laaOJ93XrGVkZpVWyVIg1EMmzPxQ02871gpKH6QYz3DXBQQHlsSXWXuwGjH5xdigHzJ
kf/t5iw76XkOzGjzZO8H6qYohFMkJ7JKQkNGLBu+ODSRk1lleltQlPuhjbPJzYUBLxWQHDPjHXEg
WPPYn9Ky3S3DryyIh71ho4ufcaJx/JmgoYlyiJO6pC6Le9m9yDdvmnocE2AsNPEn4Qg38e6ofThF
dSnBvOwxYsbdggQ0qgkY3QIZLuxkkW2HB/hwZwJQTpl9p+Pcf3KlxTwa95oMNh4V0Tg2vcsnHfYi
LwV8SgBYS0Yw0fS5pLwjVlaYce+RQG7rrsNmWm6avxN7YJ8x2eS9cJSNLn7G5ZW9PSj6sLWk7zYg
atTc0Emh384Nb6mf85WqqsXTPwq5/geAB6W34lKJtqtOwtCD5EPo7sdupjgTNLIpRHYfxfbhNcTC
Mp6sjh9op0hPh+u4t1Ld0akxJtj4gksxppeqkmCBM3h2oLsPDoha4mqCHNmycP4jbiNEvyqM2vcm
RlOqglkIHJ5BcFEqsYsDg0g9upAMqa/Kc4k7Jd3s1BgjhSGXuRqmdX7LSX9CTljklPp52FjavlNS
qyGRWWRNgJwN19n/Qp8/hXkEiv775UpNHeUGKjcnLNxI6MwMkjzvW54SOms3FZal5Hd8bNv9plhI
eQR3fwuMVkwbSJuZihGLit3cZA1aIEf3nO0HZL5eDxYO/GDCgJpFQnkWduBoS8/vLsS5ma6M9bZH
No3hLljcELQzZ0IthUC4n+Jr/ZnzmAf34kaNoG04clUrbKfnnhfu+qFRAJ3aaOQcyVJfldkyvsg8
fCBkfHMfo1NvrQgqBcP1JesLwZepjV8DCg1uhJNC/kih4Hd3wV+Q39l0seDu3In04iUvVR6crV+9
CPh+7JmOvYFyZHl3LkNxtt74GnZ6O/RP50QndT97NIRamxADpEw6QKyRF/68XbrourFli4E7LCM2
tqx+SUiA/iooyXWUC0wYNxFkZ7HTY8ZnlueLLoUr8hLe5IFs82BThC3yUbbHbFw0PZVdJRNlNJj2
RGAr6y6WkKKEs0KHln1mubJqr3vRH1NmjXY+Lw2RNZOBIQKoEpruv0EoobOuQ65vdGP5j5gjRp4W
59gCbDTioe8CviKN6x4b85NvajcAI2bPc6+6MPZB6Qx2M+DFf1Zmn4RpwRvBDFACGmZ7D7mIHs9K
c6V/wl5Z/8GnIsGOrbiGNTK//gebC1dWE6ZOAxbDW22ewoU5EDo1joORDWcPpPIEXnD0UJWKjSP7
UpWsf0DAKSH6nS7lGLrpeU3EmL+NIqPfCLzCeqDcejbOs1sNH07k/WSmkie2e9M4EsxcX9IEvZAR
dtFWbjZyIYc/1wCT5ZYgCgr/DQQj+PZ1WBhO4P+28BGWGA9dOwmMnf8U46oq2nVc/Y6XV0QVytBL
gwEUEXi7Kw3Olw3BzkldS6N45xpxJlLnQ7E88SHKh5VAe60i7Ejxw8CL9KjQ7NUqMbu2quBEuLb7
Qtg3xRS5781xcEoIZMglTrINN7HLJeAlaZUBCOA46+xGO0szZ+oNj80lEu6c1S95TRmxLzEdfUTR
+XahiEVVTMa7WfGuhfU0xSBqZTmRv3WoLpk7uWS2uoX9O5uIQprIz2Tyx/ETUURCFzsI2l6PoMQG
03bo/LBDCLk2w0+dV8kq1Viix6z0WKQCwg5BDyy2MN+Fz6Wx0/Z5aN8dvK2mwr04KfdZ29IfUNiB
MDJ76s+rMHfW4ubAsKb9bDml0uYoIE29mD9LKWKvw1++jP40hhjTc/ZDq2FOhTGZN7hrRNBq6rIZ
9wafxrzcP/t24Qr+Up8TjLsrcBUtqeCFGNk2g+hiE36d7DvXToQsBv/GPbL4GUHUcs6oOZkkCCB0
uKygAcE0Nci7cReU8L+4i+iWOTkMk3ygyRnUsJIagih7AQ+DZoNDeTB7q8B/PHDKRdKEzaaYuEO1
9Jaf19IwrsUsWaoPagBVhiwIuWDoIM9V9GQx9COoVPFxLXUfqnt7N2fAel8m2kOxLQWtuoV6BWsp
BKAi6I/tXncu5EZ3X/RGJY8K6d8UM3RSddsZ+JFsUkmQx/KnqN6/QWbtii6GhwoaTJK9VNyVcYW4
fgLkELWbaVxbYM6UCskbvqnDlry3EEnZhjXEiIyfI94neMcSfU3s7O1VDom7VhO7dT7uys4GZE69
S5QsVvQzb57KE9aO9oMC/X7hnnRIgD3LYyFoBD4tdpJTiZsflweKuBV9wxxgnEB9vupclzk8AwhQ
gLbeMg6E9jO5VKPJhlnlNB033RaBg3easOvZtMqn4M9s0SHXSmLV3TGgHzSiLSx+8fFaRbag+y16
zg9IC4B219Yh81wZbu7FrjTgbgZc6gf+PxjvDnAj9HNwrkt+DV3JMHA0Yad7hIQajgGZ4iqaN1AG
CiJyCyUyL++Of4zrU0KH77vlEawJKMlfoJc9OKj+lqQbxgFv6ylen8mqoO1Dj8Guam70FN/+I+iD
Z05VYb8NAjA947UR8BIQNBEhn7/een5ETZUdxMpGO0X0pu7UF+y3WxehRZY8XfhZBdw5bpL8YW9y
91U9/t78vrO5qRzWYmOMm2HyRFXkxhZyiJL4uylyi/Ys+mVjjNaDNIPaake1bp2WQQa64y71nwrj
ZUUJFT79cscbWAYBPSU+jf9RhbMyD/INhbhWZHRuzkSlJAjhXoD2Xb+aXTZbq88E6BdBfGI3iRjr
GDEoaUYDkofz6NXwymxok9nxx5ICgj4xC/sECUv6LRdg9nswqu8wbtiAAhgslEG1YQIeso1v8SBt
iLgkikf6VqAolhYGEPtXM/g9i4QLh7hSfb+5N7vkzG2eNm/w4JFrKkL/b2gVwWMNUY6P/5wVhLB4
Om293Y5wS9zBi+I5x0dDVWU56D/hQNqshx3SAKZXgQZwR0tQIKAzYxMFcsKX5xfsMJlY5JcIkCad
0BvZpGG288zz2v/aFI55V2LQhDCWRCXfo6OIFXfSGf4M55s9suhzJSM5fN3q0F2Sb1d7miJNj3Lz
7oa7ovhoeAsWqTypopIaWpsk63yzl5vWeg6j/chmQVX/TQqQ3GBsQla2bBkXZwqQCtm4SDbKOOAQ
R0tSmjBwhBEjqSEEqOrOsli9HVO9mKkDnA2iP1rKFpu+/ZOpCs5kDHjrWo46T52/G0X+ph7xzDB7
L3mTJG7nTZLRCjlRosyVyY0WEwKTsgg1ce6gF58eh1bnsVmleFyTT1Su2vypFq+lqSGj3w6vEw0f
/GWUj9or7Fd72tg/BZVtAQRlE4iDJiGcterxKfcWl3TStR4bmCWqPftaPRV9MuvJj8D7Hwt9WKaY
MjEz8gv+OguAiOcfhvMIERMQ2JOM3JzqfYFiXqDEAXhHRhmbbif+D1I6eynMtqOCzIYb188V3Tcy
jD/lINL4seLylN0xieNHzr8bwaaKlhhFRDfYLPon0IZxXGPdQaPSi8GAGJ2EFvCXTYy0aVWcCrXT
m+ZkNU0xOpKSwE9qjyV0s+KljdbFaV+hwOuDg8xCwnQZIheou0YTFdpg0REAmbHTFGLiIF8Sv9bX
ilqurniloJfh0GQ8afyA596mw+bmG0fsdzzPbpLAuvwN9nl34UhK48sEaUNMzwtrYZ6VOSLCcIFr
7Vy9mS48pmrVxH50Fe21ibZlx3udmEzivQZngLEw+17e59u/eY6Hz8T6tZgL2J1El4ExXud5UNtt
UbN/O5BO3QDgYdhC1H2sNx1Rmriwx731MQ10RJx7dvMI1oKd+dpAKMjEBdUXSHycGXpi/YmaTNZk
qhI0jzrsKJIqU4sBi8qaV3Y7rPA/cDZCqWB784AqtASJ3NYyKhqz3UwAyN5M9J4A7ZZbNR2wkwOM
XPn5zVY1O3GII4En5+Fpl8mI3mKTzLDtVA/N2WGnnNX+/3OW2/oIpD67EKKz4JGEDj2GkThAtlMJ
0l7zit6P1nURX2FbkqNJ13Lb9BjMoVJhO1L2Cs3kj1whq1JDlTrgiw9Kng3qqRzGTCWVT2wtYb65
ipCkOhFYjOgxyDV3NceZi9PcdSUO7100Cntk+6Q4SmsWQvhm1Z2aLldm5EozaCJ53HR6kj/lNls/
ynggz4lU477r0EiIoc3MLEovjNKyy7Ts2hb//gPk6D3Xkqnsg2jKedzTjKC7SIRzfoi7AJkzY6Cl
JcXf9pR+WeLUu9Lxr4BNR05OPEqmrfIDwAWx+AHyULX/CVFUYf7X5seIvfI0UCND816QS9s+keMC
Ypx3Y2GJGp/an60aigjKZ1+7tMQS5AxTITLsrAH5152oVSMuCeYxrAzDWocE1AAONJ69bpOJW9I1
+guUD36uylXW56i+F0s1CrxVr2H7n+zO03nDbMgyCAH2stqJRSMsrzVnRiajqWWIybD9s6e4flfi
A7Sp5ac7Cm8smyAxaTXZuIUuDF6rJ2TtO0uPiKiwTF6AdOn9wwXcswUTpSrNsMz2IwpeYq7z7PyP
HhXRfRtNeZHPIGX3RWCd7VRdAOPix3jxTlsuYFwfzUf8mWNyWAJkutEK84GQuBPuDAKl8KgyDXhX
KG//Jo9bxAHcmFd3ZIvO0tsmBUBJXq/ZwaDO1tYPFMNJmyE/PwA4edYrlqH3/xqrs6uFzgAYLUZZ
MQsUG9K5xvz0Nq3TE6itS3fThwo8R6HzqvJP1HHaJOMMdqEcaYoLKEXZdLZMNMrhQPCWvb4ItiQw
xg9Gss9FeHR+/9CxvLLieESa8wV35kJ9DjWhvLJ2Kz9sFcIBq85nvXg6oPYl8g78tED93Hxgmy+W
ROEjK3bAwcRpL5UX+N66n9MhRuMrJv6rLp05MyVIvvCjvg8DFOYV0fUSoYTKaGom7m2F+4pQsjR0
Gqpq/H9d2zDJSymeOfBB5KmpIXw220iHwoCbhzoh56nkLWoYfpZzUYNGNJlLjLrME/B7TwAji0XK
Rd0tezK3CeZ39aQCtppCQdGUt6e31BOdPKKrKP63UYp+JSfdr6JmR4F4tMseNIdIiB/IpSedJRn1
bJG4Ri7Oc1jvjoBY79Cj7OJhvQ6XVbJB5F4Jh+uEj3hxEiC87qvbhCK50GfgIZJmz6R+LBln+2FS
qT2X6txrBgUB3TeVVmpA/AaD4mkNbx5TalU0RT8o7IUCrcsIEYPWC6Ez/2NZKeIeEqpCXlyeI0Z6
7+lciTXOkYDvFaGyQle15hLCK3GoFhlzd9jvMlVmVHs8d3Nb0bRMT1kg4BVNLTAksLcR4kQyT0zN
tpMV4JBakRy4fCwxUnNzVULM3MDn/Ll8pd+4WbGEROf2WcpFK4MrqHDdbTXNe22+uOGKZglyQJ+x
q0bG7atzBaxK82bwPoDLO5b76VvCPewhzgIf3YsvqnN3xpE3obXTUZjAYz5sy2O4XIdTUV+yhol5
r0IFD1kTLvWg4qtiJcgLrgX5IRTDH3TxZ2ZwU5OXj67SdMh3iSibgs1QNNfPdKXDOD6pT26Dl6ru
O/gxEncIODExspl99tewFcxnQJ9mTN+OfkRZpM2hpirm/v05dJOgE4026Y6eqDziO/cXf+EnfWB3
XCD5KdS71qVsHBHxtdOVb4px7MCq4gGW2hfI3BmM+qsQhBki2dF5u2ownroV+k/1Cxjhq20sjpIz
6PEgFpIO/BpKBZwe4zT6A7jWUH9+qyetVBuINWyxe4eE5vcKdoUDAUNhwsOBd1C0OJ7SrRYIhSMU
Cq8cZaVEF35BpmYLUGhQ7h49P9ndUXnPvvRoaQZK03iju9KpQMl5al9rCaATgPlyIQJHy7OIZPzX
z6Q9veaVqQs5uGX/FpFT0B7Fyy7Vj9ciw3OVPV+eaVzKHqgk8JTYO2r9NuMwSdm/s6qrWPGFnKBK
cNHKohjpvqHObLPcQCVwq4mu4HQbFan4uccMqK45kCJOrqHy+jdqv26U9167D9iZWWlDYusAnXH+
h9P+evPhK5GJPxyqijsxYL9W6pI+Pn5MCQZ4RSSn1hdLLagywUMRRCOy/4BkC+nk/ffRUm6mjftg
j2KMjOrgZ0Mr9bSk6OaklVUOH6IN6AqU01OLLchG2zWWm7NzgYaii3fAoe64iRC2sGBhmrmC8SiP
m9PfMwRDgpxW/9hp/2m8L4+H5YmmIgOFGMKtiakN2v4sBNbmMRvQsqk3c44ZeNEM/eHyETrgTQgh
ZTGePECLJpila8XM7KEDnePR0JF+FEom4Oqz9nKmhBIPLuwLD93zKSWFzOsMaFWL9sn5EdUuB5YO
hfwctnFPCydUCcpWys825UDOtaZ677k9pgVatBEVhsv3ZCJNNQzvxxiOwCms7qeMFA3OuIonqCsr
UPuo9to+/CmR2pa/Blq2dzFtlYoR2cnXyJk2IHS1c2Nwu8IewxuKxufpw4xKjN9nBMg1kVT0d2fN
qN0ASP9kMbWRPsa0547+sU+JeVhcf01YcSp18YnPHO3ZshQf7BupmMjOptbRMeHRKTGqxdXDh2jS
eigQVrUetsNbLaJhqfilhQAAGMXZVa5An6IEQOUTJpyAkzukjUcXnAnsNA5t6oeuxrBvs7+EOHOl
WRCEjGrSmcS7TSwXUBWnlPX4neMNDUGOpHnQorVfAhTGT6XLWi65Dj5aibCVdMLrB3TvP5lF/Z0v
WXz+YfI8U6LoatPmP7OefHlLN2JcHahetmtutea8ekP5DHNVmXxWQvrgjZPrv+qBFWOdBKAnoRKg
Fvie+i9lI31s+V1/9VgzY0mKThsWI075hW2oP4Ynjaz+7tmvZGWATkjtjsVIE1X9/kEof1oBRV3L
jekti4JRnF+PqWpOPdxFgTcIqGzMqdrvP0Np9DAEKyjULLr9X4bzgRCF2Ub8F0HpJTg/5PM3MR6S
yGiFQg6GNNhYHErDtEf9FN2AD7bXo/A2pV/zSJvZyjSXCH5/4qO5Hy4s5dAqyHooe9RvsZExv5wA
RO8R4uuk7FrSX/7+fHtr+O+UJB4gLBVVetH7gUFHAvfcgq5TiduXKMAPBAkH1gKSaf42Cy2ul8uV
bDxt0/DKB+jWU/8Hh2bA0Ge5SF+6GlL38hi8jIpe0cRSOjEJHcXId6lrt5GInduXxkUQIvFVPcDS
bML7YqgoqyXCmrCO8wSfucogiOTg+ORmGCmTmUCCgaIfE1q4mQJbPvHpW1k/4WgN0n1ZrX4pBjKB
c24m0Oub83XMs9G5Ne608RQxZi9mory2Tf5mtzVJ9rei8SZGx75rlCXQpeoiOoagPJyRW1XUADGU
ORBMInCPHHM8e4t3K272cBmNWlx75/2mmml9GCyZVb48UJMEaL9coAcyrChy7K935cU/gpWp7F8f
MeNaeFXiKfC01ZocmeGJB4y/VnBaQ1HBCDFrdpSgMe4nrxM+1EFNOnGKhFkbp4RWsh0bYr9Hm2Np
kxZOda8yuinevAFj7iREpChOT+1BM+pwEWu+hliLSMerxFH/tyLm3XrweZYf2D5MShfpnyehXzo5
DA88oJinEg/3VENF6VuRAQgi3QFO1aUicMP9rjeT82wdXyqNz2cwkj3cWSDIaJ7bRkrPrT6PHz3S
Q4VYx/swJlemburW3XI1l/I/+Z9dE81dYmpK9Yr4Swd/Cnoj7T7daeup8NtHtHikTiOFrJXa3bBr
yTX3GMg1pP6Nrl59Y/nbl0ls07mAHv7KO7eov/D2o6TT5VMYLlLX4xYKb+g5m8gSsfMBhP2nGHrH
UOUNl9dIsQ3SYdOY0RlwflP9hcIGNxBBRkzAKo/uG+OjhMH0acT1ZqyE9IP+PdFJR3sAGjBJCG5q
0fwZLBOpBKaCczAzUJ5qDGoXXPEH6LkHUWfjMWkJIiZ3hqBkwS+XJtBFFnlGslS11Yrzk84AALPd
EsqABv2DKoGr7rF6NyRO8X94RjRqF+fiKDc6/BSw9sjYgIVaq46B6uL8+26d7esA3Q1cVMI1FNFP
IefN2kjnXN6LU5aGvuPdLvFZrSeb0E59gZ/xdKWH+gof9EdpVGSTf8VBiprNjoEVstgpyOFI7jP7
wRtUL6MTRaOqwpSbYFuh1AOEr0t/7H9TWO3RC71kJ/2ezmTfnqo38ggO1CcfxhO6P9yA3WQ+JSHT
oxCY6Z9h9DABPqe8uLxIJVPUWPEYvnGB2TkJis46nrREn5mSfYz34nleCiUC7k1oOeHYjNA/+Jfc
fAAOYjLoVpAfuPik31Vs0TbywS2jcmEB9RLk8a/CfCPowiX23iNr3IlErBcL+OF3YXNLCFtxKnIi
0mtBQeI6plXrIHrNRQL1JiVhbBXwPF4qhDG7Dcdu7EsCEx/kpcJGqrIX09Si9tbrY4xrtNxmmNFc
kVvo7E8BvY2a6ALf0GUsp7BFZzOd5AovdtnUe6xyYmaUeO8ZNgM3zWWU/aGHcFKThv/Sva0KCqrv
vLZItRwNLePtOnPW1qi08TI3cKb4rPigrfIHTQatICWyT2quxf+betR/3rELZKEa55GaO+wNhe34
mq5Kl2JYUGz7enUwFoBlSG7sQNnHtO285y4+AQWuKxBXidUFJmo9725GSPY4bFx8SW6E5F+rt3XK
e06u60OdiNW5I6JDAQQrIOjGju1ppxd87ymdtRyPm3pFWipk9HG8p/W5Q8bwzh4PZys7JFnrhZD+
y+H9Gt28RnxWPyM2XLO/+mQvM+67GLR+4XTB+2qdhhVnAQqWKC6X5WGOVOZWm2axj7/vQSEiTzK1
hHu+V+seGZDD/zC9toRzlnMTdPxv73WANOWx7Bx1BtTwKiQjejSCLwV4bshWxcRstEwOL9Qj6pEk
NEHaBkG9cEiXAC89ye9bc3yg+JNNmRMfboLYf6BPkpqeNaFeV1/yJqBNds87JKl9PKs5evFyg+L+
mt3khvCTsamqTR8PFSgKu7nXSidJlAepvHHo2BrJWkU93QQmLoWRT0NRgZAmkGxUYOy5Erp+35Zt
gtaJw6vkxszS5W8d/EM0Wr+kW3FRDJC4+namLawyc5AQ2pfTN4FscvevtWYkXlMw0uDuCop0Xz7k
5oU+uxnXbJcq4HK2lBQ3gARxXpGdpTRls2IzYDo1eaULHQW6LY88JBZ4KI8w3WmQJGi2+bkKlXgy
z61KYEuEfC5NeIYZ5W+rW/Qahz4D349pDcPJSn+hmeDrxZbBbDRQ4VuldmgkxKJXu1L3+49qZ9mj
z4j1A47O/ZdvzkKzMQXP2ohpoNdf9bOGl2Pwyed+zLJmHaNuzrKMChMM937BGWd1zEqWM7vyG7Ow
CpVie1mdM6StzR+dbllKLF8BJvhP2yxx3sG0m2ZIp4VORDAyOjibF5blMaQ1fwiOnL8NUjU8EuO0
xypRZss5ZIkphNua5V6nEwGHGY/lD/U/LLAhl1I4oDU6LRIlirzDBI1hCUZIRLRad3Fj1nxx3kwb
RN2nFRF7dLRzIlHuDgr1d2Jb5As2Dy/OV5k7PQ6FHZzd6lA2Rdk8FEcXwG6LZz8fVetg/3xy94lU
yBiTtp+KmgTzxzFSLHZb4MP2O6m7iMS3g637NMKsLeIIi4JMEM3ergBIGztMZgi30qnsBxP50yAJ
sanW+oFAqBlbsJlBynkZfTHyfFUv+BrQlQDgUVlfVlOWanqjZzSISVYwepiIk/WCiidYPYuJNxh7
AGZ7BHYAckS0aZkQ4obrRKNWrLVifcXDGT5bsu2iu1HCQAvK70nmqIqo7lKEGZQ1aC+5gK7E74vL
cgHqyZWXQdqQKZ/6tFIJNb0ICnOYRz7K3MmVyh+clufr3iHhu49wQVoDSZJqAqATVGoX+uWt36CZ
iH1SqjXyDdfI7rhee6+q/UjTym9u/intL4EvPv0+oQsgO4S0zK35CDeK1BIpsVs6QCv9ovELsCyf
d27kEnNPzyGKcgso0cRK08IFDfDEhX57PtTONaGurdAOPB65oivgqsM2zapa+BmO61rPo2MLHfW1
VY3IuDhYQ703TU9XOgbomBBWo+jjbB6kMdmaFgd+6C/eYhtu80wj2TC16TVycfafJw3bdUNTd7VK
VxLahVtshbk4nDUzer2jt0JLK/MhYeU314vJx1q0NLsySQ92GnLrMmmjB8lXQ/jwOpLFQMMMlPNE
lGOoDo7txO01TkiN78TFs78COsrUB2lMQHmlizZI/DwgoyOCKmDbJpqbKCwZJGpvhSesbMTEVOcy
gN3zbxwyfCDITkE/9sgRVwbNz+0XRpUY3DPD1wq2Ro70eFk0vhOsqU4bTX0fGsD1xhZkLW6Xix46
99qyoNwt1QgLqYMWxxZLEo4mnAXWhcWMmoO45Q69HbmAXKhwobrAgrCNXM2rLG+lkI4v+xxuHuFV
ND47DjWb/UNgFYntRLb2uPP3VJXo94F5zM5oQk54O05s/1fsoN7x1krq/0p+ZBTbuC+vjptcbEvn
Cwv9aeudCr2Qeuu+PIAyAJPbzXqvdyL7LR1V+ojm/tEyLi1eDQwDv9UNIO1dEB7qgXNdCpRh7Kxy
lupqV8mJzNSni3NLeRYzi2sxCZxwY6AO/+W+UaPuaDAgtkAyAvXxdWjfY/cfvAwZK6y37hfaMb06
AHCs1G+g2MjrATLj0R+IjT4YDnRnBGqDGFXJBpCr8QeqPW8T1+4iWYrDFYt3DfiyfLYBqNgvr48P
0k6NkBjizvCe75/mTdXKchMEbh3WC0670dX5sb2gKFXFCsX2SYQZWRb5o9gaq33MRlSaUUpD3Rjg
fO2BcfEYhMbSw4pw0BG+Bxy9dD1g1dFZgPJAdLgwURYHo0ugXTARn+WwJzPWtF13Kw8cTGhmjWzN
8u5cwua20yJkrMM0i/ySYRuhk8ByR0qMnsI9flNpUiJuO+FmCaTaEt/WR8Ib02g/Op222Xu44F5s
ZfjPmqIIcleR5Vzq8cEN5gxYuTdezDaeK4PJzX5kK9Zz5FYeIIevT3K3IM+xdISo733Z9yhzw/jK
GmvTwB+5JG0o+VARYuNo5LtBoHEkl0VecVmopmSCVawxvRwOJvnmxF/v4xatYf72bUKUDVazgwcG
ypJjjFYcZslNuH3KeozXPwfX4CU1HqBCSa7oDF5MRRi9R1N5iMPBN/UMyZiNLNkzuXqcsnX287xa
OqhaZZT/lfSFlB0VS4yKsq7xHWxuxCBqJFaLiQ0JYTaB1ooV/Mmj4RyzQBXFTpqN9jncJGZb7wRr
uDQJ6xw40WKY/7msSrE0Ng8DbS0iA/7RPqDObgd2HlvoRFWO2+5b/aL9/iTtHQenbR/eHaG8OY/s
pngCl9z4kE2OGmGZeeI+yXE+Dp1OOcRnJ9Uy2N+fvWYkpjg9kvVAJiY7TtUyf9Qln2wBhJDYq4WE
swsOjZn8ohofhBfs7Y0kpZ0AzgeSNIWxLdBxoNt28XFMkvCcp8Yqr5RXOdPdS9Xk6sDlP1gV6y3N
fbg0Oecy0mzt/e+YGFxL4aUFzvdpvbOqKlX0e42u4DExjB+dJQAxd0JYbcOR8P0Q0izciyStmQfw
m9tbBGHO1H9Sok1yMJ0UOXuJ5daLLzD5DT0kaz5jsdv8TaGvvcSLghaC3iVDSJKoWQaxkqKfuEzv
R/2Vv0MA1AsxRjiXAfLjN3W2ceoJFX7M5bEh0HfBsNyR+0jFktvbEbzAWgQVyAxP4KKluYViJnCx
DhoeXQP6oVe8TUmPZhtxtxAbkRitWQS5FiYIbZI5iaBheNkkYS6SPOcB9vEF9IxRGFhhQCZXX8Ca
anHaThr0R8Vlk2t7M7qKNnK4G0daJ8rPJ0Dl7zZ7flDpoPi92Hr9FBnMrnvwXHvl5r5U9HZVlWkV
UgF5BoPoM45TOMmN6cm9Qamxy7Ov5kMho11rAXPouZpJrGb6DDQznEkWDAkvMeFWIE9gGfJap0wh
6IyFDOUijPHI0vpa2z30+3EStca1VUhZ7I3vcf31LcSRCU1bxoa+rZSCEleDsXFwhzPNMeH6QARW
K06zBy9f/MvUx1xSZJ16SMvwQbcaz65lC+woGfYMyOMbtSVYDgCCW11msM6xE/IRtxOL87oB0vu6
fUnMDSvHsS9nQJ3PH1JUcyDk0yddwDFjq1ty+leoVnR+8C9W9DSWWvCzxu4B9mMt3iYmhOjeuh21
NBwlPnMybfSkqpeCINW4K68uTocHo9reCC8iE+brNVg66vsvTPzBQfUQyZGVk6ZrlsDmKrbgP4xx
tvTfMgpHNYKHBrWCt8KRVFQ2lwKfwLQ06eCv74fBH1s2+l/FBQJI9bYNAfVPqT7eNYH53va7NtaK
V0S4KDSwz9Pjx80+PdXQf+Jv5coatYmNJ2eSVN2GWGgBK81iG/w8iMLbRO4iFg5QEcadGFpJJR2h
IAgod/B/zTZeycI2H9qsNC8Cs6MHjAyWrSs8NKOWsh0br2DbunRyUdgXUuJB0Rg/yLS9pNwt1FcR
f2GJVNE+V9T0ubIA4heLMUgGMmyr85Sp6lRJ2PwQ3tHkJH/HG6IQPSaU3+EF2LPODl6PipYx/E3Y
Rd5gV4TS7VqRXJqc77P6WuUcCqLYB5ntKYKJBuHsro48R6mmdKWej2Iw6eUckk/OkJhyJzPjnMNw
HjlEtgeCbj/VHlj0dBibNdJTpkYjhWQ1pBPp/DOQRSP2Hi+Wooqfxnc4ZcGMjx/SP8vSGTn22Dq4
VcbSBnKnJA/7vEXUpC11oAwV2ceBRQfdXOKbOuso9F6gu5Lvpnx0GppyXCZVjV0yS0yfSmWLn49L
KKsyrsyQ23svC0k1d/p2q2aLiWONpcc6oHG84ql/YMBLH6MOBvS/ynXILenwccV6soUl772Wo3xa
0z5RDda2bTL7xcxrSPXoWuGw7JhB+y+VDwjKvZyF6sXEouyO/tJ6dMRHSUdetQB+YYaEIOBOmZEP
Z4BhumrqMjia/iIAJ9SuOuy8dWNtJJqq7VUr1CaFVIaIfVMMTD1ZUNm/Hux9coacnEP7OWlzpKnq
vwus7MuDEv+Cw2f9U1+9ObKpUMTwreGj/VUZOZUmNJAs3lgKNxvF0xWPWM1VslmMxMpsajeGxB49
JdoEL5py1nDcBzt1pcJ8zPgYBuZ4EDodEe+WykXcXRs5wyJsh562hF90B5RIu2jtpsCKxqyWr12e
YZLHrT1+HcLI9Uw+Ct7HlAlzVF2GcD8Qq30HxyPK8iMTMhRhhJ6r2TRPcbO2opRSxi3sq3DaU+2j
RYgX8UWTOUwA7P2ZU5O2c2lIGF5LZcnMGBvcugDfxuzwObMu/WHL3LTt8sacxDEbsfQR9dVdIvE2
3bWf76xvGutjeB5eLkZ8HmZ4b43fefzxtwqpfLBpQJKnT0lQnZ1vuItKSHUXK5Cbk0sbYmANhidb
41lS12O++jZ2TL6h+J2hCrSNtk4xDkjzLWRpu75vLp3hnKKYneR/xH4ujrQS40pSWN4UJeX89JM2
rJLj6+2t6JDy33GtRxtkNR0IdMByp/LtaFtS0Ju/FkkNym+0bK7BSfnHmgio3kUFmFL+Y4D09xrA
eLRBUgw5tGxZY2O+FPglaZZFtbGjEZip1ePm+xiIZf0pOYxgR85U4ff2t/pXNBnKjGaXbam2P09J
0c8Eeo0D+w0RZpcrPDo73X2aGOPqQQ26ZZNB2oV3ajldlWYpO0Eu9kgLBlq+6+kBnt1WbC8Pm3WJ
XeS/5Qzz5P9taJQxkD/PVAhPi010dCqrocS13ZzKjCtNf3/VBz8UGePqXl7pidvWln8B+fdZaIl1
xXDCSYuzQ0yOh2Df7jw4FyhgIkwcLKw5d88VRXp9MpkZnjxYSSc1t6iPiVH26oBZCopSXX7iH5jn
3pQAcx2qvaHwtWtCRHgatWv1f2H9IGxh+50DTXpsLzEbm/Tn6VveloJ+P/HSp2AVeV/kwUdbRX7I
BcofDSvF1W5zU3fCpQa3Bo7OleeFFmR1e0I0CN5rPyLM2BsBdTzEi52psg6YaG7nfeLxfYJsTWI9
onO/AOBsFbtHiXlex5Zn7VyIZN55vqpskYEHhf8pcQILNXRq1P3tXjlyc+gUaxRUctEZ46hf2hgn
LBpYTlqQsQVw0qwnCgkLL6idhIc/IdBtsTr9zEGO4AjWNc/lyZxBhlF9t172+ZT2fEBMb7iJjwJf
fMIitkrY8MI1DB+OUbZf5zNrRTe8vDSRf2MIaSXxgU+OSSOQikarDRP8EN5yUIBuw+yXhQRwVy3f
1JFDxkpvuWZCiz/UImo4QONo78dit4aPTcChlhtxiqAp+4/sLsO3oVyOsO638oJahSoSxpZRCOSN
EHB/seNzU0kRDWCqlWHTuS++bVIP1/rD0VSorF+5YHi1ak5cD2uPZ8sdjzEUgSafIpBnFfCBdp7n
Gzx1zLjLo5L1ZAWMNKHxjjfNZ/pIqaK994k6MORyy4hvTUxI6kWiz+4Foj7yMo7rkXg3Vtqyesi2
0ZTNA2zlJybn+IEhlwPKlQeeTYQSe+oyF3+4VNj+8uHTIOlNCTmI+6Pf0vUz783rZZEamSz8S3a0
EAPUkRhB8n99aZU/yy5p8TtPuj58wLiUC4h9sOpYyx5sIUa78LGGW5AxYq5x58YIfwEM8ZP9tzw5
jGvEuR7MhyfH1yU5UiEgEsfjEAn8m3Nmm1QXcLWogXzIaxM2sXbPAb9Ul3zrf4LLAzCid3ypFMVp
kPvfzABYWAwD89dBkRyGxDGgy/gIDuIkhr0HFifWAD9aBY6n3v/nojwyme4hPE7SPgU4aYSE+01s
HBSTxVjgHMomd86XqrhG+gXGo1f/nzTAV8gfbagPdyjBcMuXUGS5VbgZ85zbAvEUAhGnArD9AFSJ
41aldiEi+lq9FxMgeourbYtzTcyh+rRao855VVt+Q2en/Eigx3NFqd8GB1yz71hTFGVZL9zlphNM
YW7hbxR0RjUM5okn/JPa+a0B8qQM+aknA1OAUoU26isbIAhM3LKtTt+uO2CqT+RucxJOgefFkfFa
ohmYS9e/RaU1odhGO/2LC/7RSXs56Tg5zwCuBSl7Lh2fMbErEQWbghRXLdlxw42eoEdNKBqfHsKL
MUxp/EjMEKX0YX0lkU3ZsU3zmwoEB1JnHLUAYbX5Rm11M1P1x4AObq0lk745gZbxs2BBQcL8OLZU
4HCXtc4NKlWS6epeaASgAikXyw3Bajrm3g9VjSzwq1zX6BfnctgdYv5WTMrghCORsDSBb9Hxi+52
WIXrDc/0JBOqry0A5E1ZIHBOURVWWBojVgfMO5d0N6btnw1ectjGTPGWPnYs/qeHgeSWJLjUIhR/
8tNhn2Kc3K/Q6RHpRin3IdE/nFrjwYmmcGH+xfmnrdvEKZUjg1SnNFEPnQP61EW1liid6ILiHQnd
4jVrmj55M+kvY+pLmsq2YqJQXVoslC+pLqQbJMCUbZGU2SbbHKuuY9f+1fK9gbxy+aJG1WUm8md1
rpcvoU1AnUgbTO3QTfr9oQsxbc5r8FBJUS1ID4ByjA1hi5rpkENXFtIESvegZnA6CIT/FkYVpGRD
6g32a8giEpjzvZUTLE9C58d0YY5wDK6Hl6YRD1PzVd7fHArVNLhbj7e1yYzX8iIQK0NYOKcRQadm
6MH6iUXIIY8F1Z6wBcP7lXgGh4IV8lVInvtD4KdLBZFDYitJBhUe/7AVtAkx7Q80dXLzsgZhTSSq
4Uv76aF56Gra4zGTt4Wtf+p2Re2zoi9ns2EwwonHR1Fr+F19Iv++njMafub3tJkAeorVhvQaTsz2
/nnNuWGno66pALPRrIAmrTAUZUX3xyD+Qwxs8SamZSmMh5iA9nAxFmNMOHFzNQjKgFkSXVx1Rv49
Wt2vNK0M0oLIcua+B6sn/L9dNCdLR6dFO5mLFXFakbTUAROVAAEkBFvQl+aH5ho+Gw8TPwOXMpYT
10aDV5tTu5ZxSu/QDcenfyL/F/Za982eUYs040kx05t1EBEuikb3S1X7N01pfjEA1qt2hqEDAHwx
VpkBZsgf1XpnzaWRPhFjyBW2+x5c0qOrbkfVH1PJHWYs0s0AADU30f52QXbo6vVYODBNo4K/quPc
IGLjuCvJ1/n9KuiZr6MHhsXlkMuMaNKSdgqHNWKyVZpXX7A78vA0wv+ABFU3i1dFLVFdsk2iDTQv
MseLs1xwxSoJh2JTJpKjXPHVG13P8IBkQJlHleF6C+S2EgqlgBVfbLfOH1eVczXtpIZoPsqP4GRU
G2xHS6YkWDGWVGYQwiQM9En5PkVVVU5NeEKFo43VDiuMYJ/KUZaU8cMZOL8WKBSoJBUL7QiFzUb9
2xkULvJVXYDT4auOzJmVMx8KwnMXMIyn9zJoQinQyPTaTuX4t2u+JLqsUq5seZHKQV7MdTLlhZjR
q8uoSxcVxvlm4CWbtP9qT2V1Boc+4yvlso/eTF5ac78WK8cLZUrnSQONpqWTg+me4eBGJRAgOKdo
yCwE4OSk07Nxh3Ux5SVGWLp7+OWTmI7coFVpYytr4Zmb0GLVt/vDag3FF1UmD29gyqg8cOlafurW
p1iQfEp9g6LluyFhkMjs23ly7UKfACf5/Gj5hr0wxkV1gjk/muRvbI9X2ApJt6qy5rN2ls0cKBMH
Pr2owfW3kqQuA0adjTLFGL9tekGAYXqgmw8wmywrjLzWTUuK4ldXWS64RCjyj2mW5/uFrjyA+Mib
fqkM4lBmA3Ybw99T7yDi+3pEg+eTeg7BJcGNh7pP13Vw+RcnaDx8U7AF/SjgoYTGIOimYsq2NSlh
VIn5Tti2v5FO/CyPYLBR+0L3dDTI3HTB/VDplsY1unsqaVQSY80uL5x3ekV4FB7cTEyt6ie5m2SB
ADfAInhcLx8sRpzkyNxH7cRKTfgAxu1HRhfS9YhgVAJG1Jivp1xkejZXVDXAzYmRx+VwqQ3vXY8r
Cquq35CwHlhAeW04wEwdKfworMyYBbfTq0myyyTpBH8nfB6XOvzzh3mNz0kDIN3k9daKp625hRwh
Zi12SEpccTigmcRcbSkeVv8+usfKnz9Ewck3Uh0jJ3yy7il/Y5g4vxZc2Gip2TbzDENrAzq3bWWM
4B3emz+Bo4jHCsHSNd+vDRyL19yxPUQTXxXiwoSqIsON4yxNzoPE4GocqsNNglpZux1vebF5sJIe
5sB+MqaFde/IyuTyZoc8tYsManaDjK0PCI7HbpLoELyv7HMC0i00QZXYAjEAiswirfXKjm6AMECG
ruK3YcSuKcfHEHO76AysMMX+EoJqDJnMnvmfNvfOO9lhjL80Q91f8L9BhAiWv4qPLEUbHoHyhIlX
CDeF9/lUhTL+lVOwy7qD4w1/sZ2mgzL0F7F4t4o1rM6curvXtkGKGz08DQHHjoWVP92l0Ysj5cd5
kW7j/JIRybA2eKzAlFYmLk03Q/GsAHOoOWQFYj0bCZdh3aJugkfaet4rMOhx41Ttx7n3lTZDGf1Z
StQHTqP9rJcTdign9XSeadeV0krz3vLCZ+42cBniy7iOM8Rce68EMt+ENyyk/ljd8QNUmKF/1uTf
IFBs07iGLts1m9yy59EdQCecR/5oO5ekabyMLYXRnsrDcrI7UVJWePOnc3v+0BRL00QsF9T5PxH4
d7oy9ZWyJma3xz2LsAOYsU+iJCJXxyxcIWRvYpyNixybucFOLS1m5lJ3/lI3DSIFfEqLIDM/OigP
q39sxsyamNMmVc3JyQUi55U2xd4gkKsjGYnhfybznkqScWD9Ya0HxcE3dnIsK0GHzkcPGUiTf4gC
NUsJenpfZk5ZcIPgkd7EP15+d170EcdCnZl6wvGdcdC++sa5RXr8b4Gek4YN0wbcD6fcOxG7E+zb
5E1tUMK69Ubiuf797RpZzroS9vZSlJYc1W5/oQSN3Eznp8hoa/A2zn/ltH9OasePkTMjQPPIIC4R
NHw1WCGxFYR/AdE+fXUkCZvYioKM6unIokUkZeBV7kOZhdg3/pLQlDwyQFi8xmKcNw2sUBcp9zJ4
aXA3nO26KD+0bvywNupQ0rBAXGUHJqJoA/vKwhWwoIGQY4GAbihNMTqKLPuL6yuufw4cVXv3DTNS
nbMI3auJsdtMyACpZHlYTz0umvIQCcAtZTl4/AvFwqJOEe1vOK4+XdReOFHU5DDJqXgLNiA0n7x/
FOsaVcKWK/d7bslXREKAIZeMFv5+aTD8urYa6SO4iV+I07x9UO++mboxt0uzC1Yg4Ij1M0zXm0l8
K9ndu5+z5ebkmSyyvIlRwyUcWCHpyMliLnX00GWlZxr3WzjJCgIcf7f47MAAZO4z7bE6Z2fPufoe
XTr/CFelwm1+kHyWKIHc/BlzfilUhwHVH8Hml8LOyh78qrTRjXYdti8nevkvGtMP5FHLeV4XV/Dw
gvzaeEEWHlYChvAVQrYnKsXcBVLMFsNkZWH7m2W/h7kCI8zSP7D2HKzFKgINY7Cv2bbgFftnfEyA
4jtbxbe2/7tVW8g/tekK6Nd7qKM8RcVuDbla+mfqWW81uvR0w5wuIPY3rd81QCgBNXyPBAwytAr6
0F4+7hQq6V2FJ0nni/OwxcWygCilQI+DgfiAo6+njEX8j4if/lXE5QDm7sCZPPejzOFmMUcFtmnO
PXypOHAH5h9krRH7FgQzGZ+I5RvCbKY+fJjVlhKnml6JPtZC/4+H1Osd5QJGRrb/mM/zq8BhJRg7
IezUwVSFTE+3StS+/BqeHWSnqqKFCUuY1zDwsifdzQ42FS1tjfCh/P8rVyl9hkjZDAXQBFvC/2y1
psGaJBSciERV7bAUvOTfDUn111mEghsfGvzyLr/zziutao6YRYQIhXnweKTwdEZI4wB5OD8lCj4Q
9oOYTebY5Kbr7YESxN/Ui9/j/dCwv9yP6yuW1+vyk2nRUVupyCPOj3QH66bKFBgyhmHresbMDLyA
3cbe18R51Uegii9SNxqF4CkZPpCe8ZQnxCAQBzdwSXIIxlL9R3wgtkgjdbnPhslrzm3k5amxZpfd
MLXqWEyFE00hUV+WCSDswpU9o76TuiQyZJOBizEiWnTk6oTC6nLcrM69oiP+jI2U7XlJpbcyuHX/
we/v/un8lQBJEgmIk/PCna+BJIwOwbvKNGuGgD7rOb7SOMbravJfgAcW9Qdc2mYRKQmSFoqjtdnH
zMuuiMQUps7lNtkMDMFfOXsdod9izbTvL14Fk15QtRNDRuDu+D2cxaIxbuoEVitxZElxotuYTsqS
aaQhO9k7wwBxcM7T6gxOeOSgq4goQXDs5TU3nwgFdDBhDHktzQLlCpa95pCXkYRIfb7h3P00EmNh
ztRaDUbuWEp/L3gyYOfraTLuXez8VwpdJmgqhUQ8RyMg8JgPMKlGdVUPIdA9FE9b/ADdBujdGk8I
E3uTC0QtnmeIExlRolTTfagTAEmWXDYtbQkiAc0ln5p2PItokAyCiTKeQlbc/jvdyUEaut2sWaPb
h6N8SSHO3jmQoz/J+atCQ+EbjPkWZC8XxVlbfTE1nMYPyeEHK4fa0SKzKXOnqeZ/N2zd5WISfRM6
eHwVEFG4LxQfle6uVLDUam+QxAnEGRiy4g76qaQt0tFQ4uvU8CsPrp7jVfEZFqc39tCzmkitf8qN
oxL0+lr+cNkT+4UVcWV6QOghn+yO03m39hj48x2oSK+o7ySD4yxnJALGzXRUeL1DDUHTcAsmjkA2
8lo81gLq807t3x+rdkXKZEmS+PjmtddGwdNAlFY2LBKTJSM0seCjeOAF/eNKdwkeP+X6gYtkSK+t
V54HcOR4DmjeH53AEdJms/7hvaH4fzpGWO/YobYQ38afST4dVarXz/qtZQQIFC6FmZan7UinosD4
8tCuhHhNyAOvr3eYu2wYIWGXvoyYBXkd7JfPBvM2ZkVI2LekG81O85daZYPax9uPUTb1hORP2vBb
Tl7T51xoLqRKm9AzSmsYcZgdVqUc04toDWxumehPfstR0QeSqXZc7xpl4b9Sadzv9ygB0ezBq8Zg
X4rbUVHkqA1yPG6clvU5gIBkJfZEfbzc523USJrODEdZ774YF79YVzEMkXASGt+tYeD24yy4jf27
hgb1PYhqJMP2aGrZoiCzjzyQkYTiPFDXbHfLh3wkYxcBLV280e2/vEVvSbRmU6onACQ+Jl0tG9z5
uUDy6sA9NMNzTDYl+Rr5DVfuczIVECtQMWTUZM2KJfkI0rDqP0jMv1MEufIRoIig6p8P32R/d9Tm
lxN+eJWY4IifUNpcElb14npGnE8428NEkWlDju0YagDz+DWun2dinEC1JZ6wcCMPyC56BR2xioBm
C1+8KsNA5HzW55IIViPDcJRT6jrQZAG4mrlrfOYqpzCpjzmpBPH8CbntFAZSSYG7IgKCMWQ9Q9Vz
dV0TKaLJHFWCnqnbNCM6RInhjSJpqbXz4aNSux+aKbMiF+bkcudjW1MEmCo31RqtjKQy3vFQIiz5
kOHnvHRtzam5ZCPTQGJdpGANZ7ZIpZUVONacPjZlFI5ZjlJyuF7h5Mborp/kLmGvo00bpe4XktHm
JLNdqJeaNxY7xpY4fc1uMPrODuQ9Hqrjd42r3w8iaubVKg5cV/hSXMg9z+uoxXP04E/Q88iW47Bk
SUL8RVL7Je4pByhpR4PgwA1RvfKBVlAPQW2r3dbIonwr58UOtpB5oyyYhFi8FC5Hn5v4y1dRMkF+
gg9cGyWMLCEMo4pK3RqaH9mxSB4/FUCjRdgRzBiTXXnI0PQSgSRV7qEF2yxyGOlJV0KkMzWGydIt
olTIZzy229oX7Gp+3s7kImWqJnEhW9u/qEOGwOdf89jjyQn/spI6HskAiD8JsBGHrXpj9WkdtRrD
B66IkoAE+wQEVj/IHuYE2BgQ+ga90m8lO/KQTZQN/WAPHVPKwMJ7+QKmGCyN9Jy2MLWhyWoY/ZXB
fBgjHM0loAzmPY3GqpodUGT3GwTvVrJieIVhxdRq+NP/Y6/4isRaYHscVzB4gN7xrQPjOMON8Pqb
gQvhYARcSg0n7hEKaemPQI1fIx8fkOUS4w4+mHT1rX5YiM+ZfEJuY73He6k9OD66yHv90nkZUkx5
9ZTxBKOm9btPVNHINjxXsXaHV++z8sZYxqgojINeh95GqcbLjk6cB26xnWaw8Mu8rF9CkKVvHV6z
psO44FY+pBqxtj8QZn8AUgztSHYUW9r+ceF4io9Oi0Tjpjxu562UOQ82Q2Va2BewgcrCNReoSs7U
7rm5z1iV30QeVEQQdpMwOv0W1RvsE6wGDBOxkDSLxJzVAFyFmY/+EXh4cHNkb7AllHn9pGohbhkM
dMb6Ny17TQOy+dH+5yDZ40XPBNzLEZft18OU/twiRS+av6lVlZVSDgePzYftvlOd5L7jz8ihBPN4
/Z9lw6tF+NRKiew8IXnGYtRTWcCtNmYj0H0FVBprSetA4ek/F7AwOLksGQZuUlVYiLG7ZCy1Lrpg
h/dmn/TCmd1P9zaT6hQR1dm4RhnN0GydDXP6hGHS7uGTeruugU5PKUcXo4l8aoo8wGZhhTxTEQz5
c9CYKi+TEO+ivq54yhea7sCq1tnwuT2jHzzxfJb2dB4fzJQjX8liKTfB04aYMZUEP774Ty1F8wjW
RjqVXH8JAgHeAzN6Kp9XD1l4eSWnQZ0BMaEwYHqdOAu98YuXMu/BB+tYyVFSMGiISUnJs07m0i8g
P/GLCYlXaGEG0fgbqI8OJzT0vzb5idU2ZfEKH4ThnHsXs8mstDy0OX+j6no+/rWfYQ3I7BDYtht8
g8CT4fUqNmLvsFgZAeGMpP9x07okynSYC/sUMgDduCGz9unzkQw+eMo1aUcr1VlSbIUxtWcIoMy3
W1VC+VZuovqEW2Oae0LMIfeefruJglD9xk2wM0fmCdls8I1Br8dC2AAMdPdaw7A0JTTcj/K/VHIf
E6kwcbMmH1VsU0M69eCsjqAQ5N30GugXEqEFEEmeZ92oKrWG1A0IWHNK23GkFXwKXgxkrMfbwbyk
kOos3BzO92yPRvL1TZF1ln6i9/2MKKaXUaLaYaaRFxVJR+a544uTsDM/zT10M4kJlXwn9uRRaEyT
+4R/9WVMzEtmxN/zfZoYfneEBd3G4xgqHXD43BBzN76/A/Ker0B+D6BNyWixHcGKkA6ZIE4bm9ly
FwBSj+49i9b/vaidc8McHici9h7vIsSiPJSqiB1E2AZWev+7rMWph8A0HkyNPKDswi9JqBNAc2Xl
bBWbHRupmcXRgd0X1a0JfjsNFxW83zGmUOOsheWLO5Ug9nhUbgOL6bnXW0gmmQCEwLoEaEN6hrFs
PUlponwiXHLZKDx0Xm/lQPuj6+HRXW9G6aqje9mPEnLN6qT2CdWwmR6uQ8/qQHvx6riuH2Td9X96
G2Q8I32wCh9dSW7Sd3/clgbKLkPTbOp9prkqmpW2hJr/BBpSp8XjFTi5O7u+Ipu6gNgOvPoa1acF
HACJH+tQ7wHp+NXPXEGnjhf3zIYLVkR7Ge0P7iBQ5DMbzqRVY9ZiDU6L6adSJR0QtW7MSZB5s/tH
YbG6Z3fIsNfEtoYXrV8TZ2zh3JQvP+pnVZLAb6BS4Ds4nByoMzzSDsFdtXIVeA8IREGTQkoeoZu3
bEezR7wTNgwdRKNytZYhF85aohWh8JeO2F3xG11kIKQoklB5WC3iBUX9W68yNs1iBwA/a+4hX7yQ
lZAfnMSy4oLT+4NSxKb7KJFR3Xb9yuZDN2xXXliqppG3AO4lyvQVpilguj0QgemuoZxXiL7l1ZPD
Yi9GQA3WiOwM+ua7afm8QPKHp19keyJ1PiZDiXwJmDKRK3B+LVIwdNyd528YiKWNZDkefwrssFHr
aCZHWNCDRsSAYsKG51rL+zpaGUXo5OZge9UGtcokD6NJQdMUOSYzEgSvNz3up75NKtYYUt3By++F
HYJmYNdix3DSLzfvuy7BXNjJjbSLO0kjwNChZ96MC2Hp588Ag80GC8+m3ncr65dmgQI+JnmiSVNi
FmmIXpKbrxMxaOPn8vHQTBLvrUo5tLGF/JWm7oqiB0v9X7v0qZux5aRM25XKze0ZIwg9jAHUyBUT
nHb3JbozfcZUXxo+qXo7vU3JD9ThK8wIAHI9sJdKYt8XcgYfxtNuJ6nq7/7BBs/8p0e/DPYRMHZX
JYskkGo1qD9TEMXtPG4nmHsCMGaO0wOpfJZkEMIb72E4dvlyjURzMZ2Qy18yOohc5k7daqt9AMFj
BrJ3nua6+FTirrIEe+kS1nhP5FM64ynL0Gr/CP/CPxexSyBfhsmK8siAMUZqVuxRA4HH8LGHovs0
U9WqumJauwZc2uzr7bLBjVk2LcGeXd300MgIi2czpY0jHvyBHbhK5AYXTZolxL81NvTAZHvxzC9g
csR1t1KOSsNmECXES5UpDzcbPQuKci16XRGSuTJ/N+IiMHh127aNpkXlPMUrNf0n5gWwdpSeD0ch
9t2wRxpP2DL/IGvPGIiy3AoYVv9ut00bcwsKI8YkLfbvZwgxgof2ifwyhyfA81KOvXxjODtrXIZ0
fOF86aI+KKY7pfK0hpnn8L4niXcbOsBf9Do7sncGiUQUAX9RivcVeIhYbPoEI9rj0GsFzCl4rPFx
Ia6Nf8VcAoDRe5lJgeKWJyq7dBtN9mxHyRbgjKUQcpODQYCys9sbdU859MeLXCEKtkHFJvpVgw98
eWbHsIIcdp+GqhS9jAWd/7wPYSbG/gwyK6kMKZu0Iipx8z/HfGZDvK6vb6xbm59WyfXwJ1FcH30H
g2kyXy0TyM3ypBHo18mj7un6T6rgoOMnskpoJd0VSuxesUS3ZygzixQrq5d3czxEgrIBow6vU+Ig
QxlmnqaxyqfoZdniv3nhqU1vY08jcsKAXGmrmMeDXf1W/b/Y8BjQAmopLFMWFApF3mZ6/N3vgElb
uWMM+HtyqkI/qVlcYC8BTrNyA61bgIaqaqFa4EZKPwE/FLWEgCthnDlfJ2Hqi0Wnk47HBa8r7WKA
pavrKYVzm9mlLjADdFqiNJ4paa9MtRY+AmOzwlj/NmRRd134BW+lbjKEWloufpBK2SSJo9wbuGSp
eNqVJLxLEQpyYgTjzNhSiAObJMyyppHuYqd4rCcVAOx56B6HxO/hfAG+hdCd5MV90tglSu5VRDm/
Y8w+8CEZrbg4+evbOUovJxjsOE8SrK4fJdclX1TtuKtXqukOK3U+hpkLi18RAn0bQFQnGZvBLwOV
NB8x1xAo8a1ZcgVNCuyaB03fq52adp4tf0pJlXriuMmXfl+noKeSCs8TUu4P6JkKecyCsRoJtD6B
lVKSLadhUP9SBvi75NWnPM9vOKyHrIlTO2NWDJdk13PVLrtZPC7lRnu5xCr8o39aWg5eQkFhV5ic
jnDTfmnuPWqkNdee0d/Gwek2UUXG3Kul/UNrQCVrMZ4N7SbH51b5q9JFpABRpjf9qkjlSKOzj0Ij
cZGRzgM+nQLynm3uWRO9KZuwHKolyk0bqLV6KBCxIn/64nIK8Bp4quuSuCP+86J0r4scZr2JIVmn
x6SlhhD638NWmqdX41Gn4I9EyaD8oWQYqtc4WKapE1hDYfamT5C+QHsmIfNKcqyEGGxSefdr1HZW
IoD2i94r7dXTbHJ3U6b6cMGJrZWrvubzYWzhX3b5TlBbuXZ3AWJPkUqv546a3GvyjT0Bag5jpwYv
4dmwaRoLtSSOSZYGJGsdBnxbVtR0q59Clq/0TvijoRfkRBUKr0zCV2gDYla/OzBgoWa7V/Ba3Zdb
ZmdeK/MpAKMHtJ1chJbtDn28pM29CgDirb0+zUqlicGmWLfGK8ZvIPa+gyIsmkQ3OjwlvqMfYErY
CAM8Ov+3K2nqRzOW+wPSCX7FloYS6hDizKb4zSHhRgOmag/qJeJmwLrWfarYJAcBCFwhN8Lah+6v
TYz3s5TKQs8Fdiwk5ymlTKpuZ/2BUGVquomqXzt4FzE9hv+3jrMxUmG2tmJg9mSquzdGJVeCOgng
NwK+aPyfFQUhRvVW+WUI+f6LiWSuLhOXx6Lql+266iT4mav2QWJ50L4xILffYR/G2/Tv0qTT6Af1
oWTc3RdykI3HSeBRDyelr2yVSSXpBLgNo4c9h9XDT+FLiZMEZZCMgCLvmEZ4XDRunwPhlsm0eF21
W0SVFMtqGc6PwIwR1Csl2fNOMJzvYhK0O75hu0QkxE5wul+VGN515h9OxDYmflhWvVndfwWBDIDU
SbsBnhnZV3YLt+20XHlQ+tbnL7M/d3EAogqyfop9EyWdT8wY0CiJZEC31dV9dhxVISEIqKCPN6QP
5Z5LDzBUljR87sOnLdPiL9XFmR0DvC8v3AnaznD+UoI9eQjStgvAaEMrGsV3b7JQLT5113y0VMLP
qxU8mKIelKSp5jE1yI3AGu3Ep2t0Lw0RsBQ3soJBvOW0eZYrMm+chSNPmNSVeH4er42jFuZG9b8C
j4kvRXi8TmUtCw3Yln3yC7Nvku4sQGZZjCE2CpRCZzfNG7135qvizW3dmNj2vnag9H6Qmllsn5gX
9tMcTlQ3cBm0bBSr0e1wU2XVH8hbQWRW7CQ6YWGgd0pp7o05f6Mbq8Ahocmetnn5SsH4a5b/uzgi
eXrZBZvk6v2QJeqAaYe+TW5beqHrHHMUmOVIdtA6fyuS5W1yt+8JN5n6Kh6s7zH/CMq0AYVf29Bq
jXsELpVyBSmd38IaYUghI29CmFpJ+HFw25Yik7h2pRnnwxhj5wC2tsvQDrjlJvap+df/ESNlrAUX
Bz8NN8pduzCp9lj7m9xOJbmc6QHFjbrt94aGa+mz6qc0O0rCCLj9RZF2X4n1vg5L1M1XMpmRsiR7
tXGJ2trerCtg9uIPJce+9jMOsaSRNeEKe+PzeHeXNZMpsP8UimDvh+fSAW02/GzH8/zHajpf8yGR
g7fmfAMPl2qcZN3MBufyh8/44OJxJ6oEDc/T46c1MqI8MPWCLOo+YBvW70E07JY+QdmEAESXfXw4
UZvx2W+Nn0AD1Fhg3z+e2cBw8qza6f9vQVPiZP+Rmd8nWtyKVRb87FqDVEWeuWqBqAls/AEDKdtg
2JSwdKGpbN710GS0c3jVFjCIlVRzFz3+a/7AcOsK9iW4gzDcuDL0jNhbyA4nnzSk3A88QU4npo3e
n/jg6Z3mU3NkXoDYNaZHrWQxY237NdTrOi4pFk2Tz/eXaLJg1RQXso58GN1UESUSVjYqWqod193L
wEmEsAAhsmH0sDdLH6kANuJdC11vRQlC3w9OxTR8OoVy8XtWpuOrXKqrISxrJWtw84FOX9kw1e7d
cgOb2Mzs0SIgQ6YbpELZsv+1gbuzXxNyXfh2oZUefwD49XqJfIgHFlp4/plC4oGLrkXTRMLjEjqM
whJcoYAtcFrzXwXgFkMiPm/7jgxJvZ2cBnCrAYnbo9XI5JQktvyE2LkX6fCGOUwyBC2vl3c7VFRy
1nt1kpG4s6KNoWrNvcB7N9zF/W3wlFLslvNG0nuplZwOqvlqqFsGTp/1Q0iXkHnhLBV3KpqacqLa
SkNHyBUfJJqPbTzg3/Rju/0+I6fNshcu+mPg/aUK8RH0w8RvZ78vLIV/YEGloOYoCxhdgqwpBpHU
JcDv6PpYCeraHTZ4mJVfbe9aY9d0hKRJ6xEPqK6HJkTbIGCnlCzMSCwGijbOMXFM2hWG0XgYay3a
eIGdxW3poxlICPKa/Qu01gfMyO6cmSMjHy/S9SicHQDraI6MF/9kJjrirIbckYo7tGQmZ5tc3Poc
aRFmg6Ltc57WUQlUrwMYZrEicqq5IKzuolaDNjjyRxZ1st4ZNRw6kRgVyESV3G03exqkxke9cjpm
zE8zyz9jCyhHpKS252ZPPRgQb8KEoq7IKwUmCxzf8A0ae6/cp4cHnr+TGNAVhFf1BnBQcb34ma3F
wuDRMzoXbJttMmDgnNI6WsNSb38XZ5lTo2/P4tKZzOGL6Al/1RcWbvxjVXm4ajH6muvZy6ECFCHR
XmYLWLQq1YgVQh+fhvRIvtYBXL2w1/7Eg6qFTanxkDZA2v6e4skJ5VbUMl6NulLsRA9+1Ih9t+Po
ptIuKseBTs1WHUyzns2/tTdiGV85Xdoe/IwvVcEDsI4TMJ2v8QWTCED9xlAxMRVFGIwT7f/bVt1P
qiQ9lPV6QTgrOUoAwq79ToXbntwLz6xg6fpyuSd5J/pbamkojL1mT6uykohLBTwe4IMOBOHkODrn
nJkoy1zJiYGBONM8ChlHOSBk3ewD+eQLVp7PhjnaRdveU8WxqreqeI1pZECSSwNRgLC6DSwi9jd0
vVwomJoCrv0CgKrJMe4urTjvXRafmzhRW0RxIxvvO0ZbV3Bf7TqtUsaK2uUAtgBS7Mv6NoeuAeBU
jqgAekPWQ7GDA7SnA1GjneuJLDCbqu51E1pbvnSmxZiZP1DGexO7cd6JYzwq/UegXLqnz/HS+i5n
o2Td3JbMWvVHniGJ9SWa5zgRpR2qH1mbzVgWIAYkIFhJTmTDuNio/jSkkEawcdb0FmJAQc1bfBYc
/Cgb0X9X6bzIEjCMYBM3/q69K9xcJ+DJEfH38po7x/h/A03GJBRMx7nMWAE0/ZbSmn9SqMhh2ecU
KJJBpFpojKQJVyagjHYEdnW9EcOg2f2T4NsfPZ9qvQmTRQ1fFuYL338ssTdxo4CHr+fRzaZjUOXZ
Q6PGIWW8vjZ7HrN/Nr6lr/BcDiUZKrUivCx8VX53e0h2g5n0LhqF4wwBzWp+utvfSD8NKM+vSk6e
DcHGZ3y4vc1IRYHJeupJ7aHcHflWA9OU77kBpoufCKVsC2Gvo2uRygWAKqGgzbk6tzrfbqVAFXqM
luXI4Xll1qhlnGf8n8zbEBseUQyh0rU4kRqQQLvoMY38PNY+ajIGnErU/yTQy95MgqyeluUP9Mu0
OGnKkak35uquyOhXa4FB6FpXD9EkhQtIkx5PFdk38PjeLkLOrNwopLFXFE78cCvGsmTCy2S3itel
FjRRt+ZUSzp1MOee0QE0QqWjgKII2e5fG9JBZv3gYIiGRW4a4jOu9OEMV7nWBxsNRgWiLY9znq5X
RLIgIMkdCzE9E5u4v6iBtKTohAEZ1qa8fvQeAGnkHft0slazKj50N+2ajeMmFyG5C8crzYwJeZkC
bJf1uV5llULpMxMYkJ80UaMy4B00Qy+ErC/oY90Dz6IZY/qTTF3Un+eueZ9vNQmF9UYSqlZVIqaq
x0sZvVkydhQnYwnqIeqV4tKYFfUPQbXGyb5/fcGO4kn1QQWMtTuwPrnB5UruzdBBUGNMlsdn+TR1
MVt6sBxdhI0+N74lipGrhCdAcH9aXpaoW9n5sxDJJvQ1iqy8GSUFd2JoclESoLGmePFNLnZDyb/O
GYLWVjOy6XVIGkQNCHa6OH2JCy6G4+Bm50Zk3LGEPu9ae+5c0LG3DdaRfLqerM6uXuqxQ/c2pHvG
vlSM59/xDv75/0eNOy8lGBggw0J6UJkCWh7lOsqpOpzCdVilbjqkZj36FILouzhTrprNuA5TlE5N
XF++RSTqkbNGNWisarPNTI/RLLaSOLhHyvoo/iVWva9auL+3U3OJSwCbbG5g1M/hjCD/33NP0eBE
ptLmimOC1kCDEH3QJetcyf2hBeCcmguZ6nnn+HMqHkoBEQ4xWGegNZpgxQrli7ubSdmkXPJ6+r1e
uV80TrRQXnpLamEsQcehY8i/rZ7SRHLq6wI4Io8kqbfGUJMwYhu+qMavyekjovhaWguM8HL2O5AS
49JOOFpnstCleWYd4Fu6oDwOe8hZJC5FE1vA9IVmqBX1TrDvXtNRWyGGoAtvPTaj1kOlC2WysqCV
Wop8i25gXJ3jKOOCTHuKUBBbItsqSZ+qWfF/1pU0ii0Zn/tmR3az7nuKHMUPcS5VLfvTfFBy5P/l
qK3JYvZiaXDSoLiXT572zciiYRVlpYXSk+Ah+wLrEP3UDQ4245yZMBiVuBeHk06s8jiz4auvSu4l
6GRlCyGL+nAxU/cRzQZDbVDjwPDCyyidycVOB7hs7oHTK+vdzUcHjyEN5fgw9EUaAbyT7sxnUVYc
mAEz7+yOdj3LNiEvv7dJdskZWdIZs9lpZGLSEKXfp5KP/EhT8FIeh5m3NWoOPAj4ynEEwLMf2M1z
zIxfHW5NRQ7lOmWgmKmgTgj3XT2MrzH+ozcsyvlOBzobxcnM5AVlPLfDAuSV6J/7Xo8SdszMlyjU
3ZuphYpxOM11TSk+mv80pazlgDl+/3dnCvRD3BzjwGWiS5OC+vv5cx6od1Sl8UlsnYdx7kyUyPnS
P9NWMDAnSIFiYaQgWEiwH58yWjZufWNoIrzJns11ja9fmCBjwbAW2bmUP+P6F3hS1+wsNz5M5mtu
lnqIrY79cFFrWkFYbjI+9J1+vKXAxfhyCh/nhh1cyAx3i42oKrjt9qXqN0pwTTe8cAuhKriyK/Q+
d0dO/2yWQLZgbsJ7pELvx2KHHIZiFMG6hsD/vttx7s6mNyDXoBCdDMqPlsR1oO57/ohBrRxYz84g
26f6+VxhHA9BmxGhaRrx3qFO6NtFKMDkKgwLWHgKh05Hpy6igdGHMfJsMQUAGonxp3uuJSA+uguQ
N+Z1oTmcWrqQtRG6VDr6Ko1+UJ6bcBTVPHJXZjDJm2jlWvMdXay7it9CtmlySsowBq9zU7Iqf1/7
VeLtPUgQswSxHelK6pXbqgvOoJgd1zPEkLWoIPcPgfx5iEm3OtN5B95rnueEoMOoFaenx7X9hruz
Q8Mgxq7v4yvhNMuJAGgvBAkYuPiIYIL4UTtcu4QBzwxCS67/nVgbTera/BXsGhSPpmJJ+RgKblRZ
4syeMYTmN2NoyGW2n+IjDjdn8Cw+fRGxjEXsapQZt+oBS55jf0VIAjO/zZ3BuESf/X1/9jg6Lfdf
Z6N3FgxHSCtTdrjUghPdRK4xCDQ46ToZsWU+Gih0bGVHTMiXxLsscU05lzZ67AFNweOHn6HU6xkn
OHD3609d/SBoOKAXGYTe1mhNqCg7voVuRP+3bNm8PkFweX5HlbHhs35WmPJmAuedV3/5O7krb8S0
jqtM1dZedu+genQxgrTG6sFGrk2SFhWFu5VJ7Xvj7kXp6hktGqhaYJVDRhdH4MTtrP4yXwseWqpm
5KYIjymBKCH0tqm3hZcO2Ycn0VgCwLBZrWBqlSauJKqW68wiPadYl7Fr5BRIRIL/cEqsD/moM7Ig
UVO/EK+Et6x3Q/cf3fI42cIXLtp3DdEduSSHhT02aJor6rJ8voftBxdJKW20G25PjbJO5aYekw6C
8f4Qytkse6pjlXz6+yDl65vUP55VnG0QlSUnZwn975fDVsqXqatzhA5geJeh0MQM1qi358UJMteo
gguZak+xGM638DxeNfE+OUa20bK1Is3kNmBZCT1PnQOVD9IqpVDpDaoQ0HhVkXWKgLEpeVOAuMBY
W3JTZOplFeSSChVo45u8oSgOiKlRX7ZVCE6fqnTPtsb5jOrWKmhjBVNH+cNilDEKwZAbWTcpsHr4
z/ReAebO7pdjhfgv+KF1zSOYnGrfZuok/zfA1TKJEcWdzGJMyl4zRT2Q+rRbcI5m7n7LLo/dH9uw
5FRXiOTBAqpnkhiSZBTfv/4tsWXjXu5gdGML/Bd7lvBmxsGACIRWjy76ObPTXoBrJjYwA7anw19G
U0NOTzsIt8ULtEbS/PuIAGEDZU3oPcSLnd0CFRbOUoN/0stSyGjin/XXizBcsrZrY5YZKZNdHnba
/K4J+RByYlXJyxeQNquBL66yX4IjTBzhP9ENpXEMXxqNEiG9CGIvCLbwI5nWsEETWvRd+Uzwzg9G
7du7BTBxRrJXkQ+/zQnNDmQujq+e5azsQ8TctUiWz1bdNd2HarLN9j8zc9SKks2FhGVn3VCSmdCM
OhHq40nwCjpxIhPoDsDpTtLmlIX9+fAOA94Y4u20oh29X/G54Ky3aIODVdplrIhC+9mcVoF3jolj
I9mmsH5FoGz+gocUt3cho10PD1YYnhDCBdxTuQ30YM/WzMXEND0kUJnJyrm3LX714iv6ME/PRTkW
YP8hLVD6xq05t3FnJo3gCZb3JZWGmEeAKAuFKop+O+/u636y/PvmWeGx3f6FuecdHyR9nK9k66g8
McIjai44sfKBJ+wMTbwyGpsH4FHuTe+G20sTBc8340MyU5SqW3Yu6TkHZlnPL5Ln98qmgZBli4jD
7R6oCkEEGF6tdMT+SgnuzryHKonIWQSEE4YZ4U40lUkG4eKgfnQUJSnhq7W3sWP9OWV+lKr+PhHm
zKNmfnP0NHID6drc1dFHIH9HVB9lquMBbBMlGalvMt9HPlAnMU2I9A9eQB3QkCsvAf93ktt2kZju
SvgPz73pMXJYOJc6Fi785BThZB4ihrclwB3xG18JzQTaLVuZpGmV9i9G02X/uHZttyersHS6e3af
aH5W4+oJB7OG4bjL1TmlMtcRgzzhVzL5VYHZYmltT8zK2Bnyd6ra2ZncZ5fiqgzPqymXrqYOZAor
mpBJ8E/p580CpaW8Z+b1sI+8P1y2P0OOrgxX+x4CfU/abc+wBbmNXMaIm/cLztwWGw9MGBjM/ncd
FrzXbtTjaXnzcqmfe9pJq5OA2KJqQzXo5T5MuPrU88UDJcAI3vlCD1wqeLTvHP7yewWR78sCZ0de
9EfP960XZ7QXWojqV1om+lCI8xK+5h1YmF8nIrP9vmI8gXvecvogoFABs07KG5jC81wLUr7sJ/dh
OBLhcvy6XrqDzrR0VsWCfVE1dD/RUcijHsnKvqh96y1cxZJuKJZQYRcS6ZU0RRM6/rw7o+NogOv0
KuayCtS+ak1t8+aSX8SHovKztIryU3qjG6R+YyH85GfKzVssXigy6sAfUk1hh10lK4Nx1OD7Jgok
GT01GgHUJ0KiMkNFnzIm59Xrq3ybtz+zr+FCIwycr9kmKn8tH8HGJQmZdQeUg1YRT5Ri0lD5TLSM
GsvDcCUvSos4Pk4AT7bZYiHvl49Gsj5z4PrvLX2AQAtSONJflk4IWn1d7uNxkWCnXyL54KGg6Axa
L9s8bqoglJMou4eODjdBpUG+HWpxGlhSqar3k0r7KmT5Kt9QzmcWZrkgu3LIre8H+dV36dtA0JKX
SmYzNEMFDkygJsbIlstrPT1gcJh7Y4oMUkg4eCXCaJIAryL8tUk7ZwcLVp9w64C3DrLUvy8Rdfvh
vhC/7HCm/rKO2v6yW0eaf1QomKwAI9ORVxSArpRYcAj0Tz5jsCp84oOk3kxAKd5rxIPPZ2WSU9Xl
4IP1eAtyA+EhnthiINurcNstkwpmHO+B4FIYhjU6Q0YFQP92bSjxMGHLi3c08zbaWodoxta1URX0
ES9yPx1mVv4obF/FG7Ag8GpPyz84QqBluRgVFA7Y2xfSUshetqZfCVnexv3y3Fkb6SutTqyxMjtB
XQOnu5j53xhfSw3S++MY1KmM9L9DwsXWSKPLc1ycGk2MpuQCi4gg9DxLzWMnk0e4aqCN1Js/dSdy
HKtoObPwn8ramCKGZIWM9dcMpLjVlPeLWALrSfDyX393VNgzqO8bv4lEtVsaZjEfLe3g0CNmy6aX
59mm1liTrQ4SKaru7PVJWV6ubX7GD+Az2tS3sRRmVsPiLk8frcSN3vrDOTAFUVvjQDEWBA2t0WWN
BhlXGPZCWCf4BIxQVJj69hJkdmSOI0NPrhsXf+VCswd7Rw40xq6/C2zgD0QmO06MEWcLMRw0ueoI
1ElMfSo1i0ZNE3Mb7wF2JcLez1rWvtbBpgsd23Uuv6dfrgXL1ET4VH+0Cs3IQhqRM+FDSSAqu/nA
X7QTf7OyxSOpvf0Q0M197QnvzcopJbp5PAXU8Nzm556FFN2ej2lFGeL2FgHmW41x4amKIiYCOm9o
qkZnT7mSdppIJrmlhmke2+1RKp7l8co8AudwsLcF4x0vFbvT62znjR/tAnYXTN4rvqFczaZS4niB
VTghnlrvDKE628cWy786oAlI8nX6ZCt29uaxOHmsXopWD1J0Umz/QE5tomdcVcG9f82mk+rkGCin
oUa05AozMzz8thBbqVBjMXPMxoJxYCksWFxSFOmQGZ3kFdZEjERkmy+GmzgT+nvaxfuvaEkXbk1l
KnGFhNYalhdGmzALO/FIDhNoYEpkxyvz2Vfo2pJ/Gc7wGPZ7NEUTLIlJwzJZ9VRlZTnZnowXdQEg
ss/Oh2GnvwIPVECU38Y2f1CYDDoy4jVX/mSCxKqSq2b9SIdQNGLfAGrgRhtytzqrEiSeftqs3F+P
rsyh9K0UaeifckZjtqvncHPIP74OWUsUwBj/y6ggSejoiX6+qCKOjRFlARbpNA09F03RPxmEvFqp
Be2/9SFbr2AI3qlswSBVrBoFaX5xHDEWzs6wNev9fVAwy9L8+tvpnU0SCln9iQvSsIfRJ8fvpGuZ
hhNJQSUB59KnwGWdh5QLYBCPJ/DgB42cHAeIST84DMzmLeZN3lfQBns6aCVilgBIW9OR3Q8+Sluz
fE8ZQhDN4DwBa8t3gCq58fCi5Vx2UX8LhjfZEKR6ihRw/bnj1eb1qqOX0+z4qfiDfnEPY69Ywch3
iIMPQghMhKzEFxWQ9hRfUs7KKJIwmOsB5DbTIl+sN/NnGpOoZh+KYgNRYM59MrYFRLg+o9M+iLrF
A5P7g3IzyVp0fbCvJ5G4Dh1p/31usfNgQmeDWdkcHh7SNIKmvgZJ+PrpUroVs5eoKzALk7IPHCJ8
go8JJayeZcjd9HyAI/eYKRn0q520RRwSSreGOlsaqMfCjVglxO0HnbEYPSUea/oqZ+zI45r3ZZws
P6s8uaZDhn1Vwd+eBF3Bux7XwDDtf99b7Z/UIDanVrrCylRnne1PbmdBiAQh6l91cHrAMFSW32CA
rGk3H4hFJ1y+CKNzq3U+MO0Pm1j/MCtsFxbDNYP+PuC2K6yTLVSLjoZUVARv0VuCT507+0s9Ewkq
/S0VsmxcsuDPCM4M3W+C7SfCb4TRXNEJO6TWiPgSGivnsJVfwCBX2MA3PKnh5DxhXZWEV9cRcfQ4
+tc69h7yzqxNNWOBT9GmTv9wmlFwCQx19epKjP3yEQkEzkPteyJgMfZfdUQ+FRWA/YbjTVMuXBO4
LF5ozrkgLyaVKexicV2RO+K4YbbqQzkrYh4v6YlRnMSWuSWNeHmTQvsw9zI1AAR7N/4Ab2fkF6jO
F51z7L+gU2SVzv8QmO3JEziMBg0Zmm57Jg+hqSNRbqKPkkyIHfb6tFYKMuMiDZlK+0YvrAJAS+kg
qzwb8+SfkRNZ3iKoCR79U3lGob3KVueebdo0Bdnt+1WBXX1F9CxaN53CDa7pfDUQ+Sk0uTVfzWhl
VuLqKNuwAiGazU3kM2Li+y3uP446crMQFmUQP/XngOz8ZUksU3OcBF6XPBa8sQcppi2I51hG9ZHn
iY/sBGoZIDNSddvykxLftaipUb4VEZBXerC7/SdY3m7z4wN1Hz7xDNPozjzxW6UFXkk/Tn0E9Q1l
vcDrYsSMN8mNHktPavjlfmldcfdpHkEh9Hj5Ic7ugxNdKvpy3P5jNuhNmDpsqgJtWrNWcCKWiXQb
9gQRm6QQY7W15Mw60r+8TDjZh/oSvyINyFGJJUzko8+e6qD5T+iqvWFlSlYTJzdGALZB7zmxHn3w
Ik7V6/AHoflwKQAYCDRgZq1Pmjrx7Bl7qUj0VDEzyXZo2F6XD65K1dlArdYqvcYscrVbmuLaDn5a
QqVQX4i2a4sa4ti7KhgMqMsbxTqawOti/dUlbFBMnyLgop5yC0FU3dr+Xr1+QqDfO3f2ELDFewMC
SDTqq2F28uYoab7hLL/ZaHQvgvjUs8U4DpkMS4UO3n+LNcs80vnB3QeFxAl4GhwYRI/PxmIWsb6P
E6GaXOyVHSpKH4+fYjWbtG7c0U81Q63GGFrwQh/teLbpb0swqE++nn4MboBkzS2fWxKLwZ6pdC0s
FT2Gr4Wafz0XUrcVSF7GC4G2G2VaEJ2+7hPdofoKZqQYR0cwfRLwYbcA/1rPrBWxdHFD8BqeB4M0
TlhMgz1dr4LYJTzYHIZhnUrRCYDrHsfPCvK8Jgi/ORMk9dFu4zeGh5NKIkksOMzuj+y2X8+qvPPn
4ZMgwMbSz4TBJ/7iDcU5/2HM9JyH34OhMMjHJimQsrLHTT8Q9PKvotUeGjXtPsq8a2XUAL/Idk2Z
8m5YzabuDgpwHKq3exvG9qsrho6sMq6p8vMYUF8onWot9S8mgfqGHNg/q4EAMyNo6o6xUT/g1HvG
Vvb16AWEP2fs+ZMSeuSfhOxSgZWvum1hqWw4VmHwCO4xi/qjfk4nXVU7BXyjLIleoPi+8linqTTG
mMLHWRTvCFByL7dij11nym9ALgeMnywOX1XQcwBu0+OO+xn7+cAY+0J8duDjJQySJY8VY6NLOiDy
K21puIhVeIJC7tw+WWGz4RIDW74kdv78wQcl6unSpEUoy8Vt0J7UODslrANcUa6cR4qYiGEnQJLX
xwZDUunqmb0de8W/tjK6IEzJKLMSlXBN3OMoA+uxUfdyKt2FWXAb8Wo9QM0HxBRRDZeWVPTHfXHz
sMBT91LEvCfUBwL8ByIWgoDSlCuq7FQDjrblzDt4uNz3eczNQWGxRFtjuEISasplxoGZmy+rA0k+
m26NhR8el2KGNrhT3V5qci3+HrfVhdlJSQTyeU70qsI1Bk6p7F3FjGffb0PQtoF9Vjup/geQQY1F
D7jUdCdZa7+hgFM1SgEkp6ysov4QetISFQ/rVVIOCRP3LlegSs6gjzLyjXyBa4MLMsxwVwGXQ4rJ
AWAZY9TX0ZYCz57ZDqiKGovc/CQs4RGVPzW9OHgFt4pq4Pxq003IJC/BS2RCUDib8bmuD8hd6nvA
3cmT9WPmi5u0ygCOgTwekWX+epjkpZKqf2+kQdEEjUcVAUfXWmtOFesBwH0Us+6D86vK7aYwkB8c
WDD5f4JFYHOnv9+VOn0watNChJYxJDSkH6M52p2HwXX1HDjHFsxlAbJOfYApg4NfXN27gEVeroiJ
ma3eRL7yXcZnbYr+JIqXzXC1ROClVCD806empKufIIWLH/7sceF9YxY0DGYvyO9YfifZQuLEKD9N
rtCpIEKIwXhg0FXKTwJkrjyEt/9EIkx3EGeEUn7RKvz69Q5YncYDFjRXmeKhhvyNhjm+Ii8266Tz
D9uT2dPCZFlNRiCl2WfuVF33j1QNXWPL4UHSKYSRzgzql5aoo6DNXfc4Ko5a3994UH+JnTeZ/nfe
oe0691nRXroq97F1ld8EnZ95cbVVTr3fOTvBL449nfK3xRc/91H69jiRt8BbmiVW8SJU+Db6uZ+Z
PxSM5gIypjCH7C/5HR8s9xV2RtupyJIDOzGccPiqZ9YXdw3ozl4hDR6jnRDEhnY1/KY7V315cr/w
q69BFXRpwcTk7rga8xGLb8HvDC1liMy/myi7aVe4bcVtGI6DaGc93JJnFXzRxiHNXUBgmJxprIPj
0VFgDdT7r7D/tVLXczeIHskEhEJAzUWTAAEkOyPhVD5HY6tCJwQtWVeEnsucuUnkDvkPfOdfYEbV
NK02XGmQ/7nOEvYZDWMYhlLxDWMRq2Q2TPClTbSwzhDrWvZT4zqV3gBYi6B/DFyWHf/VmDtCbLOV
MArX2oyx7c0KGMCs7uf9Lx8b7a3Gc7Z40eomhBwY3utdZvkH5FKq0dNXXCKkj18Vvg5FrbQQKxLQ
grYHTgbh2IHFq9+jE8dKyCYJIuW1MGUQowCIE81HpagbF0jT4uSPfzb40uel3S3zNvjGpa6EjE29
g3oonQzrCJ7pfbWxAnVMrdHjecSaMalhxiy7hdXfkMOQGjrhGMba50n/KaGwpJ61WxjEcmW52Xmz
q/MOrTbDoVSr+WTaf9DieNx3Vfa31I5o9eQ228KYtv4s42OUqjXo9pgh8JBN7c7bxn3cQhxSUt1d
iXuhtVZmxDmP0cRTJZEYPE5omuNwq3etqseWp6Hgt7X68L6YSssVIfl2HQZlQ8r3OH08ekXZNyKw
7oVcroBtDmcQz3pgM+odGhWFngSV/LUtuVZq2sEoz2pRpsQ6vcHq/shlxr0WMkXy3wnXv7kXUF9/
psicXDDlBGdvpWjS5qUCQRCBJ2C6utyW6YgFLT7JpFdRCwCi6SyVbD886UtGJ9QfeHDRDzbKrEQO
eznGX+wFggDLMlR9gAUlc2kE1rzEAD7trdr0klE+GuGIFmsGHUcL2wIG3vDoNHd92pQnVfFOH66c
tSUngUDPqsL9Bji2xgT2FBrbyqSH7YeeT61Bkkz9v9Uc0YF9LZF26rybBF9TA0UHGSC9Cx+DrgEf
BmS+3zZr/aly4DboccciPhk5sYjBvzWSWgZSTFbvZ2D6Ws8hZ62xq0MK/GIJRR9cswr/WAWWyi3F
II2yRoTRuuvH6j88vAq7LOOpNC1aUFxBSbyWEyiZVrttChAHl7ks9a/7xdZnL752Rnm3LYBfbVw6
ppLgVdZ9gzqLMqEirLbFRmWiuwDm8vy7tTBqN6bw5uSVBFr/vOq9Z8a758Po8u+l0aLmNVbehOAD
VPKCYHLx1OOZUSz2/7pB7enEixmujC2spavMqHhOwDRSvNpMq5eTdaJWpeCfNdwoJ55rwA9ekJmh
Sv15wfj5VSKAG4dhIlMrQ0xlxWv7yAiapGKKumYXiqBZZmbCuzzDosoptGRroT+ibcSPba57Zj46
GZY+ajtGKCglbNS3uNACBTi9Fn2/eKjGqubDXJ4qVFiqRm0ReXXpE7fPdJYpZrRtjTwBUmkskB+u
nl33PiuHK+pidvJEmMSHPezLTyo1K1LG9UFphtsHIAX8EfxiK8/zWreDKhXTafU4uNlB9IO4SgCt
7ZzOJifHU7S75w+lOmsLyeeSkELLmo+y3+R1tYPU4lxUvVao8CA4ynZG6+ISaNqDEkjS/+MFldoq
iVwCaiZwYf02oNNYfbvaHXK41dthH4otEMnzzk5QUDN7a0nhNEl5wJct6tc0XRYg8WpvQPbn5fPB
aOzXmSPVM8SDXEYELp4oQdh1wosJrl4zOmaCvTuFSyvFVvzJkOzEVmvQvEMT1N9jSzm2o+8shEy/
dmcHxLeJOUODkvSZZfsj1sQZfrlMOH7LLiyV9wOiKc7egtCI6XxCivBmgq1vFsexojUyzLlUZ6GE
Unyryj0ccJPjf6l+fDOKO35RW2UO32DzhA6YEJBSLNF3FwvBILfrSBDUdZCMGqqNAiYTwQRPxDvE
S89Zmt7Eb2yr3uprdVbmHPF7iyB3JO/+38/tTuGX5krIe3rZHQBiz68ZwAbXP76NecCYHNFQo7Hb
m47tdOcrDzv4NVGnI2V+msCH12bV+tVdxXqzvt6rosLqCkSFEbZngu0jnVw9rB6+hRzxU1i5DYGB
P9CYidmXIT4wUFu/t9CoBaMhu559QutFcw9tDU156UkY+l14FxD7LmvtD4DJl06AgJedzf+GMwTv
zEpxYMIYewiQ6hzE1uJSDairPY8+x8/4t/+29yxh/u9+itbzkDuemi08rhj9tY8GVML0CqF1oq4g
B5l6eKvcdV8xm4noWf2ZaIt6r2NppkkkXfJRWtIxxRa93WpKXagah+pRr61U19JHDHQAEdh1UzR9
UiERaDJHSa+jy6n5LMZnljVBD7G8U4EaN+OQmTjSnJBTO/50m3fvrLMdCDZf8u7rudPtwIOAxxxQ
xVznJI2YZl3ZUG1Fi78622b12OluprG7NMDmttJvqLyiaw+aMvs15RGAfnvm/M6qaE3GXZMW7qoj
fedaKPQJw+KQia3NUOhqLyfSJo44+dCBfGEybu2y+6xGoQbVSYlLYLhBti+UzkSA/j1ym1hFXb8A
yWlTwFn8q8KnvP6s9jeir0F+CUjnUwV66lFEUt2AK+PQwjzl95mo1DVcxF5DWPMCYVEigyBd5mto
QKOKa5WRZps2AA/YQ8t18vtImmWFicDngQQNZqJjn/vMvRhwkjU46rs/EN5h/qF6fPVk0oPnc6ZI
mD9bHXbz08QCUv2Ddnq7eQs/vEugQTL5J4MiHbjakiIU831y2QOh59ZVpY3H/qH4tTlthoB9cjhf
US8Z8A1Ylfp9dOURewLjhmoACKHpdz+MHSBhhf8rVJmo5hz/t4xmj0SFrIqFpBO5WWOpg1u8Wf2B
upWA0o8R3w2DcvBoIaJuqkHOgMbSdwrsSd+9SbyinlF+4+DnUvh5Bf9vDq+azPZQsyzVz1aRryGd
4/lwkkGk8amm8LQmuDLPmzJkIOP8nTYbMrA7hgKJUA17bIhFWhecZqFZtRwNLgpk6dejRCbS1/0R
4VFcTPMbAql1Hd7tJoelQS7s7CsLO705XbAf0+cXmsbGccbfBMCaZ2YuF/FFHm44rN7kjbSpyKc8
3TA9nsntZz3ludN9rYnwydbC1j1preUaOZ9K7xawQAj+RyQOgBPNOnagvQEAgmPCRxSbQIRtRUax
ynoPq8/8gNIyv8mS0er5/OyMv05/tChELw41q9cf5hzHDVK2Pd73giMAfqWOn0pRMluZ+ZRYolEO
dafnF+lyhm9FVdZlPzw1dI4DoCuWkiRXh/KhY2pgbc5z4CucBt6oU4Qi2gjHn8pbDzA/2IhzmSXE
93B3mTMhMkvM6JmjexbfuRxnxpnXkhk/axjvG1v36A2+CUPJ62IzGhNG1eA31P0AQpmBZAbcNibv
x/tHFmktZ6UEmxSwK9AJx4hbDDW88uA3ffc80+c9NuJMhmbM788bBqHbpfSN0fX7v4F+Rey5cL+4
/DYaiyL02jzs9Y/vbCbru6UvCyX50UYfxghURcFPrD1t7psb3useUjxNx2Hvhq1QHm8NV+L/UqLI
tqAwtd8Slt/RGb2OUKgqOcFp/A97i2q6ZFJCxiHYBLkmy9CVqNBYFpbPgVjWOp3KFTubUtKnlZ4g
CVg4naKIotXFIbFzMKPBYWJ3P0j4kt7pLAHxN+jDg+vgb6kMwz3qpJ+cs9MLYAxiXcTvZeVSWFV2
Uy/XrbSXMoKCoChFp3dGjojVVD5aXZN7zXFbvxnVvno4pxPpH0jeTYn+LiCYz+r8bhIaCF35PuHZ
pyBwZUDOW+sM7c5eBz1IVYCV+Bemghezyftm7ae7KvOI211fLKNVVa41Jv6h02ln3RsE+i53Faoq
RZrvLJajBT6d/7RQFI0LoYw3daQqU5VHof+JJi6coWd3wEmeVvIwzGF6cpJ694nra1i2MAfydWBO
B0NGTiejYooTSYW7yPWAZPYjLD9d8qxf5lyewBTw7VeqAuPNJsIbPhaxVIDwxn+VUtWu3KRh7Q2F
a8Sk430XjGdFS1KAzU+lUGaMYBcDYnQU0AzB2ZPU9tLZsnQvSMZ5cqcZB1xwOkwq7NL89vgNir5+
I9DiezNgnLDBbqRX9bD0ALUkt78uLgT/RGkgPmRCoqoSLiV4/cYSgjkVNg17AIZHtHNAUKqC8EL3
kNN00zdZWIrMvpxDRPLf/cyn9oUzTrQ1JdUF00fgSfCmDtnxr+vqKA7fF0ojZZq+uaL+r7nVD1eQ
jhd4Xw+n55t2Yk6Y8aJrJjrDrYePmID/toiLX0duf6lnQWkU96gn9HVUdXJJpFPfpL/IHumgJdlh
yHMt7fKWvMwyh4oXTkSFfVSMRdzvDL+09C2aw4WrCcYORBQjACtO+UhGk/vCYGqV+M9lyquBfk/F
rTgLhLGvtD4pJIgnCbXLEgxyH0jg1KPB6iQ9ygMbOQASe7rVMiiuGdfPKzV3WCnknCrPX9htx17q
acOyb+EHOm/d1IzkTMdr1KLCyTtJs8b1c+OTAx5uyMB0xS+3qifvx5LyfBzvlOZGGJiotIzfZE0w
gUN27yojhCx7kjPAw8huPp4YUTRhTZNkBmSJsZGJObixiGFRPvx8ZIQd5P8AImyCo5r3cScwL3DK
dwRHoO0MmPcdJXJdDYaTb8z53dUKWvCzYxEOcqLfzi/18l9L8cDoZih8eH93u5DDjqsVI3GzghnF
j0dxmfb9VEa3a9PD1RQPgsOV13RbHk+Cp2t8Sce0ybHz9EC3xfzBnMWux73s1DVzB9uqdbRIemgL
vCRux6zwGMjSrsWr4fgYASvXu+oj8flEQJbc5lCi6lDKAHc34VekpvNLdE4cOMAAUBbQRzs3e1PP
4F5yAyaOfFI1fsovkN2Ke9Uk0KU1j7nJeU+ii9fldutlrnfA8d52F74zr1dDcy5Cvszt4iMMOjk6
3l1ikKJc6q0mhvqrLsZhxQrSalWVavTQxfCXDstDFj7KoU1OQ28yZ/dvBJNF+DCYRCc5xfGqsV4l
6bRJry3xkqinoYHJN6wOtCJOfbXI816myAwcKhoe21kfuHCgBTCPqJedcnIpyoy4lPt73YIvB33A
V/PvaDaFybMpEgOOwr36HtSszWaTmhIHiYu40SwhbqYU/cxzskvZk3HkPSFQUw9o/MCvZ28P3yOy
e76JiQ7PuFHAAjBwR9Viquwd7vpx547eClKyReD/Lq/FwtIZD1Qjq4zDBWKSzbeUf85ull1R2nnF
ssanOeJv6I7OwE4hXM0HkvyuE9u/nYJUhoXn9ckeHQ4/UFr273MTomkPGkCn/8xGG2k9ShfbHuyr
b6j34fiKxcQ4kloDcpRhflUd1zKAEKr7olLuqOBZydIoosD2OlTxxlUNUyMcH5VwpBoX/BKdWVgh
Qkm2l/bkV1G0hUI+6HE85A1nXE/e5E8cmpWXjPCVR0qmuAKOsP7d+Y/zgNWugbuRoD1jjQzLzipG
lpkwyGwvjHZMbfUe9S0aw7zpq6RiNmCHQBIDWW3sIez99Vq7avaM7pDo2DxEFM/qHbnRlU8vis6Y
w4cLINatc2Z18ZZ/70svkzMZ2L+7c/ge5niV84gmL4h0NgFOwURf4XxtURalPmeXGudUE6u90ssP
stAd6KIMYo6cwIfaPIafza4009ugQhkDqAfQNtqCXJH6X1h/0yR+8tuvYHHQ1h9ymIYh9ip7t0T9
eq0TrkU5nNPBdPVLgWJOw4736YIvhAnLGQskEtA5lYiEA5XjMos2A4j0xo3QTmyWYe9Kg/MKMHf2
Funx7YWgN9Sk4KvQjBJE+H5UcYr3ZqjP+FSLI/FvnSfLq3SZkumSxVqHvVz+RJfKFn7rh+uxR5Sd
AA99Z85BObu8MT7w5mY5lvmds2Fd8PZuD/BoWteXYd6EmhF+mo2t+aLaO9BwVS4QfzCin6zX5U64
GXvsbd+37IP4ArzlIbJNVhW1ML05HEUzOEeQP6UGwzfAXFfFCLtrrzm/ggCzmw3qinNv3j/ElEJL
94mp0oY5AAN2u2SHLANbLFt2Q6eaB+3cayk2W2RMCimNSFM2iEtHMk27dPsSbux4KHABbrZ+f/sM
f/Y6h1gq2063AQc5mc7zlDbAaPdZd/RBogv/Ok3IvnzesGz/kIiL5rs0FtLklYftVOUTtk9Ae5BJ
npivRzsHBVuVrPjWoQj55bx9pP5x0ON/xIulr+RL/S0LfBxQPiNz1UTn7svbHM2eozb9v2tIZBwc
EVmm3JmLVqD/u2gc+vxr6NV13tgOfvQA70mQLDXpl4LVG0JnCoN1q16hgIaFe5sl57gj8UhgxIHe
XB8fs3QjUjYms066VL9g2Uc5rm1Cdo0eaH53s7pw1kvqCgrtmqjM1CgBBu3CXwx4pjftG+ezfeMD
nRaOR9Jq7X5ksMkHMDYhSWa5w/7Qh7+Rhs4v8NT3U3iB0esqYxzmLprlZLBuDi8x+eIPoLImuNM2
qF680s+vtZAgGYAPi5wWKPIh99cRZ8Tv2boWmu9D3j0O2hrlL7fODKjvh4q+E+pAwuCR5NqUkFnT
IZhnJBKyTfZoRXLuSRrhUzRM6fgqJvhldXnu5uA4aIVilZmGCd5AUSsQIQ5H+/ascnLXN5sgN/Qn
BjCzgYdzesvR6KKlLF17Cv23aa4MjYF3f9ZlK4uLGe/GaUCn8I8J1pdhyKvKs94QOjFD+dtlW8cD
aXFsxWs3aq6gtR1M/uGfkiz/8G1ekKyvfSAFXzZZeW3+HOQM/sTKbzs66DReBxMOqyN4ix4U5/qf
brRTpjcFqOYeS1Q8TDyp0r4l7Fl3qlIgVJcXPYZe+WVvhPvlxcrw7Yw4apNEhGy497ZT27w6nWdq
DvlgeJ9BianVRx2Ji+HGhEpVq7VBeRzj7fePkXTx5m+4ObSiOXqNXjsHjOX2KpFDJtoSusL8tEaN
WVLy+XFIQcjsnoQ5+uVaTCl//SCWOE5AVA4Mc/2VT+2/CkI057CHeleNc5pvu8J050KKLZeaTw/1
vcVd3D1Qi0BfGfT8oHqCOA7GFvvX6IS4FMqKBDkmfchdOXs92j3+T+2lJ95M/KcVKROIGUYrYjz3
6ZDWagu8d5PQQPIPAa2YIDKjTb9+iIJcefxegzoB5OVLJW8MabPl/TXP2sIFUgXvkY6bgAWoYPmR
fS25ljOoqI4i4YjDC6DDo8LFnJJtiqng5ZZV4ZdTs+JbyE2PCvUXxUPUNlJrEsIoQGzDIdyvXm8g
Yfd1ooXm5oe4psa06AHR4Q16ibhdaxERvxPNkgxhkErLAdI/PuRcSObK5ka/IBTjeOxktmHaFVpM
PGxOvzx9du3Bx7yPfQ3BZJsYtLTjQ+QbhSDnLFYUK2QS9UWeu1jF986HZKQVg5GMfpwajKeAQ7Pc
4WArCuFOapcssDikTTbB3xZ4Wei5z7bDZlxRtj5YLkPNKcYoKsqjuKNSqRp5AQV+T10u0k4IsM8P
lFB8XXvHjv71yDNa/bNS4kKZ+aoRh97HdPil5zxShviaHajPGzRxrFEuf8TpYdK3+NsBMMo3BBKn
ETut93DpCCHX50/GXmuk+YAV7Gkr2nv5zGrKszQ7JegF0yJ13EIDX6Pdo3JIg7isMPdt4IHsRjuB
QTFUcl6khLWEf8Bh2fiXklBe+FzE3bMaa7St34Rd4wWEx9Ej8+7W2O/bGUgTfUQ6RTyVotyWsKcN
VAtmFHnc9OQ2VU4obPxII90ud+DWk0KVI/ioXsYyrPT5B0ZWA5bWqe+tGwDxutJjsycDzdoRUORl
vuI+PXwfNvMtAWDoLU19/f2j1icoEphDWoUYpLHhtnQbPzFzd/KU1CoGpYydt+WGfZLuPxR+yyCq
DOk5YdmIf1S1C+/Xk/W1PvGqxkrSJ5cUYhJ+Gr4sVoUHxvzIyOlo/OtlpzNZ3fCobcnsM7vsCzNA
kxsFYWmO67Pea1K3ICdENiGZQk2mLXOuwNSZCV2WKK9cnLbousey87y39TqNbxGrI0mYBnuF7Kut
7n9j1qdpgxHTDKY7nVhcfwEkWAzIruSjqkgrX5+1yET8BoFTi9IJp1QSbllixQRsNeQapig5Z2SK
fIUkuJz4qTUZOoCdb1V1j6CyYEcJzkWTPAb7pajn48Z+1vDusETNCleJRslZAzbNfQUd2PPnPx/D
xkQjOZQAF1lMhdmn/bDZA/u4etR5XBzu1CVAAT3ZMNMlb63XkPXsbeUnyV1tKgXAy8aRZdqIDcda
w+dhnL3RLfdZdB6LDaJYNjMqjl2Kcyi7fS0UmBH5diL8Tqfyl3lbWdegxR/8rihxzntFK//IP7KE
ByV/gWlqsqDbPUjzjEc1/R4P6D/AQII9aKdrbZAw5F9OkVlf0JMCwSaX+KBO/t+RIAs+VHXUREKm
YdP+W5DBKl8bME1aFEyu3X2AuOGCPJeAvWcPdlmv+RuXEz/ItnkebHOsusFEw7Y1FPt1H25QRFIy
c1vi/C9NWdq/IzCRuz25qtWnHyAmb0Aq83kwqLn3OLCx6NmkemEKBw2rfxuegbmaXP9O8OpWNb2s
0IEgURzZJsQU6YV5M1gu9jcV1ixQ36ijOOfp8MceqkegeFGhWzIEFv2EVQ462k4VVqqE4Tgah9sO
pVxVHVHtZ5W6Sg2qywGnJeap/8xSZCd6TFxNuK/OgBxbmTggBInkVB/k4MVj+mlGUwJrqBueDYB2
zDLBIqu+rIgqYq3G+fqsqpi2p5RAjnLGm54Nux/NTyK7jB1blGy7ca3Q/fZ7C5ogD+IAUwex08ys
VRWhtk4ENTH48WpYe95kZAn9XacymQCOcWfAZMiI56kjyITvEdjmHpSLiidcbIntp2ifrKK0j/iM
ycKCcYm//sp5woWMNzSBmCQVZSNFEcmQuZ6ABWW7bSHArJPMMcxyxGQq5+SJvIXFC745HpAGeb+T
LeaXenfOv8n2uYYn1SSALZmWuWZg6cWrUdYG6RHu8mpZEXhD0dRSeo2xk1pG7F4LPl12kgeXpINw
ObDLZKEv2v7IXrjywrVEjOfQSisufM5+ROfJThXMVqZO01VIwCyv9ZxTRVa++ymGc98cd8r9dS4V
+DnMGtnd72oTkq9ifvNKpviSOabGTt/m7J/8VKVBNh3TzXNwwTGYR6+9lc2jA24eUP0Rat1OtRQd
HJ3REw4eIwkY5tZrL9h4/nk7YqkZtPVOtE9cLdHXuNl1GzB/makQdRL7Hz3Yi+h7k5w99re0tsrA
Xjfq+R8fhckzkrKhxzhR3x5/CfJjU541sLcaqwyNNSoUfbqStQUPzR+RRC54NcNbroxApagm/OyO
i3a3VJ8RhAcT9QAtPuWabOpg6OY8C53PA+WNOZbBFefyz4Dc2tGWePmlP37GF86XK04yj7ewjVAp
aSVNkUSpwkf7jSUY4MStNediPJ6liysEFyj+6ooWIcTXPV6wj42wogth05o9togcUaGtrqIdX0Bs
4Z+LPBedFhrImnGy8k3PCakbuRp+D+fuc19j4Au+XQRB6GlD+mEEMOnELFjSBHPOOf71APoaGEUG
7dAbw1NSfPnGAXFKdIBarunXgfhoAkG1JpaPxCDy2QkEyM4gDm6xr7Gzt5kS4uTtgU76VWoUorjC
1FMqz8HGsUg5Ha0tnBiffgtX5ZK96GplQhHLZV32KF3Lu9OPsN4/gL0WWh2sINadaSelHJ4ad+sb
3V7uupMuWS1wLNEXSClWp6mhFZtayP7DwWMjOzz//3vBd1/nWuQAZPfXQfquM5HAxug4mN7VrYuM
JuamMcPNmltOtGmnFlT5IkO6lUH+bBfL6pSmCC7eFQOqGNoonQ+shEM/zWu9WBPUHWAIM57+fRmn
B3T3eG7P9TKwirS50FIptcsoSIL1QG/A12J7eivinULK1JuAjns795OU7w3POSpz48TxFne7zxaZ
52Iro5X8FV0GDGrouPgFi+aEaIjtvYvTag4ZpEZ0BZgPp8Z5BX8Z3TqblupmvIeqg/Y7noMqUon9
VaXTLQrWaW1k/zVK1Q58zI8+ZsIUZhZwgRmzx5buk6SQ9perhJ7LnDtFym1YoDZjPRozz12TG9rY
fcKrqzjG078jCwtnumqsZOE+nJOQaHJ35Kb0tN40jHoI6kT3vxy7BLbRnJnSmujrGbzLYmeNZlDH
CI0LpeBJNA+pBJCVClCRf6+LUk0xhfYSLmEZ33ZctOE7ESgUZKN30p6XX2vgd5YoPqHcjMUJPEyq
Ow8y2+VybKbqyBfP9v8Ah9CX0OPFUH/+FGt0syDvFQEhRxYW1Cg5jh45HsHQMTKnatdw5PFXEQQp
psw0Vs85KYw5qLzmmzX6W1q9fDKWozrhqb4xOiRsa75VKQaLB0mssZq7wvaJUeWZBYedo1WFYRK8
UbdI+bICLdTWEH5mHEqcf0uV1r3RcZqfwj6aM7t64X8PX5KMzdCUbiA2BVzZbpfobT7G2R/wzLbE
tUerDsBKRD6n2MuHyIzd5ERlC6qjukXZEE8eeQp7SKOpZVg5dTUmYpfskzOiLpFWLDsxw4FpX6T0
/ZIbOUmSsXNCgLuA78Dt997FgNJG0bmHCFUD21B3aGqOFTV4IeaGes5RHKzy54gg21A3GiUNgdKS
2N+Lwz+DoSiaRggMjL0OsqRjuZLV/EmSETUR97LK0lH452Makj8IulGTxgIfLLYWy/xPTuuqaBFT
3/Thq2+aQuXyHsQFAVtHGP8WcuaBuJ0z2UaI6nfOzhK5fX1+emlTv15fvW+6rJNYUGoDRFYZiBw6
k234Cyp0HuBjctPg9kV1Lhr59p5mBhKQx8FO/SOEK7qwk2clRpNs/JIcJZIkOgRrb5/EMDpxAZ1K
sCPGZ1UGtA+YSkGfdwDhHqEN+FsGvlUVah/2PP/X7ZbOxf0Q7boLGFx5GnI1kLzc54wrqcfXYW7I
p+o6pWpdla9iKOmj52ASidBxfrEqoHrdhoc7L65Ul72vmPM3uCoTkNMY/ENPUzJDsgAScW4Q1FP5
NiuRIvNsq5XJwEMWak7APJwymo05iurVZRLe7C7DCKh1CBTNcyiF2eGfmbo8iMb1ILm2R+tkCp8R
s5iiuTn/2xTD9L4FOxzwSTbRFsn7wP9e2RQA1O6QFO9lYUAe36ljXctPx+DuBiTBxrkhz3PqRbNf
40aDNYF4XHBRjmryXx96C08my6/YrPJEW0el/Jq5ssH/zkjdsIy7lrGIlB3suuHx2WouIqRUfC0X
10cKVa7oofkdFTheXR8GVTQG1A8RJyc/gLfJEZka5GIBKIff8Tw1kejCU/Esh7N3ShcEYUvN12Ng
SZTwo6quyQMcZMvG+zn43YFnj003thyk+3kK6jIQHOEF5elZ7s6fUJNaqrs8tjc1PXitbplTLQUN
I9D/abmMQnzil+O8RzFaVpKpWYzNrEJRfl77XRhuTAwY1eV5d19FYbdkB0Zx34etVyITn+lmi3Im
iS/t4cMm+rVIf3kFTu9pSpET3MksQd6qJG8VhWmKdpaXWkDOobDNeRDLYl3JVr+C316oq8JxuKoV
FwJqu7dcBxMa8GDtgVQ8tTRSRnrgTYSSKDdifxq9Vy08f8dLHTNpah46RqVsaAkUJZGJOR3tk7uY
HWKRV0flRJE7ASN5BS85VfBiLr6AEf93hMV+VQSzhgzrvwZa1k7gGG4b3iJ/Bu5LMzkyLmBjmynT
+EFSrFE0pW2zSIIv/sfiM74+jyXunb6zHwp787gAiUJolVSOhUIim1ab/Nsbn4xuCDhJjT+V7SZ5
gDoFWVVPCtjOGmGP9NKZpF9lJrRj2GIpEKWUGzKBwpFsWac0twzWLM3iNZdULnSfF+xkU7eePbqC
+Nb7QlVUGgIV2/UE1G/PbMXdp8pa8I1XfwD1ncLt9RKojwd+hNPXD39oJMoEOHwLQ6lDs9/8Jz6d
mR91PWAQ9JcGnc5p92Wj+4+q0OJntyCGW320wuE75B3iFGPzl+t3fFPDyQhvA+LcuQ9JnIqntWX6
p5nronZ+ZrURVnneMzBLIKZn1DNnacp48qJ1qj+g1KBRTdOFrgDdDYsT4o5gKqwjn9SCQQgljCvX
gXiU7Gua07vWTxSWf6YJo0hmxVQbt18kBkr3qLWCksmShqRTeP3H+Tp9ofjNHpReBFe7ftruIAgR
dEHVx3PYShh4wqvLRphZb2D+WcmIHFDKzb7+XPWuXOlD1sO4Lm7N+7qM1qmdNgDVm7m6Gy7oX1J4
DcEQdB2QB+Kjp2OWQ4SCYZL0o6tBj5dKTzV90cIM6fcQc4rZ9l2ozpopNakVTgCpINDXE7DKWO/M
0DtLtLXpiA6rkpaTeAghVbijeOPNPtqqWU9ahZgcx3U0Lkz2pEAmRA4Cag0t7ejG3jK91jBTNsYh
dW6LvCFBGJTRoyQwoKWXMOi3vH6Sdp/G8X4Q5HvhZWk02M2Q71M3KRIOrzD8sCbJAHXt3auasQ2E
HuWLlA1/abcF9asta5Iwqb4aJS//jP6AgGXii8q/MY0wNupB1dst0CSlVaw/MQBOxHkeaE/VMeJ3
WHxC8jqqVT1btzoZaIaqG60C7MjhbF/DB0L2k0e0xnXpL1mg8bcLVQzNUalKiaQ9b4j0zfiimaXF
M7/KdzqosJlbhAsLcO1OA6hcePDA+vwbJkRtbDrhgEU5mch97Wp1de4p17Aq/gjHF0TXMtYwmh9G
6Wx0mzrhSmdCyrFGvgIgaLR/7RBDJF5mZKREyoCN7zQwragiOSsMojTqFc41XlZj/FFPW4RC+jzD
qRMlr76GUWuZklPKfaTuccOJD0dU6Q4IDDHyMMirea5rA4F59RCRBa87RKPiip6847/+uKpol16V
m859e6wfDeu/S72+IejEcNrQ/TYvZufF3DgKoRQBbHzIMDTnPVe3AWKs4nWJ6n3FbRy/zPJi5vMY
49LPsm1U0UdXcJDWGr+YHDg/b0gn24F94TIMqWFdgBsMIZsVd0YWIKMRcnMHLUrfXpqa41g/5Eli
ebdZCWC+EnVYfZpd2YvIyr5WMgadIGsmQuB+yzZQ0KUpgynPC38mezzIvNcRqjPVomlO+HITeoSl
1mBPHeESdR6FpzgT6W79LG/QkOghg472qOPXCVFiXcEofrX2T01VAKE25rhJm6XNAec4k4TVr6BA
xQ+hM8BARR9q6yBRYh4kcCYcWtrkcIcewZG7eKaA5NsAj2shQhMUQpEisUtfQiPt8IgsUJEMz5lv
Qj2eNbdSVWOTtxM94RkHHpaZ6CmEwk4crMyw8xOQbHVMhonQBSGG7t+P0ivlCKd/sZkrfR2U7sZO
+ZybHmunI/XFgYbNsBh0VBKBhhTcfNJBDsdiq08e9/Mra1ZvieMqOYFpf1H43ODEhUqfJgUaOlJ0
NgLWSzp0zIJS+AgGtqvc3GFDOEDxvV6IVHYwAByZINUndYkT7pdO0QEuGkmHu+3oQXhhBN17Vvlt
shfO5rap3miSKzwVnjjwdiH/ed8PCiDFqTS0vUg/7znxvD8vYz9Okx9MKxdZgQoYaos0AxnaJRGW
QASpdhXgxUsyfzGQUdAy+ZG49CxM8lwUHvNao7e3e65XLJWRvGsFvkEXH5PD2rG37qxKPs2f5jJO
cYU2uNLNtgZXSR2BpLm1p60agLQsmp4jLmS4EsQXv5/1H3axb3h24Dlun0zUg7I0Z4Pwp9JT+34n
udYIuLYb0Ib6JnFkY8k6MhBLpOXdhg9m97FkfFdAFPMtSLj41V7kMiWVFqdxD+2Spyy94WfeWI4i
yjHuOEOoIK/qSEQ64XnskaTzt5pE1eQUBsKrEDPQPSDyDLY5DeYvYHuXm/ZKIcnFwNjTtfhhlOrX
W7nYXkBfwC27E8W/Ai9KndPegfFSZBMEpDXxdNZpgZmhqjopO+Gw6CnOS7yJxCQZRhMWvPtPyNKX
tlwL/+CmsoZi8Ens+4kv8T2jNFxQJiqLgDGqJkasK/Dw1HC9cuvmoiepK6rlzuQNSWix+qNwZ8sj
k1UzmZINBLLxd7yROz1E8ICMpE2Ln7dVIgZh8mq9zO2IcZJ1/qL3pEeFhrGqdmmMGsH7LgKYLE2W
ZZl7n5rQ4Oxl3J1LCHIwgFvU0fXZBWvm7WSPvlKpl0/HJ0io1ds3Z8hkfHQjFIEM9VkBBs4n/R1q
Wc2uhjBKum7KoaPD/VgSSoInVdfFgIeZ/vQPIE0w2TWGwWokG9RRxlj/Cxf9GtyBgfyZWFEil/0Q
kpVvrVTpvOsJdluVndOwNU34HpPeGVniUpdw5Slda6nRvypJB8dD3+RgUdWqxZtqDSfOM/gC5nuO
gzkTN/nNGlo84z3MdsmAOpfxLi4H2sf0Uf+W6zeyzX/qAlSNo6IJ+EyJELLroke8RPfFEjyRiOVH
ujr1l6o48L/u18aCMiOBB9Sjhfte+1wk2HzKrBlbsY+o5EnSrAelNi3rMy4atbleUu0vf7iR+tnN
1NIo1D7rZ4OF+dRg1EMPqE/NHRJ07cdz7gZpB43mZUvWZowXRBsgVRWzlSHyVsN4+beZTAoWpg7m
V2v/lOWVZ/k2F3r3rI+Zqwg8ktEUDkfu2UoyuDMs28rmNHCt9kuL+iAM1el3FHhQjExDJIffS081
mKXvJd3YOyg+8luzq+73C2zb2WEIbrMbaMqqvIukK1k3bPTpoXLoRGet8zYfPzXVfIAhUsLeRKFw
oqjM8DPj4HCaq9Uw6vR+/sr39tbZP4/KaAFyV/oj0z54+GzSbTNcdG2/yo61BnxcDsUQUuDRjZLs
Ei6ZvhHlwjOlxzDDHe3/V5q6N8zX92bd5EVo9KjX89b3BRZ0Zm6/v3Yqov5qeXuW1AqhdTIt0UNm
1kl+Ug6ylm4O8JwdA0Sdr/HU706wXG1EumujBtxPjvApcZRIgE82G98GuCuim8fnDmQ4tK5ybpxt
kWycibHIjLv/Gm/ig1jBic89JAvncdngpuaRvPAJqaPa3UoGvUQaNkh+U1IRcepy+pn4ykHJA8ME
XDjbRs+AtkxawaxamelNYrefLHAJl3QtBf5pyfSWqIYmLFjmZFw0RXHF2EsqcIWTOpxGtM6zOI8E
pODB1Yzu+yGi87WgBekdgXOMS2WdhMrebzON3xjxHjNq3ej5FNVQ+x6+xxMhBO36ilLP665NUspD
tZ6iS19hrUt9oL/GM9A3KbDncZoOv4LH2AR+vAnsIanm2Qp/TRq/tIeFN4AJze4wYpja4QAkEVvk
LY9pj6LGO7wfJ9Qoeudzzf7BWHeH/CawgC2qIR9NkL68yHl5TP0H8GN8FrsfcC2LRhvaVjI2zsPZ
I7CKQQJNZe6aNM5D7I+4yZQRqwibMY7mGZuhytK7dY9Gfw3mySLSWe92EVUNMOMUBy++Ni6pETJ6
HfSRi2oOPSpekCgkk4fNsYnNA4ubFJSh1LO4GEV8ttpVio4+oYa+faI27CaTq5uge2Eb8N6wUAql
0sJXlqooShS8PTXdEhiffwQSDDB7JHm8d0WJS1dWhG3Bwy7C41Ls+gkIcnexldrugmx8lQiNSsLk
ZfNAAbwiaQ7Un9i/ck0NUBL5XRiGNtKqsfpK3bQL9Fkr1/ChyksARwuyEc+v2PS1OzlwwTmsKYv2
500oiXYZOHnoiYz3zH6wurImcREErhmbR6yGmLN47xcA2GOnlVI6a+IRDmu59UyxgrlYWb0mfm8I
Bu7zBDCP13lavJ+5ZalHlAmo/leZ3qQ/hWR0g4m4BMPNH1ncIIIlix/GdEh5Fl0ZEraP4LSNloW2
I08INjraEsyKPNf0islJM8MRmr2VWPUsj1Nk4xyQyFuIcjzVbLxH5nvxltRR08RIH/Rvd/U8E+EF
1NInDxICwq8XmYXxdTas/8W6E3YqZmNQErP9bNH+nKMOrEAd+r2HH5qZJOELur7uNgc+ZWhWKBKR
7OlPuY0oND+rOCaYbbQ34riNOBmGyyxroG1xTpI/85vWPBnS+uOmxcTKrQ995v18gQ+tifvdnR8X
TwLSv0+xFNAtd8KZB7QkpXpZyPGae03Lr47ai4lLjdt9Icvj/ILV8rv2gwOtdPhnhYJZumLUfx39
F/jkyuswuxLKXv1XYnFOm+z6vdyZJJZnpzRXyfgSCLkpU8KiTw2l/Zry03qKCqWQ8tYu3tHnvu7R
TcDNLuHxCbTlnbXdDSh2i5mHnD4TVaX23t+/nAf7WzNCMdDF6odzP23kb0OMcinXFe5A/s60yww6
8jtXWbcdHATjySigR8M0EqUDYqM+roTj3oJ80xilamFPPEhl1rC2FuUJa74k3o21zcIkR4tBIwjg
guD5ibr+1rKoHQLjxPCblqljmVhQPFwdFMhayX7Vo+8LRPhRQuPryb3Ei2xC4agwkJRbrk79CS1Y
nPElK7DBYatDTEJ/DfD8U1Z5UC31FvDxMiqQSuTRWdK4rlj4sAuZB7tW04j4LBNa0zoUC3a9Lp5Q
8HJv4uEn9WwhcLNZAZuCExwLO0iyhRf/V4/6fZGpaZKqHZan4Jx1MC7GvIYJ42bB0wN98QhmciXB
HXHROi+Iyq8S3iJo0ldRbF+Hm3uKkprYDpBzddDXqhJZdr00XANsNMaIpJu4oZdks/3M0WWeVfkx
RYu5XVadshYr1CGceBP8ITAMjshltQwvsHicOAlqepdjtNnjSyl9/UzVBXIGP/pIfYxCiJLJuP/b
fs3KYZRsiLZLz9lO3uwevpbLakNDCQWAz98rpo7OM7Ook2wxE6WllFSMuEGGK4zx0zTy+/3RzvQE
ZZJOGWO1yQoLzVXW6YI/hbaKeAU7zjV1mW4DIBafnvAdhlHSAt5t9OiXb27f+K3jn/sujvU7iY7S
TLj85Hb6nVBc4KTzdtQ19SsG2eZ9wOuM2jmG8OSbmtgm574vo2mraES7Gqm7HVStRNanwjgp1kdY
icXHuSoiCFzU2MXm2sLp2HNA/V/iVooliMiNJ4bnywDjRhgwRCVrArkVVSXqO/sJCD3VNKtFLKJP
ZPnjOVCvylnnnjEqffDP08Yu+mABKe9awwnlrxtVaFSA5gserBFcDDjw9JOmI10IA+XCjJ83g3vR
QlJiP2SInzin9JHYGX1ALirTUB8nuxe1Adj5qgvMx4L7gvAsFJxTQGkA5ontkIh8CYXoFcVOiCeJ
TfXHmWBGsBDiHBp777Y4AlUmDRojir1oOI004c1FxlIoS2lumiwuh64TJxfk7j9Is4HM2TpS7U8r
DYwhIVPZumF0MZU54QRgs1fMQTxXubID7qM5Ah+Mmi8OIaHrZzrcuf+7DbJZKQOaCEpGvx5hLKX6
iXEmh/o4fnFhI7fmjSF5NnX6cSaBPDTiD6hJRPAL05Q5JuUyTp/NdDgNpTAYcEepaZtOWIdvpN2D
YygwhvTug8ywgMTXGEhyY6MhayVYqq7v6w2Es4ZwL92gCJndYc9X0DoI4mcpp+rIrX8Hf/zc2gYw
049zkCuc144IAQ7ShlyjiqT4SWeAAWdpyGZiSLz8h2xHJlECtcolSSM9SRTFzd0prvonK98jJ1J6
DEGravEhfjjRhcGvUTxkZZjUtyqEvUSPjKShwM5PCIahm611Z42HOv1Csc0K2awiEZO8AizmUCjT
t9FPdMnaT7WBapDDQZIm8+8pOxmD2TIE5gDmIePssv7p3ltpPiAUe0SW/em3LYSYZdRgD0LGkHnL
9tEIOHFLIEFOFdTgcOOyChJ6WRKITFfvJTghcYsz0cB6HgMUIdDFQHGfLFAaPabYPcsmMa/5J1zK
7w3762Gybo4gttzNRcFtAYNlSjCLo3K3c58FJVZO1OaxRMx2i9DccsCIARoZ64I/ZJmxmoN+ciDE
sxnNL1rxh2reCDEh+fN8zhbZki3RE7wDGO0mkP4bMaO/jn4sHcffQFbI2OmZXuf6PhG7gIfR3M4v
vqZ5pzRhtodaFvVHnw76/l0fB6wTOeFlH2x2dtw1Ksagep1LQ59OUpVTarhA1GSAFwY1j1nFV6Lo
6SRUPNY9ueTZtXgoLX6lGla3j66MjxZnbuF7TT1RiVqwuhRg3Z7ekPm6CLvpJl2jOaTZIQm+WYCL
yrA6ZzCQCVv9ZuB5c0SUBFLKf/pwStQaEteBuTeEmPblygPDR1muBH+noxwVA2bTZRmnhmRRAaCi
ZCgyE3kQLCuXq7kfV7nQYCRUuBUd64xV4txefpXQ/TEr5nzSogdSMAA3wBmJd4ztQqbtde0cvFER
Jl/lCudXZSr2uu/mxe9NHCqqRJXzCZ+IEb8YQY9MIhiuG+HNCN4otRLr3G7XIfl5EkaJjw+noFUg
DmJqRH71fU3IVsfOAWSRqwPB4xSh7VS5xZLrJDEBDkKYie/G97V93hDr+qcimCJAn5lYjgDWW+yx
bExVaJ+QNBW9QnVGGPjTFZ+/0IQCyHmfI4tScd8XWI2ioXXVJcLkyJ/wq+1Vy5Tx07AIkGxY/Hqs
lNOE/snhl/OfeEGLN+YpRh9EAnjpCB+blSpJk8d20BeMUGZV7DCHPsAtsZN58d8r6VgvNVpXt/S3
XL1PeVpuRMAbV4fZInWmujqvAjh9PAIgXZMsaNRWvi2yTU91AVEShEwTNthAFolXM6SEcwuz8QCI
aDsCmgrSRCWEaqKJyDC6UpGwhNbOblc+5mx195EEeKF3NjJxV+E9mJUkW+xx+idyg+9YldEdGCx6
KfGVYsTGAcTimntWBJN1p4zaWvCj44/XEKLEcrW0jdHuCnaoSBlIMYP2Wr7cMyEhfYAJlM0uF9kY
1AgXdkalnqjg6NCgR3Q1cByjuWHFZRNhF//nGG7rPHQPGSrY9gQ3LqzavpaFTSXDVGa+xd/aqYiE
zRy66lQUMCYfAkjFUCx3ETkDg0F/KR6PdsKzWR7tGKblplw3hSP0Fnycaj1FDYD3vjiJjMCyWlID
QW726YqAh8Q4CqTqFQ8/9EiIv/w7+7PpLYSkqZXBYITN8dHeL/Gks0b2C39DoHtizZ8psoJY8sWK
vUyhCky/ElmxfT9DMei6MSD6+0QN+q+VjS9ExGwT7gFjqoFRhhRqmEzvRHn6Kz0fAyNOVvO4flkF
IiqOmcj0MOkQNBX434BxvYvnQCwnDjfSsCM/8cbXI04rYRMu86WG2Bzkk8hEBiYhgiDcgULr9bhc
ssHIcmZqSypWRJh4r8RUeuA9cw2VpisVmINxTKfCQ+nSI2bUtjaAfyoRswp7UTFNmO+zGPJKMKpt
6vxDceSIX+DMS5gErlEttjN9AyIgZuonaApYdeXvSAhYid0UwXllcw+TFO2i/RlzTk/aQE06i5ad
Pem8qKDIuymlFzlH2jH7h4DxjGqcKEHPo0SZJTIMp1x8SjJbQ5YPg4RcqXv2mSsN9qjFuAYWvmL+
JwfwxM9qjNwq85cX/KB0gWxmVcVAlQXBTS2zAfqFWOxOVmUrXrPhf5UiR4mORG1J9gNksKV7FBr6
ybaQuQfwa3jWK7KH8N7A1RhXGgG3mj7MUsa7AWzyDYsN0bNERujUpKFUKRJmd6MwAyx9nDeuEsny
0d943bdj2qVm4Kv/Xeh5vH5DmEhB60kUEoRVAgiuQ1E+G+6LpqsgwY2Cqq6zWoYTfx7boQZtonlZ
gdgVY6R9+hAncsir9uyYTIv5ZVtIjb+jPhvhRkqq/kbuZPz8iGTmdMYOSXwroIpaO5w58vpwPnls
Cwid8jnCYIGGZhNO1lWMYJRlAMpXIg99L4xnfkHorI9cynDOrYoOt3obhHGD2wv8Rdt8fVJg3AO5
p4a7+gcZYFsgK5I/+K3PNBvye0mDtsHUFcqYj/4bQDwGPOYHla2+iRQ+i67uLOf/+Cm0nnqUe4tV
brljTIUSTtv8Zxy38ZaqiAOJ6Q1SD3HMBk1cBJ4TnJERAFRiIZfuKYhtIIFzJhYqLKCVSxwucY3n
Y1QQ9JQnBzdQLFnt/o0NjiRoLjlbTsSNB7g8ReayO68+pAi+Kw1fyd/pLEHGyM9V5ig61dvAScUx
XShIISsoab8QIxo1R6GsBhHirBjrW/sqWMOUCpJcy3YWXzVvR9TPrt3xu92Zxizjj2Bfj6DAIr/e
y/a4oSRw8OXVdctl3aJ5pH/xRNjNpiznzaGn2i5eF9oij1UQMyr02+upiC756U+RQiht8jkVhqxM
f28XRn8zkxBxVAxfqTH5lK1YNsk4JcL4wwKfPeKEVlsckq064nPbtI4VclnibGP6yxAbT5X1VA7F
tAF0ViC78zSZkTCxw7hKVw1rok/Yo2Ai6rRm2b462aY9sfS4GmKK2lU/dLJiL9YMURi4XtLopMl+
eJL5KKWVoB1UX1KDZc6Jq47WZD5YBWTwdHOhnBni/59WJ98wS4HMWmv7AZ/36aaeUuo8dEHLsatD
/+SBNefEzeVxlNfR0lAIVq3C9vNyNv8fw8Bvkc3tonDFrrvxKCF3QJRsy3SXhBFy5D4Fcttd9Rj6
GJT0dSLbtT6zF7U71a8Yk4n4+pzAtiY+nG1P8zDqko7E4Gh3RHmEpdo/fsINsR0Xh/+4ErGVFaeL
QLfRZNAn0rV1pXCwh4E4gwyL4/8aIgWVQ2ZnKjDjHl7SjY+jnORrYV7tnX+R4p2jkA1ryVgI+a63
Rwf8TEZcSwJH5kIUI2dxY+rBL1JHIMP8OXnH/O61flJgTlAndE9aMDOYFSaXxuShWZDhHwBJXxgH
XC2HKSCHnenUheNsAWaMJvWTiUjkgXi6UOqMq3ZtGP7C6PfXlonAdFLPWpacY6wjSBr5U/OiN+nB
iPhj6iA6e1qD+83oHodVnTlN/G+KrkI9BxLjgDMZjeFxIh0fd4JFM0QH7mtOEuKWS4UT7wjYwy9S
LKosBaTllqOvjVMHY/vObQHJBUn0JuQlQsaikpmLnFdvIB+snt1hMFs3DQIBRcn4++eJ4mevI+mw
HZfxCHz3h17b7S9ZwjJlXwpfKBL2/uk83DEsE0dVVNsoXnfzviJCXQQWmOzpEVx42wcBpa3YJOFV
0Me2YXyNW9kWJBxX1pz3MwlCX9vNTGjTtWayTbYsXTjDRSZD+Se7nMEHEMxRMfGkYp/ibI7UjCNY
BCjEAiQLbSnfqhc6KinzATP/J4yN9fK7YW/6qoGG4wLOd372uREoltkMVaCZ7IzGltcPyOyYmnZR
2wGWFzc85zSf1Y/Q42KLLTflTjBVlVbGIUqVIJ2LeFP3wgMTmwr86G0IL2V7vEbrni3v+3/JyGIa
7hAkDTibR6hEtwpssfmtWKuLuWBk89M0VXvSU0W96a9elEegzVY8lgIPHg9AbXw8/yn5+TK3U00G
ue4RPTztPkVyxnzAFLn1QMHF7MoHYWKB4DBw1Z9UOuYLRzsMYaAITn/8sHD8avQgontfc9/ZwS7X
6U/9ve0Ti73MI1op9GJ+oF8ssVQAsE+5I3QBCkkFcSGItqNZJFXKP5V/WnfDHzV7KmCFY1I17fZU
ZTV9XRitOlmE9/vkOXhisRHbz04FU1KDtBnRX8VlOUIH7OIifOSrv/F1fxNMJSM/UZL9n97PDyLW
TqnKIgPsW6vGvKi3buyCT0zQxgq9hqr39SPnipZCje208nW/AqZ5xQQHeTwPVMp1mNjq3eQZPiFQ
2lBt7E0psZs9mc3dSSGYNG54YOC1Bc07bl7GOABk+aYmwQpxfX7hCsvKgvAOozAxCSVrJtRf6kCg
7n14D+1rXisUyvRCcN1ZDiixbR1sCgwwdsbfDQVwY9failEJHlgeDOTJwyBQ3P37qIn1UE/lQh6q
bZUel4ngge1mYe5iEjWWQLcD/dd79LMikOxUEzyJ7wSifvYm75BjQipthhZc97O6FCX0cQB9JpDO
St1ELdWoJcpm/ipMiyf5KrHRTeg4aqwy7rT2iytWWHz39czacjN+304tc/gY72niNqGYJtnkIZuS
z6ei2pxDHvZ+hcJwL/5hlTApVfNHuqeW4u2+9iGh+ZToDL2t22mn+Lj72W8dRWJgzb5u28etVtnQ
ht7j7iVrcv5qopb1KZai6E1xQLmweJH7WsXGWuCUJ8voKZBLSN+0JxzDOZIWKBZk/3pLpJAiw+AW
M1Z4Y6LI5HfENlCLQ+TXtk7ROoiTx2xE9/H8+pLIazi2wVbpPBn+v2t6I6Etz1bwaoXInWR/tfuF
qIP0932aFNrzoH0oGJMmoxkebCgaJ9YslBSWnXOjVmejIDQnki1BihbN4J2tyFtDdchNLLlRD3Px
hFpZMSghnZXINTe33q7u+oxg+GqL+5P3LaVEbY+bGftxiK/Vn35HERkkkLJpklKpXyd78cBDmfr1
FfSq3ogOGibVJboSoXsBSt/K+KSL8McPraLXzGmCZztwU5QTvrco+kThFFfGcI7Z5DW5ImMRGicl
QK5GpGCc7k9unEopBYdwo98Ac8jc6ymQ6QdKFFv4E6/F8pehRnXNrWvjWDDRdy2L5pQUjF9qyn7n
/20mmIccHgYK1+PApZO0f/ZBfZtSCzfzCXr1IIO1oIlaTmauUn2o38LCqe2O2KvMUOjqIrVjA4z7
xdwwahJguvVrKVnqJIHIpznTIw4M4fOro+WH60qdC5BvHYsB5XBQwQ+Ylj6kdydnUj/0yq4QcJiZ
pDavNA8DScgBNKazSusSXo2qhPIBzAbtwQ7hBZ0VfLW5Omo/VVpDYtddyiO0GwCR/TIC2M1SQZpz
qfUDS/R1u6pbCt8oNuRcBCtO/adFfaLL1MxmPD4t6lWEuJkqSq/ZW0GDBcWvqhCHanartptH4LPG
dkfCcK/YMXgKn+Qx1uiTXG1NTkdxjHqc9ETTaPBba2RYxi6BvFTe7BbqAN1utog6fV58NvosI5sS
rhJz9hF0OzB1RUyEPkvR0acpTEMujHwRSGuLzOsLKWgFwXrZELJ8XD5PCts7IEN5rTUpfaHAJjK2
aXfmq1Pi3Sb7BcZx12Q/lQAPyS6VjHWPpAJ2VHXv2cwoKaiAzKqH2sBfpolsgeWEwfv3buUA1QBs
pCm1CHPGWV5XjH4xBA5pbGUtHBrlTKRHUD1FPGrsnJyvwOlk4yWRCl+X/CHtM+pTetPdmxGwvOWt
6OLT8tIRSLLS2itphJRczNhuJ6HezL2c7yODQE2oYCaCG9nDKR3ZIoUb3BKsAi+brZ0fjzhOmbhx
95uE7ChDxd1PhkaT2ZXviuYg3SHtQn8X8R904JQvonEBmOk26Y74oteECqAWQQE68Wj0YZRbACL4
1z5mSRbZa/eg3uTm1ixY5Re3LlJyb7B6/i/IbRgP+r1Hu3QfOtjz91q7TJDudNUwlki0afpoQ1g8
9zRY7zxPlqfSAVvXxmQcLby9kfFhdzypP4Hp3BZlq+Kn2xo5Al0VlSxxuYLrYT3vCW9hNyj29Zxe
/eZR1yXQ4skECSNJFXJwgz5AhWybfzq7bcqcOa8YbfgT1yKkTMLCQwjNJH1ArJUsyZpL1On/k1dt
YjXReo0Woqko7oNTttfeChwaCAFQ+9uF7aCxZJ5fprRIuU/2wrwd8PDI0vx6o4FOqtb638KIYRL/
GORXhzSeNkD6jgO+9F/IMyO7uYA5en6V3419TkL7y+560f8EoeHWU8q2/OK7KOKFHOWwjMHkCU0C
wasIg1MhVS/9hivYVNrNYcZiHqJcILfuXsfeN41O04a6aEVqUo9ZQnKIFRiama7KSpTNtZ9flLd3
CVZ08ZSy1PMkiv8eP8Q56dcrJXRwmk8dJV7Kx0Y72bsJ3YAYtQHIHit2VDTbLQsTLwbn2dV5Nzn2
LcQU9cwxiI4yb89HBw5MPdOnzjYHL35UuvaQnAcDLJcy8Ab2QA8NxBFGA3o32xEulQCoVOvXatGx
1W04AMkb3ly75oEvngEsJai+Vp4acRmAP0Nz5PyBz7dq906BtuZl3QtheOiLpmAsVlfE1R6nCNMM
5lm9HRAm3rk+HlOgwBXF3wEyQ1JVvgBKU7xtTvFCmtqjhMgDkaiJKWyzq6qWp4RVSX7sUNxm2yfU
WmFiUxapqk6xsXINAV0BnBayNfSWcuO/UdWR7xszDyJpB67Y84WLycWkr7JhA+MNJXZAPhQ7WweE
zHhbZrY/6ZOw18haurrQvXzQDtPtXflExNMqJQiX34yDDEyi0itfDTNDIxikcTI9qfSHYFz4vKpt
6y8XCSXangTRuWVWZff+4IOsjk2MKYDaFhz/GpP52Ynzn2nFBRJmwnDX9lYQR7Sut3mtAllDq3GW
Y/o5wGlmMa3iHp+CW2+jDshX+nnw9NyUCwHxwDeXP/eIm5AMl8XjRzGcpkV/VVzt+mcTzDi3q336
ERokjEKQbeMpj530KliD7osPXC33lnOOhH4aIHVVTjXNnmWVQUdhSsFv+9mkU6bIW0oIsP/4FMhW
JWv69aUxASGaWeQXJRYW57ZIIzdmsj21+1de5NN8piXln9fdGDMpcDp0gA9uXgUpbJMS95HkPpNo
Afx6JyYdF/rf9igBtZp1X+haCsaWldnGfGpTLjDzsigePnxSgyPLDWL55VbCvgXm8fQXyaEH6nj5
o69RKvtvzx8mm7ApjIBRl5+jGt1pYOvlw9fI1s8Ikb+vJZRYSb5hVgSV6reDYNVe2RTLOqPKGMqJ
3DHWZx2//qmoqjLgOc2lUJ2WDeCCtzcug8dzH3k12sYFb/+COuu9kr2Blk/pWisUN26zEe6S7PCa
p2f6zEb3GuQlHyzu56iTVgxAqHBRZ8zJdmLHFdo+N+D5caF7PrMlczSALXVinPeTX4d6cgVbCklv
3FhsT2Ku+piKb0B4T8MBYNFchd3aUa1/rVvde5m9oqtEFaekV5wrDnCOqLuGqjETUozNS6DNXhVp
jOlAQCdvbsX8B0l6Naegvz8x8DnTmUJxfuvz07rr+ZzogVQUj+YIycK6hhT/3mc+ah+2nktcQuBP
+o9UC/MUc+9wQNPUGRQT4JaQD79KDMxARyJlDOHqdX61GS265NsJfVMsGgpDbborAUs+Sr4OZV2w
Bs+uWwSnPoc3FFzc/CBAEvc6GC9QNBIwvGKu+VNMVoDdOPh1DNRrcsWNHW+uoiQLBrZQOJZGma6t
u474z5L6A5N+tkqK+SKvwoEUHF9dnemhh2rv2fsRx3AQLyWe5srjN+3xVZNXZC1B2Fek+wqQb1X0
y0iws14EaJtlZXoMfcLTgEUv730tOKlgMZRdwkzwlB2yuwvYv49WV/NBbrx2aD/kpwf11F6QPA8G
w0UY/p1La1aIFW0qCxDQmmTcbLwMe76NaTC1TQBUE80pm4Z2Kpx3WhwmewTGlM+1y1jN/TpRBp5m
S93Rb23Lz3PY8N4IzGXU+W+J1rLbCgSVr85zg64eTaKq6tZ0JwcZ4AGhCTbvBT28zV0tFhBJ0eW+
jUfZVm3SrmyKcZYge+2OYLyd4PPsDBwNNOVv0ezrYWosjONjlsDkwrI74h3iLTWWHlbFyBRn442w
SIFugpTDALD9bL4OknPA5wGKpgEf0IhwFR3NOQAa3VNhUmnmHhk8WT8uPrCMrIA6qv8M3unawG9F
WgPSI596/1/OCIRJcHGTyYsl+rNpfKseuQYejsZ6b0eT0OM5xJEGn97jRbm0AxnHzdVILlU5HJOM
8JuWolUxkcUVbcCDmzj/f82b2rmaXVOvRYGx/jAx01vkgPDBxXOX5cN4Mxdj/3+CTClAENWlTgnv
XSi5aFuVVmADEeU6N8hEjuHUr9T9oREQuFkxrMwVkHBtzGPZrmd2pAPAOxJHVJ3P7E+yM5R7QaXS
m+wORkI7JEEY0VjHv6ZutgVUo9dHNRMKfgx7SlrG+tzjRth3ERp6hhiw6B5pXHiseCdKkhf8CibA
PBHLqYxc1lMrSSDMw3AzOKQ9qcHn3ORugdV+oNbK/I7MWqq/0tHYeupXbkhkv5V0hVZJfn7KSQZm
lAYD4HDXoRr+2KK6WhAIAY5QEGx2xsg3N93mA9ViF/T5K+BBwFfTCFvx5FcV11xfL9zs/YbtD3tl
vMayy/7fsrcQekx86ZAm5ZHF2SoVYPyTy5K8LcVg0Inno0oW+5D+7fQsCEQmJ0rzR+aaMaDgYwUv
BprvfBlu0Fzrn/w/uK6BcXKlasKbpzXgJo6KbR1FhegKSgwUO08LOpqYzJHexGlbHnDY36pEJCLO
stjvDYBFKBryo5/mFe8P+U2KkGW7yV88zFShAia4+iDvTX7xHaoAUDC3CJaSbC4Kz6XKgX4WVFwV
Qu7gW2bABvU/xZ/Y5oyzMZq65ELJ2YncMQFKUXcjkTJFlHD+Zc2tavS00wgYH6Yqk5cDSx4CLL2M
EANSuHv8HkkgSGIRvwgw+E5XvAuZq2sOcqv2ULERpT5G1VBuEg2R/dFDwQ2Vbizu16TdmGcEUGMY
91Ch5EwDKTm4oH8CL6PyVPEYimfK1aXk0aUmj9BOnvzXAVIgD/8SrTBjvA/GG8IwfdScd25yX7Yu
h4gDqOgedFxa4bISz+6WcQK/fpbcLUvsyKVG0oPEyWk3XqoGwh8FO19Ha6ascAAvvGLQz+tM4CFv
bzjyDK1G7QDDGiFvUZ5dha8TO6gL4rM8Qt6aUIHCxcojW7laCfPVUGA80YXGCfiO2uVTA1v8ffXb
uA8loP+NGkcRtEhZAKP0DmsVqeaSGS1vqPv3PhT3mcbK6ZF9ZpkOScVN1YrjNeN/CDYMvDvbinP6
BbZ0m9MQF+92DCNUjttYiB/mpZKojWN8xB5iuP/8x/XwebHV3rT6w16dUBUQCJbPmLxHHJgiARGv
4+KZG6viZKlK6TGk3NP6HdrP9HSf4Ma48l1dOnVRU98ISgfDEWaOLlBs9URxLYewVQpJ0dnx4D70
XkHqfez8YhEse1U/8/OJ+DoG+0xbXfMV961qKtsIRsXOoRBIK5qIllcc2gxfs3gbrxFKFJ+Ccqpr
+UoRRACH8CwEW0K9a8NeT6eXwqZB8AUX59uK7jFv+I5Y/Iq5K8S09VbdevbC6g7LQSBAQh8ZFJkZ
3CrZthx3QtTdz2NbJZpJd98vp7GlbbF5Ba1Da2ncuLFO/DhVRKboArZAC72jTrfyIaQjepVI4zrF
M1xUHDQLsEA2Z2AR2vpqUHZ30WW7eB6ATxA75OrOmVLOzbqLYhG+e/I/CZFQ39VdM2YxxBpMTTtS
B2+37OCDmN3C32cvnbMxbhYu1LuEKmAE2KAvY2p0DED9P1d0HSul8A0uHDbr0l4YX3ImxvdXtotI
JN1gzkWjXw3UGqyxrzw5vt9Y7i1AGqsNiUCAG90+POqAqDjXe4q3IZKZaEutOv30dLybT5cdFivS
gbQLGSVbpxw4Rd3U0GlkXO2GDkGOdrKr+P3SyxkKIdkX7/Q4ILe5BJFCPw3nvqQY5uFgAGLdR6ro
xiDoLYUxDw3O3rl6GFN0/GHsUyA95S1g8sZ2E+233q9xyZO9dLb1lOOySw50JDt9JFmgru1wtBMl
0o8mKLpa/1fVzrAvf5+HSPhF1dh6NG6I7ECUOuDOSTIQmapLtDp9I1VLw2s+DOJjphjOKvUswDlN
IjO01enbEs7UAhO5E0/fD3hgOrghBLMokroW84rqg9pNRQ4RIlWCCQ5jMNDiAk95nBUJ/STgIvX8
+sPC8fPfayhY3d2dRw830nphU1RE94HpP86PCamBwXUATEzTtFXikkT/4lReuqsNgS8ZPXA5VmL2
A55b5KccVh0odndc7it887RZHQ1hI8CXZQ3EcBuD78+ANbYUPFVY447AbUV/X9DP2Pi2yUA1ztEJ
2qSgXGDGbf0Q4ED8kzjRsfDAT9iV5kOIAlG+QsRpvmsAru0pvvcrZu4TwCvFYrIPBeFJ551OD5UF
CVLjuaIxL6qfCuTGvj14Nsd83xCji4p3G7rUGLcI0Pm3ftvm/w7MB/NHb1T+F9ubFcfniKjdsbXk
swUFLuCN2bFZtzlBMC9eZq8lx/Dpl10CVrmmcq6j22IMouxjCOQhNhq9TtN7o12sMfztv0JHy9if
GWx4v7RUZUCxDun027zSf83nX1GRhl+tEqnEmtlJCIEMwVRr3IcMXi82LD0/vl3FVx0SVTi7vsqh
5GV2vv4Lk2fVg4GMfx7AfFpbm6eh8fDjuGGedYSpCLTTRhBD0W4eBckr+Jg1C66fRnNj8HX6MJOm
blHzenQf6BEpCla3z/EK4h8SDlWbYULBRPD5Yohgwe+EDfqiWMzcHfPHMTi/eTWpwpqYCjXYqWqN
1N/gp2yI3+F2kQgHH+eU6SeftMmFQrgJHd2HYdxkcPnJp8m45Y3+NCKyWyyTsaVt+tUnbJuWZQid
SUV0BCRRb6tBQnj4d+vn2VN9LdAZWKIT1HtsGvrwBQVkbmIBbVlGM1Zk7JMdtSibPtlYkVwzByMF
Dg5GMxe72fX6EyfTKWiXbAOOo9FD9X0+ia0eo/iTiI6ftGgBlpYMXCDr018Bk1XdCpGO5nI67/Q4
Vzy6ud2h15a1PO4shN1awZ4yWrqsJ7LQZewOJhY9i4nnogCUYxckvBPDWkeNbZDEc63UIIQrL6Iq
iS9ev2C962xileM7XovGRdgM5JOsAOfMR+r6nSFBhAR91D/ZPqX9Bwa4V2IiBwzNrbKVJtkPTBiJ
G3XPCTukJaxazA17wjJ+WbNDCikd9MnsKk0D0ZQPxumut94+4XRWbBO/OF6qEMVYACj6oXvoN/YA
rEzCk9zCsIk5umqnqB0dh7MAkycbl/5oPgVUv+iNm0p+RZegW9FGUvn9h0aPXMPMnnj4jReIP23f
pLC5UFk9CnmJcMu3TmiT9nneWESvsZelGlDnM7SPhBFXkeu/lLK9F8PykgkE5s5RnhWBkObWE8Pp
ck4rhr5X/mjRqBY6KAWdsa/bfqp4tf3JIHxLdzY/USwJn7u2DAnsjZW7nSMwqfVOt2CAYNvrfH1o
rvQvekamCecsR0mGhT5tLbfavmVxYT49w8U5rfo8WB7mJC739dCe4v92BOketQ3wjQNumRqzrqtT
04pk8XC7NwhddDrvNy+W6slOlITu6uxMDKAblrkXxmdIiTNX7vn1yk15m4ZcjxcMfYGkeJDTVHEY
BeHILmcvPMx3FJbG31eSs8CSm/8RfQ0gqxg42ypQkegmkiLDDCdVaYKYoNZvhf0RR2Q+q4xqGnID
twRGAh8So7S0E2AyDA8m8r2mxx/mram1Bf9/IrwI9IeZEMiOv3cH9pksw/ovNLiu8WyWe/uNl6L0
EUNHJ40NZ9EKYA5CBsp/0LfCiiSoQRrcoN8f0CoiA4ICX0S7fJDNcZqiKNhvwzsT8bohPhLR7px2
c1aDwpyleE+DzvANpasPcndMn1llvaBjeJxdNetZZraRaC2Q2TzfWDsX0m9d8cEoGNzGrTrnhtxA
9OADzBBd2/DsKgTeh62me3iNxf8SdzbgFhoiAndyXYn8mMwveUnE0I5V0mwa25tdtsHBtg24fHZj
rN1eELCrHSg3cSW3F9gPxZUffiHayzDGdqhf1YN9kil7kmbn1KcwQHqVmhX853p86l31ZLppJ+X2
sVAL5IQnfmAsVyzAeojihtralwbTTqzK+X2g39dceDH+lOLT7vRZzj96DhLPNV0wQqtV0xiTin7B
ka8jbhGYI2lOpl/HiyACT7hPuuL3OQTJOXPRlrKPWYayXDPI3l6P24SsxI4zIU1nI9QURH/Y2DA2
J4AW6LNPaxAZt5T8WCprlp90fuL0l4X+63mJ7mE8q+b1qTc8NmcD4X99mPtl3b+MAu0BTyZxVWy5
S477bn6k5SA/XM4YyV6HL53kMEov6F4gyz0Y+X/YLdLhOpKUm/CPv1poS464u9uNphySxAkeWE2I
APM1/uzH9rkkAMorKz6JftohdAo9gXHK79SsX7yGe7SUIah5pZx9a/cJIA6fVrc/ZzdzIQkvziNu
5ztNEg/MMF7xmkr/MSIZFaRLsGgzjxx0/6+eCwFubFMBTLiMfmIziArvlnRPADyHbpsAw6SpINFo
9IN++UojkxkvveRE8RM76YAqSaZ1is6jQKZij1IKTCDm+t/4MykMFvNfkE2M5pqCFwpzgDAuY4yj
xfjBlBjUEGclPJprjT51DuqXhYoADov6mBQOKvat2gEBbNalP3u0n3EVCSGkuQ2oW+EPMlC6/zwc
ol282W6J2ZrKd9sTohppd5a6IzBILLmBeLOCEkmYREUfP3+Slm3Wdr0WioBWXePVMkyGu8+5eB4H
tVose5gtyc6TvVsB/hNYAm0tkz1G79YJh1fbjnXG5s8Ty1MWznoi8jlFTnL9Dflf6bq2pVluiJmE
h2TFz8xuOSGuMgIUQGsVdudX9DUZ/eV7ke8NyvNDol2EH0YuBPRewghzRDRarihsS7SncQ6rB58G
ae1O0IM1fzAU2rUh8Z4AgIxOXNEwnw/ET4MNUyFwmO4+WqWwjdotwFw9n8U5JK15qQpsO2n8r5kO
5VokQqkmrermuUM5MmyVL8e/h8kxGHggGN6Unr+Dn8l+8qgMOo685m8AnyeLFDplM8MGXbU8CXm7
5gMbAVHzP+gVSt05SByCKLjop7UpeznZf7s7NCOv3fkuPfXk7xEIDFRCysRlMPTBjb5MT5fgvEiA
89SsnkGwtxFtwhFG+/FxXw18GEwnSkCNCLNY1k10TTZT5BHgZlJNvGn/F3WTL1vTGJmZNt7FpcNS
U6S0gQgB2BKTQoi5SQWcHWzdgcMg7z6+e6p/EBCO8S7Udl1bVmkm1IYR+pV0lOsb6pHRuvU7y/Du
WRF34wAlTyBVD5PkWE1iIIObQZWI7X49Dae2gtLxdTc90r8ecv6AY4zn5/2XW6SlWqcTL8inUPNl
5A8ET0EXcMjzgJuowvXXxNvvC5rUk4dCIAq/42pDNciQJObkKcHfTxjyFf9Dgj+oESw3mxyO8/OT
rIcj3sjjvBwUlTv0NaQfGe1Veg1/y9/WKJQxDYkYQfr0xiC1ef/U+0p4EWNsrJFYOKsKTWFZGHOa
OWAJcajAfvYvxF2jDW8jGpvR/1FVUG4FXN1gWV99HirRJCwh8uYzhBSfRld1v5P9fVnNn9iRKuCT
HqBuGL3b6YPKB29p3SbKrQwTHoekR+zZo0uz8Z6X/nWsFxG4u3tIzWd4g7d/9Ct9oBHhdeSWmlpQ
2eikknfTC/2zjtFcA9MW7HRua7AMI64zIwYtjcCSeyZZRhn/O4mTwYhIBrfcl9GWSVEzd6x05QeL
A56eQck5aqPq2nhxSbaXYHXc3z5US2IP5Cdp1tOShjs5rk3mf4YZlwEvXujPpxd5ShfQUp6tMAeh
Ua05AoQWhdTL7Fq+6KFkTZCOnPYLNgdsWMgzUsMzGrbR1eOEXFPi0cavkoU5zBx1KdwfxAFhuOk3
4XmvpXAa3K2oXY3yf78P3g5Y29ykdh40HoRxa0IQYgvEO2AC11k6N+oNgvFcVk51IfVjyqNb14nt
c8m6HjBDsTJqYt1u2aPyGX43kXJ9gUjctaJDX4r2hP2UnFX1uCXaGFjaIpnhIIPT7oa0mxa5uQFR
rUERJMBLG3rmj0rWnEuemeMnXkCQOKGvnfQuztHc+ZkgAeWR9HdEiHHbakpMcbjJv+6G3T3LYf3b
I/Pac0nyaZD9XedS/0MZAmMVuKgsLqvWYWd/eLGIzxgrb19bQ7o4qSh7nXZVgsDpzHAY2RZqpcDK
LWI8phDUXtcciKH9gN97T1AdRVnnzfry3V025LYp4C1CLN+nnW5WSAJ53/Jn0GinOLdmuDQ1WTfK
S7UusS15iFakmIcVQp/oHqSA7UKC8DbEHeAOPzvXTBIhfChPf0/Qo/0Z5wp3dYSr0mJ0RwODYQjL
3+mvHdPvDv0j5pzTBjMAGCFXFbAGPvesyKDaobsdfx0Sbzek0zA+b3639zzyvZeFGTtdp6fdP3hv
rSE6Ez5ayf/x5NUhATka2orURS0AYaI92h3leoLV684998gTBrSj3vI2x708AprIzfdOgEtJANsL
Q21SSAixmGG32Ev76i+bCkfoZkuI5cN/ZzKSYqKo86aIbDub4vcLTecJ9/uOfx9+UuyZccxxBi6C
COr9IWDsqeEYRdHCcoots0fjUuwN2ow1dNfg30eN1sEZ78I0g/l7z9ytAsAKI07TnVEj0Xj7Fiyv
L4buxaLf2aE4EX05cDoX2tZ9R41E+f+/zDaCKNBxuetcYlAloG33b7otDUCfEpA+QwltWusasS2J
tPShlTN9/hoOArwHfaxGq5xlWmerf8HeVqK3Oi0QSFW7dB00WOABQgUgskOaqRCAhxyhJffmSMJG
WMKe+issoE/fX4e1EtduGOVHCPYkpdP3fMqIDvfdAKAijI1cB/lYO2+4PBrI8OuUWI7WK1IJqZ74
/lb5vriHPgg3bOfKznL0Vc9UoOQDndPOOHj53Efw9B/FKghgu8x7qzzDSJTfhIoYcKrMkPndVw6A
M9HujwWvxL4c/SZ/Yqs0GrnZCBV4qCmThnJC5xbu6NRegll6JtRgFA1hkSf4oMr6USCmGTbv5QgA
to9fq92rxCfvILLGIv4PtDoYjFtHdqOipH3XnbgWPmwoh6RHbQXyfaS/Z8nOr/OweHIP3EayCNn8
i0vqnyHTpPzqMRSoHpGTDm97DO1iJz2DCvCp/KQsqG0PPtB+0kT0W1xjYacZrrpAavyldc+lThgE
6WAgzTutOqvLdEUNuszdzjnRsQYd3vrsvfhP+3g0oxFXO1pJPFBHjfpMqAdyh1aogLA51vnv96Ic
GjfgwhK/3HQ5+1DXLa8LH3RXcm8C95VGbajNsG1u6sWa3ySmyLGh5EEhXf4FQM0fBQzXqcwlMAKg
qOF15tSrAwBV6TmI0+u4YOOxrOOqC5KNGegZ98w02+F+5m3FbgaGPUuL/vRnBK6AZBVslVUguaXy
VUJtm49lS/f2H6p4Kjorn46hbDKTnHMkuc/rHZvc4qIqOuPhHYpq2AjnMw6jT0Wcm3B7J4HbQHvf
rbCFQmRrWxiX39fh9+vsmkW0u4oOK5yLzfTf1why04/JI2H7rj+Itrqv84DuJggK1nI72CXHToPu
sziBDgNl7QKtsMEK3gi046ahX48fE/l/gjqX0xesE0pLFpQit/eIplwyLehCym5WdKOzg1XGcudR
jlnc8/argWV3owxrsHDGlSIsFvRiC/mmJXUwi0G3uB8qPezO4WqSpcAHdSiYQ7kcuxd3KRweg6p/
6STpcwEdii0A70mo3UFY65aJblEC2FrYEh4iSPeMzT2Dr5IRnP2Tn1GYVwJg79PjkbHCV+1IrFLw
JTajmwdziLXqK7VMFMss56b1CCxl5xr6hiJfqpevu717HXjkCXo4oWgndfnNZJTbcZT+MMi5FjJh
uqmbln/QchT/kAibWYyqFqmNnO8je/KV/3W7V2TlCQIrTFAAyjg7LMDi/Q7shEV0fip0JGRts6xO
hg2ewlSnQQzrgwSoLp358afumDYSfcJ4jSizYe4g278V7PUmAO+PR9DrWSY6pQGxUlI+CfW0Lkmy
+eLQgVs4IqjPQAk5JGHnKouGnwId48M3B3LZ35JBOtsg8P4tq4Hn3GL76+GcT6G/AArvb+BKIZc7
LEeSYJqEUWDiefXiGHxCav1vad03R6tozOq0YDXSMLjcJ6OkJNl19iCPhbDYSRCcFq9fChipGv59
fjlKkb12y3OWJaIBMxZaniZnk+1RO5bWWSrukr+x5/lqUbATd+WiTvTRyaq0/XQVZdKElziBpXZP
o6s5DreuzClq+0fxDlkzv5OhCOfOHWDM2gfLOYIBAVnKx1ULdx6pGlgjPd4Oh9l+VkgoYq9MMOqh
+fmPdjs7g3WypiSicPmMCjJZ6jk3GQun32bOaI7oMtRJhF9Bw+38M4Y8AiMARnjjti4Pg+6mGoOK
Zg+1LTZwdiE94XSIXtfxB/qcr7JOhqz2fsef0hl6wQ0d4suAkI7xlvdimNOO3I3qt2oFB0cRAl4s
e3e7tcGHWX4to1qEKVXcTgz+D+4i5A+jtf0BnEryeOOihVPITE64ne1qUmD7gjfYz0ADCrAUyy05
eL7PbAGSrtqCRg68aw8xalBujL4TOA7SYpfedb2b3bdGku+26JOp7sam5N4/jIQzVu3Ygbmtktpf
zYiwZ7xgaxkzFKEMaUIkVs9YU/G8pzWBmhECBdbsy3ERLmalbX3WpMFyYiOMCMlJbr3BYIYfbAW0
5DOt3wvLdUxnQlSSOSJfBr2o48laCaMysg1/tfT3tgtx2xBvo7+B7abfUw9I24FY3mgWpUnbWfk/
Os/qNjdBvbLkyYVlqxxZ+MntHNjkz1xd0Fdn1QGTZfVLp9Uz5wt3ZA7iTdf0oSbMRe68i300MnWa
2e6fvy36KDS18MjFDnfcqBW0+M3P0ByvL53W7rnyx7TvNVHm3PgvZ9Mwjtc1kFDXmAHpvOB6EXjU
rLiRCWNp/57ZNKoGMEqj2dzEfumFGqpS7Y6EEMwzQB34BPFgX/YYsS5GXQSFGJtyt5jrqDokmFJU
EZx2oJZqFMaoa3wphXWmNxc6vesOqKJ+FKZBCmKUtlcUy+mHqGPYerWMbkWxwmdaSSFciOELD+G0
9Ygu88j1GGJMLM27Dmynqaef68Hc/Tnzk2sQq85Dr0fsZxQUmRkUUFChZUByAr4XxUWIps+xge05
8E5lXrb6dcqJqbXHkVaMkl6eq5JuxB4kPWzqZ9um1A31Lb7c3Kj+N3KBLGRtT1ERPYno/EnBMdvP
3PGt1m+JsFwORSzJpv+3RksUbsqP06TlvFyHeicqripIkfnNBvdyBqJHbYlMmyuvhAJjFf8anMGo
Kj/VtDq+F44duPDbd+BxRgeXHc8wFeeZFZWwlHbJNuk/qGKqS/6+dvm95cRNFn1Gj5/yMXrzbRfQ
VKf7aWJTnJhsDG0JHjhgrRm7ZZfPK0Skj6huuiQnXWtEdRI2dnOXxOk1O/WZ97Qz8k5MRdMc6dJx
7lsIFen0IVjskVALkdY5RXvHng2U2oyTaWOeuNOMC/zWSEtQDuWmn1W0JqT51FOhQka63t/lxplK
cm9w3KeBwP7HxkDn7ORXVZnJ/pTeQ8xcAt8buXCNmVrRjWe7GRk4RysdXfucANyzDIzb16VVjBUA
8inc4obpslRjkHVQht2ezmH3zGfs2CxMWOKm7bZH6OCtCfOtElx0N8joze1mD7qutknZTVI+kjfX
Pe+/mkGmUs7+V5PpkNkO5CW8+ZRpj8Y22lzkfAV2UmLxb9HDSGeVMRry1lYALjabxtpS4TWHrRiI
LGGVXtxJzJ2DhDdu4VGE2Os5MqXCH2fBJgHEjSzodFpusIMlZCmY4j/LGxiRQwGGGSlyyWH0wjT/
Ht78qBtY4HU4l2b1fGiPgdfVTDJA8k7OYd9Of7YIkiSvzllIit+o6tAoscokxg4ew777ETlr7Ekh
rV8OHJT/wgEGF++PmvIaOwKtFiuLk+2mVVgBSHgZMl26Ll35Acv23mUUHYOge27uwDOdeltF+obF
yHy5LKxPa9pC7JvCSpQWeYerqGBnqJOwpXVA819UnFKrEdXOj4lBSVzznsIqjsELzn3A3LFROP+p
0XUHILdQG1HUwzLPIVLF25RWjNb14q+n6byuAd2FHL5jk7QY6pox59nvAmwfpCy11GV3O7Vy1OUb
ChW0x0Fj8ptZii5JdHxtCgW8qguY4+mvOcEWMGH2MnqdRVB3xk3Kw/3Q/OO3PrvBqpKGRM3wggph
NUSCmM0UH3Tk7h1pr866+IsGophzyuJ3msh0Nuy2ykGWn02xHCTfPvClE110CQXWp8V+TCxyt9lc
fsKziexgUQgpcYy0rP9Eop8d8/Bl7/ipuYuj2zLP88oNFZgyMgBsgb381N86LVN7+hokaMegxr9L
4n6o60Ug9oiamIQvmDdVUriCpwm0GnRvC3yZeBZWkOOokBZmnR574gMygLjGfA2QugFqVCX/KDuo
8z0opTMDtUGmR4mF4le5HtqwA9QfcyOOpjuUUBJlXYd9ycgxbgF7lOsvEsfIniWbPOrD2c4B1BIN
ydxAVeRsnAfvg+gJ0y8yKFxxJlfEJREfwq/xfS4SElmr4bgHiuMDVoCVANGptLzrRTQXJFP/7pfU
CVSU6BpFh2AgNB/3gzCNZ0K3V0R4KY3xLlIyWfNtFHVK2875QPWJdR1o7hpv+dTlfKl34Jaf4urD
VhBPWthlNSMC/PPJI3KbpAxw17bdxc0Pa7ye1Tq5UyFZ+GxkfsJbEjtTPkWltRvhklp3ftrUJ4RQ
411uJNNewS5Hyg/LVapCcoBYTon3hKyjsxM2ZZVlolmKcuawv7ftRBfDU4hjV07oPGC/fLdCkT3a
WAsZih9Ys1Ki7lPPfqNmwaS9ctnOVPwZn3ixVhiFKwC8guXJ7t/zbumvayjuL32ewXXUzWQrsr3F
pcLEFYV0MRrbaT5L5kllmzcg39p7n+i8hTQg3yX8xoJpaQOiYPOId5GEifci0YonVAUSKZ5uq+jc
vpgd3tQyf0oGlWLrWr9HfiUUC4JTWOth5jL8ej4mrvk173dzUvI0ylKNcICNZkq0NkxrhRYqljwc
k0tUWBuLcoCDBZDUmfLde28Z0B/5pBPIqcxzEXQ7PJ0NRPHlqp+Xp5SwdNUg0yvYEJr2uAaoJauh
HJpcccwCKCdQMAwM4spvTmpsjSCaDms8FGRFbQX4LUl9jJhhR4yeeiyJYoYW8dg+qRdx8Rl7k0BA
d1CAPu31krRQVwE9QNgSBmK4hUO5q3PS33TZApeQW3zJuDnpNhQFcG+tRAPDh3HVszuHLCYwe+qB
9IqXqxxZ/bEYsa6uLDBsErl9q58EHkOD+jSqPMRaoaR5g1XtPVctv2JPJvxp8oBAT9fmtLFbRwVa
yO28vtjt3vcHG03A3nePHDnP0Pq/PyyMuilnf0qXpf4FAPgs2tsijCNIhMA/7b5pxJKYPTjnpIFR
fiI/EMXas/NwHTvd+5jtnQfJD2Fh51mwad0vOx/iz7+iEKMrof98NNB8bvgEbknApWJU1LHNZf5H
TALywMWp3Ef9OzXGAcqAZuoEdSpdJ66vTydcswseD1KozOuvq03per87p6TFHQIF8O4olDaNwyY4
1uJcxQPyXLBJVqVMs3FRPAjQ5+/WYOHQ+snppZQeVlFu6fWKjv4a40HhfYjQYpPQ+3/ZkQcnfcXT
eeFIqWiywJjwdRt8c3qKjoHV2leRlcz4iwc1L407QWJo20AMHIG353JRV4kBm+S5Jr9BmKKqqkF5
nznDQ4htHV87wqm4owLeQmOGplSfKGtd5Mg6bSfJ/FheBUYkmz4SGnZFczIJGAaLjClCFW4qtrNY
hRmPPbj+12x0pptclyVAhPKMN9eBMUCx0cR8z8ledbTHhDnz1/DJ9MWuOHxDLK7WABoDPnV1QvDD
V46Z22kLIIccmHugjIYjhlbe2EevEP2B+VOzvXnsoxqnL7C3QoAIU3amOD0R559WT8CC6tdn9qZ7
2nM713lmAlCTjgy9qfHQ6zEWuRN4qyUZOkMh12adFpfFWPll0D9a4XW7o1dOlWGnutKLarquFvD+
j+2zhaLzj2P2oZAY6MIw5WDJNoR+bn5xaIRhiA5dKO/OZfhuYPZ9yv13grAkZHNyWqOssqfGSMyt
fcDVRLjiymqq6zaVTNZq4JnWbh6I5+noDJ0KAlCc8UQZNM3zmU4H6yf//KfZXzVKshFgzXndx+My
2RmvVv7NESUaxcQDlzpTlUE913qpMLS3PCRb3ZLLAp2V7lPT915T/L8ksUaKl4YvFkcfdQPA4dwf
hUfI+Pik8MOvaUNv2IC8YHqh/sIuRqO2GT6zU5lAlwWutgYAKEmlhRnilX1kb160Aeuoq+no8or5
BRehASVna83gpcKxHr1TnBfABpCD/C2cfMQMnmFZTWo8X/I0GUeVDNSrBNAFmmXVQycxoBIWDZs3
3nV0el6wlNGhPFMLtHFbezr5a5gtf+vbyU3Gf9mA0qeF/HR6qksRlMFijx72O7EJeRp8qa+mxK0C
QkOEXmspqf2FFvitDQyo3/skf9whlL7HYPvlJw35h6I+JAZm3gJrEnT5VjyTyZkQMMRVqPPLIQ0U
D7vuPSylI1gmvYGYd1iVUxbkjCVrApacJP04Tn2IvAEMNcCdCyCdkEYpbRRqYY5pn6KYAckvmIRa
y82J1QQAOS8zLDhgsd3FS8ZaImD9ijW78QqS/5dFULb2VIzCoDP5+9fPcyEWWypT5MZnAWQX8Vkp
+8bG8LHyZqLh1fgg3wkGEORRwWgHjZGDt52ThzYkGctRHj2JWD+FF3v9P9ZqQNIcjBxtW8FBzV9c
6LZZTPNciMvMyB2anjBLn4yMt3pto3+qDoH+pDKG39kEIwfpq5LkP+tcT1z9eMTq+y+UFiaUR9c2
k6rpwwSeC5wSddGfqk+I26YL/3Li9kig1BYAV4H4QD50tSmKrGKTviy4Lw7W47wpg2iMZvG8hX9x
EBEBsJjXsoiO1Om3y+EqyPOpvVsDnjdlMvt7XGG6Bk6+MRyiSTz/4YC+0XDgbvV4t645O5iS5Ae9
qSoDPmlH+8ZSu2ppxybit2pHqi2EO8VUjEEvUWcv5TePRwDqtdNas015p0GrLt5KGtcNf34DkCc2
eiRUHA+L+3AUkmXZAU4gWT5rRjmEGI4QTQEn4yMDClO7BxXSAkSs+lkoFCr2fDR5GpSoRr4IxwpO
DbTTRfoD7iGMN1vdoHV5+t82QrOfP1ex3YiODSO+bNShpAs3TMJlLpqyq3Om56izsUvXJyFc8A6U
PfFCAaZTNdRlhKqwWjwcUnCtzoUykoq1r8RPkT4hP8QoRv1IkM0xBjHB1FnP+8/QCyY/KNMVDjrU
7OQYCTRmGnMolYJsseVUtkPPKe0Rojswk9a9wxVZsPBt7U909W/pYvjs5CQDgXxyjh36xeYobF6c
FD/gZMWjwTIRcOMxz0yRAux/LdJ4ypEVcELK3+bMZ0ywsVzX5fSPLLaJKm4cBRQXP7TxHtO2yOKO
DffD3Ef4ApLhYd+Z8yBYpUUU94EtDYLmOnkQFN2V9omlqj0zazP5Cam/oP/AU+7DZzbqZZQLMaWg
2RDakbM/zND3ZjkXIgOMw5E3omKG29syfSt+vxm31qy+bmXAU5w2UPr5mPTyDsxDtZ+7MG6WnOv/
nWlItSoF5Ktm9HO282SRR18VoT1FRNjusNf1TGkkBSPzk92tHqX81jA2b57lKE8VcMLtDChDftqF
vTLuUEeyUyVHFBDkC9GObSyPvfwpk7Qoktd/dCbGlMcDqvtAOnOuqtfD50m0uMYmIFH1T2mXKc4k
wUQszwH2LDXBcr5qf/jiLS5XyLW1bpVbQgfs7JK74pZ2ZWVk40Lp/CAStEe3wVFL2qnZheOcwTZt
IIIm8euUh5/vhfaSFlBUJse/p18g1XUJyfzAt2uDtRUwgVZjUgpjvl4PLdaotYTxvaHoYzPHgazY
DWTV0teXo/YW16EwFUzFTQJGIFQfYEXZ6tlzG6qreRhV1V3BnbkxECt9jNJjYJIcZvTNdo/ln2cS
kbrQXWgp1q80/f1b5mjHFwtG4X6+AT+s7Q2MgTJ7R9EA4nOnRgDCCx6EpmJA0heolk3Ji5AnN9hM
v/Lcvn0FxaoAjd9N6C6Wp5buL16FNtAZfhtPk/hCsXdIhQWlSvEX/xoX4St6/xOra1/NTQPLINx1
lQYBmoXp9Ap37aGm6QUM6cCxAYIYwTxsw24lhBb1aRwuc5/BITBs0q5SysuLF/jUHlOGW6eYgzRt
gG0e2W9+M9caw6FIsgiPap5N+76+ttHCR9L9em+Em95QjIPnrAWpg7e7fd2q6prmqdxogBFjuBSv
Xbf6UehyWJrtSMkf+hiFsFfcoUwgfgV65EtoCZpB13TOC32OusgTtk6xossYhAOnr8vaNF5dUVXj
Xop/NVKAN43tf8kXC8R/23WniWqVcDTjxv/c7R3gYXr2DBDtsLuSIUvH0tnLF0WCM6gWq+HhC916
IIeHcFFMCtfYueUWJ4Z9IkXvRZ5XbZtfWwdGPSxHH3JCh7cYLOvx0VkinEQo2gx2EoY0FHKSfwt/
QZmwI8mgrnDc3lb85KdnQUyf8g6fosGaOe3wtqKp3OJ6RDTUc0/ZLAR1fe6E2djQTRp1H7y1gMB1
ih60GhfOdL5kqJizlZY8a0Bot4YLgtpU/+jdM6A4dtezDsjpNOX2lyGk+GwI/ji2yORkAeYPj8Gf
uN5i9+yiyO+32ChuePuyTJ2sBos4yYcIqtVdN8EyB3bFBuiLCiLE/TSEQw0G03xWcsqTjcH11LHj
FgcxIsS6QwpAk+lVjJgbeLsLPCFeiY7I9e9DlU1f616b9ppcewnTzRybNm7rIouQLjFD/0Xo830O
lsCJ0OFlSCQzidrARLEpdrCMUyg3iYc2geFhdOwhlbwrkiustxrpod3LfJcoFgghEf0AAyxQa8jg
FCWydv712O+kM8BnNdDmHR4jgZaKoJDXy8Lt0AvqsyvCfvSO4XrguHSxz5IED9GRh9uIT4oVHvGZ
fiTwYZw+jnSjtZxbTCvrEYnSD4ZVxPdSQBX2sVKwUzD506goBqVUAtlyK7Z3ECNlBUpCQEZz7xTv
swa4+L/wzXGXTqMTAaqpW95p8sT6+J7YQS1Mu+Dl+R/xuKxE6f25/rTaPCO5+DRX2cqkdM4Y1lo7
JNaV1/P02qCNvnlOTU5SvLTsNFrCYb7C9jPPGJggadWvGCm1m6EsA8TnrFS0XPCtP4B+2oYsWk7X
J7MHZihHfiwdDLqkDfd5aNemOgiqg1hjImkIZedOcJhhAFUF8wdX4Wx6S5J5+Y/laZW7W2WqZh3Z
DXHuzFva4IWXwaR9hbNm5iMFHWDX2GKwCbNxN/fvOL0L+yUEX4D6SjyZ13HO01RQJj11FyhwZW8P
cMVI9rhbiK261elVpo/qVWr5p4TCpeQ/YF0vUy+zdGJ9+IDJ2PHg/NSDAPEGySCK90N65RZHRhVp
DTRyremNtWMbup4du4+y6q78ghB2o+7bUNztS0im3LrWh+29beC1LW5dFUIr9F1hNk1q7dA1YNHx
DQlMO2btYx2/dfFrOZmtElBI8MoxNPhqVCA/PEVqE1n9QccJN0whJ8GIupP9D4pIAsesOmrXozX1
DFXj1UJnSXeLEI7LbNC9P74Unmq6FL+ZNL2+vMYMTH9RSjuXSHynUTuw2ep/ZHrdLs6h93j0o+oe
k9VJb82uaMcX9SkNOg0/Tk+oOi+nzOt+/FsM3xDo4jSoEpxoExNge3qt+RCsqj8jujQ/w/yk7O0T
NWoNiQ2nONtLUgv4sd2wFC8cOCfol/YhpHR/seiorZXzeHKL7di87WahcgQ3ZgH4AHESj8qJcMFm
5XXGyCvXSk9Smqw4q8Q7kX9rzvSSQS12CaxKlR5AJEch/jOGUc7Nnl1dPKwjm1vjUznxjmQuSUBi
fRA0gAflB8zzryKNNTgunMS0pj7otAHigBty7GysCW0NgrhAKfkZUnQoE8Vx2E56zHBPJZ/ud+1d
yAnHHfw4jg7V2rINVgoIkwHI3grxSH8TwA45q0W7dvyZfBR3XWlk5waqcYS1F6Qo4OpTZ5ONG4sD
eaP85mpivIxCu8A2kTuxDDJOKFypab31E0QXfcH06amOMBGcaNCKO38TMPBvPGhZjoEZaJewyARZ
ZcvY2IW8PLX/Sgu+0o8ClvkSM5Fwim2RLM5bw3XZw3PgR2wC8St8f7tjxc8420BxsB5u7qyFzUp+
wqG7bkRflcUoGKnWaqyMgH0Qz2ZBQS5tE0hLO4Gg+JfqrTYtYYdY9KeOw3tVg1deK57ifrlmcGBZ
BCWGOfnzL5SM7J7tuXQe8XmZyLWk4tUAQPEkj84ZHyD5QKJJbkCz1ykX90+s6e1pLPeYA++bJ/5i
B14J8tJx64oPoYdO484Ju+Fqijtu3bPKGFTzELvCysm+RgMcomKpsL//+scNiXoLUep+s8Cy97rj
c8CMI9CZd40bLOasoKFsm4L9v6ZOw/F6+Oc0RmWWXqBhqEXJ/nK8YvCkvxP4kq7+48qwUENM2G5+
arroyWEVOORK37pSy9ASnnzCJbs7OysGVvfMLl1gZdT41qF8Fhhict0NekcoCiv+ULBLb2RD3GSM
WDREJNsr3ahCsR9J90mA6swD+G2FcBf7B2/sWCgNpvrMwK91gcho9znok5b90rzcwAXLlzCdHda6
AqSpHNeou5LMk0M+scuK5CkryU+KsAcqmhF6zZ6Z885EkfSbboI+z/r6O3w24qLfKiTDZQ4nsGhW
S+pcntEjy0SN1DsaQfo6tNiqy6PSI52mpet9yiYcIU2vTp9QdtmejL11JlL7uAJ2a2sYaWCwvqYL
AkpFgvQI3Y/g5nvoet4b3OjymDbK6ZHzkF4yg2FTpcP1mo5wJzJBJheqWuTMXk6/E+/DG7UCld8z
uf4r/lHL2am6I2OzRoWMzppvchT/Gl0iPzPvbOAO1rS5rIacUauaSJpSxYXx1gDbKGMFtcKVCKYI
520DcjmURiCXrufxPVTNSdqV/EW3WzUw0S9cMp+M3Ygs1CiBic8T3TNoR8ZLmHT7YVdQMMmOv8Nd
8wegIsO4D0HpPXmW5R7M2vXpNFn7DkUsWOrVeC/3eaze10Hijg9F+vfVcLiWyT+3LuUYYwyk93ra
BMrmajn//8g1MVVGokcx9Cu8h6hDgQV/dfAFpTwiZphoc8av9r+h4E7m2Mb2ri1zH3AWRy+6tNJx
A71SwFDbZ1BnOwIPzDamouK1Etp/ZD9uPhKmBphOQIazj7wTpEgq6f5pdfI3apZSaBzvpG62gAjH
dshF55i+d1/ESnqau5rhNrRO3HIxt2n4ItkZkw8X9etAQIRJehTQr0Oao5s83JqErQ1lJePRJ96x
R1tXDKEhCJeBjshKUD+jY7SL51kENvfpTWli8+tAfi+l7QfE/t4bVFNYq8T18bwDlq4KNyeuurRm
B+bb5sEm0gzun+Ox6ZCep7aqkQ4EoVGtgXSawNI6WijGh+RKej8BSVgWpppDPAmcmfqLnqeyI2lK
jOmjiGRpqsgWt/crzxR/RrqhUlUnOe0mCbeGqXRZ2Z9MjYgjQ+qYFPDNKMF4kp0zyrlymrK8g1E5
LP15VfFhrSmAEHut1tw9Fa+vLT397gKvVVGubJI2wSikNlugDAuxwpLzV3XZhxWZwIh4okN4Wt+y
3IBil+I4i8dwQrQEE45x2N5ErPSRL1OLgwixV8V1kcq24hbmSABFxvWp1RcX/mSdcNzQ+q6nsBlg
rgV0yJEBsKemLq3Q4rCnyd2DoeC9ManAaloiFpilukgDj29bcqdTbm0Ic2jbysEtBhe6MvAUX977
Oqh9GUqT71vY36o/+LxKv7FD5eODx2LynQ97649EXeSYAnEIrK48OaXvRZ/pMmkwvPy3GVqrDWqA
WCFvxFfman5FbUhGx85fAgtIty+eikw9dr0B91ZlkS+qqUrYgSfZ9ieALKEq/2tLOICxBYT9rbOc
lYk1Hn+o8M4gxk1At5k2IWqIh83WXROfWTPYzTu7UZJdH/S/xVSxqfnNuGglH+22Cm7f1kdxiCeB
slwLtdNeUdS7DQz5O1ZhvdpwYW3hPTz5hoCiy9NltCfnXIIKmV9F5snmciuRhDENThqd7Q6zsQ0t
M45SRBawbIw6SliOELwrACnwSAczTOss8tB/YNw0H7bw7gaAL/O7ZPcCz817ONtyHEHyaHRFl4ET
V5K+1w87jYscGPuemhOpBrNLPuY6p6wnCr6Q+6bhLgGzBXFc/krSaEzDLhNaEeNfYpW0CNP0osVx
1/5AEF77aocGbEOzi6EQEVKfGCL1Ai4l79OgIYZRXtbXTDmuuCtNrDir2dBXoTnFZcHoY8kddRhw
bkPtNRl+uJbzlmF49rT2ldzTe2VrPZ9uWaWUOOYpXP8Me7Gq5u6qz/rnWKEjWqTKl8jKAdUf1A1p
bZhywyWT0IDB/JJh10hMoSfGITq8znCvzarWWKMwq81hZj7TVecV0okdU2Gr/JLOenw7qYi4D5XF
WDNL4b+GBlf429zull7eXPnorT2M2jzrPrM5ivvrT8khJeSNczEkbt+RFfIufL2oUkBbCftDoiJi
1eSSV/UgGDtlblP4P2L8Za83GkJr6hmgtDrV6E8TJ95HXsAul/myFkv9yrSNsEkGEHUzJ35zhaSq
XCycAfoNLM5zVHLz82S29G6Oxkbu3AOGzxhb86LrdRGGLUKo2EkkYEwGmwabsn/VBo6UAG+IFXI9
ziViBr3C49F/y90s4OVQmi9CBkWRTKsAFurw03Tfe92WjlufS+LPmYyCAM7hjrvns5hzWvivRpuX
a5jdLujZMdOM5aPRKhAqKyIuWGc4mFRsJO5a08bs9Q7ztcZCfJh7/aLUQisNhRMOJgTKX/EqruKN
WuB22ze7h4oD6R/35ldmIoWqBK6kknrbyrw/KyGd9C0l3t7SWIuRhjsaGUvjFLmDYZQ3DJKZOBoF
n+fdWHQ3ZWHUp6UZ2FYoMqrO5kgZP7QWQjvLXCGs0aVvw3KjkFRbZ1f23sh2BlNr3MMIF3GxRzMb
DxoBKdU2ESw6BoIisUY5Za3lxgq/2blxT3BPf8PSjwWvTBaqg3xqnbQHs7FbttkbC+8RCkuUBYaP
jiM0Sj8mvxGdJFJRoWcdyXKZFkkgsOE0p63n8NoT6dAK2UJ8UC9yGFigzrZYTR1nf27zcpPqiLJB
fj39XiFbi4gQMzNL5C3MEl/TOl3OsXOjvMSIOCMTziFE5jURsm+FFO3Y8/PdLRuI4pn/GrDTq/2l
X1Lr2WKUdAWS2stBqHmBCQTpXJqKFQh4FbH+86fK35VtYtmpVvSYmoA+YdJmbRSKm5ZT48CYGIg6
u7AKyJzfxCncZjdxd3Eew8Pz9On7+oSgbH1f2Pnh3Ep7sjXrjyrlKGTcXOG5y3Wjm1FHmPc2NehG
XRDx0hT4tyRR1YkzjYsge7JhtSTRB6F4Nkh9O+tFju91hS3cmyOHJ4ZmBHiiDnz7j43Gm96RiGR8
22SugLiyTXlsde4xOcn/PhS3iwnR4HaWF4CGB7MSmoYVJWYigSfSuu4uEZUNf3KhVWMsZEBUtflA
VJ7uBcOVEUZN/ommkhZijOcRdTopjSj2yiGuZ5TqVpQ4UMdeBqMZmCXJVEaFd6l2DzbUoOTBTOe3
i09WikLQvzqIeTkftVhaM/yfeXD5dnCzQGvPscCDozc/5XeW5XoJDafgSc7p/XxmvfMoi6Q7kdxR
p612rX/T1eNYyDY7WdRldmSm8n3N7CIsyuW0gR5lPMku8dpqNg61V7LK1gFU458REiuHCCsdY6dc
hSah2jIyIh4JeQM0sAZYjW3eD2j90Eolc17qDWQ/tGA7vMzt4yPICAMdv/6+A5clf2bSjo67osAX
705JL1ljCY6XRrg7k067Rj5ztZQvPMO2GA9f+b0PAWmLKErCXDSaKLltr/3jZjrZwx591RnhYJhj
+x96ftGlI2xWM/oQaNjnNkIoUK/GVEw1ldRJ+2unkEBjeIz+eldmxigW0kCzOXfyPrugb/U40Ptg
OGOJXB1wjG/rHLoFWFToZC4ojNWsNGO6h9AlxUuf/0RJ1VvsWzyZ3Nn6D6qeLM2X+Y7gK1RQ84dP
eHRto3Cwmx4IFuuD5iRRTT3i7MEqt5tEX4iFUToDbP1hfjxSwKUi1/uidXE04fLr0aZv9cDeQ1sE
QCOZHe5EQ4uGKvlDUeS8OJO+keRf9WD6Pe6EcS0aa8xqOdJXTySPWOyT3EwY50XdrYwsF+BiMIRi
POHhbm+apURwloJ7fgEccP1Tb8fYtcnepz4vBFTYVCcC8IizwlDk4qiFn7xeXEoTjqxEIQu8jDuN
n8SemegPDBEl/M9uvuYk164lnxTlE41nDAzCvChB0AlIpePBYd93+mSx1oE8j1Y+r7yoVgShBMP7
c6uaSZUIGNxI3G3UHnZ4FpP4CHBf4Vyg+T2Ueo4fpCRTwDG7l84Q7yuhuUZjRxdrE315NoQU13uG
EOEpP7u7Mp2G/reNMvR/vSUr1psoPqlkfa4PqqToTaLs+SxoNd6xKxM9mKf4kKM3ZXZ/f26+qACo
y4ldlIwkTTDmf0gckWkqLCeRql4zUD8g6hm958Fqfdis9ptUD4+av1GT5jiapevEyx6MfT7OmDzT
bUsY//9eNBdG1MhYMFC6JpE47WzIet0VDiwSD1KIorUOSNztCg7TQoH1QiigdADo1O46CGLn3Omy
4kW11yupOJuwb2KdDsD5tY2xkBsOsUdMfk/vinq3TLIHpn+lntUlnET8y7Q/v7HzAF4CqV1EhwoZ
U4jsufKIFS5smsSuCfsU4uYTGUbUd5CUvyX5K9FQ8iyHWiUokVwORT2bZPJVDtsAdu4Mr2EpiGbW
seT3uKyBKmTSK+Ltu63ClxfQa5reIK7ei0NBdsexmpkcvshx4EOtJkZQiO3qeeVeqHkJUV8q7BJX
UwDSPbPHyIBdhZ0M0OKut4SFyed/u39djOtflvij0Z9gMTN3Q7qfsuKfN+X6QBahFUn0JcnZ1fNS
cfdPD08rtPNpnTCUFse7hva8WtqX3YCjVQKC6GJrB6bSxObbhQWBa2vTGj2tEwoI7EvbdPnnWAqs
nkn50T97fyzVlkf0WwWTVBzTEQip0LABPo0RXgiBWaP1rwREqNFNZeUkCGADD+4gwGBn7y/X9qGz
vpUOPodoYtDrW3UOatrZc5z4bOSgrFhywrxA5rvXxjf52arXSFI44LT0Sv5mUfhzv/3iGjoYbu5R
jrqz6FmtOMOQ05b1HulSOCwbUXK8POjQ5MHvuRbBqbLl4xfY1q6+szPYfMp0UVybP4CzqoeVbnaJ
XgPDPEroTtKEx691WBBNAyDXsF/YNxqmUyCeou4jCxDdjZO+sz8KR9hsTt4mj+YebCiC3s698qJ0
5HqvpZkUw4JWvLxQEEfgdO+gcXLSw6/JjSlngfWt6c27nI6ShTeO9HuPZd5eqP4qXi4BexlrNbxu
MGvZ8WFNtc8bCFqrUZeYTDFL6X+Eia68iQoeMEsw3njvuzeHu4DZFcmnyoYtHdJPFPv0VfPHgi2N
sQymi3IJ/a4JXet8S+WPOX74ZBncF9pQ9EQu5uH5c/+U5AEVEtSaf438Qzs1JDkFNeJ//jfZmsZt
QoPdRE1SmLdFfVPepGSNEP2HItzEjO48VXC/UW82Wz5KSGpb35v7lHFOH0aA9dQ3yQS4yc2XqeGS
Hwzu+EOiP91H1kwtYApQjsHmYOVJYnjQWSYPy2TlwEOy0qSxZjVpzQLRzF0qlohGJ4u5ZcCWcOvP
Bnqg61omobroxr4xfZZdyY5Ny7zjLzkQNyJp7si6owHPSlDPx59oWfPdpMqu0aMWOLH37RnXQdxk
qUAFvSlYSureWCe6aoR3MLKHisc4xt+UbM2PBTsmd8vJIsa45f+p9mFK8+qyD81HMd4rZNaVxrX4
8KLT/GNDKSAgxQsKwwsIN7YTmfbj/phxHLBCqfp4e/WPZxM66/KncPmzvNmpY+y04olV8rwElQ7q
eBSJCtZYsLU5+h+u4ti+aPF2l4auzTaZO3yti6jSJs8oSJtaLGLQ1z4l9YIcT12CFmylQgS9JuWn
thFzgTl2kRiyETMkfaJVsTfDGG+fBH3MsCmkRTuakK+4MgRFhwyn+0iDYxAYcGpWU5YnVjxjrB9l
t3zP2GVPTEkpb2XMXkzAGEbAhJ+nX+Crf2nR6Ys2y0I3GItZvmk3WZtqSOpQdDHSwWSx5JZZOW/0
h12xZeAIDIu8S0LLdk/SQ68zzO2I0qqFoB7vkZs+Odey08316h2LW2rSfhDAgHLHkl8OZ5YZurhk
3rmqaJCM1DmvuFPkGZUfuIsvuS8W6jqTrYahVkWg9Ht3FbmwEjPl9N0hPDWROyGuGiUG/ZeTgVdB
xAuNXIWeWtmMeXPa4CqF63iYx3NIPv78sKOnLfnDhJOpl+hVUBnYpE4DcAktA9PQOADBjcToz1c2
NvUKXmIbSVJMRDwGh8jR1aAJ2l0rXpH4uVmQPo8mWKoxcdJdghpwR26RkGMG3yyS58JW/Rblbk2X
Toks+TykN7qzdS7nmiFPX7osNkYChMZTmrAiBawxIPEdaUKT3YthYyCJdlyHrHVTOVOAFkqu28u5
DaJMQEiEq+XOfFz+hEXy64TwYJ2DtXstcgV84ADcxkrO9ESSZkGUP1c2yJxBy5gGnmAMa4MQDKTR
4OCMOi64eDKo31+VM+ibPZFXQNRZYdC25MldFUwe2z/LdxNsb3Tx4p83rpxRk76K60cv8ebgQzDO
g2YgM7C+4HzOxE9joKypQo6bRn9UY3tqFZ0SljbTIkmOP7zEJjrLvQms9klv31Qvx6ql2bZ5UWk0
z2OHgXLBrNddP3Bh5xeCoMSG4lEuAfAcoVI86zityCWO3HwCRQxneGQxGhi2LIuwId2x/1wnDt6F
inwvLBZzjWkm0fw8DQeAg2ur+al/SU3swAl/eOzE+K8Ge2eb+4YXvr9fHlCa9vOl63qgKXKr+aWQ
jgqMz8CNYjjG35K0aOrLFVT/Jdw8QeOOLzS4QXHYbC9CQnYy0O9i6oSEZrLPswyjh+KoqWKhge07
5U241Mcb5w7+M1lnL08KlV47O+Qulsvu44YaF9GAsAIdCriXP+PVeYwhCwromo5isGFFw0gK3va7
gG/0W7RkejA0Qvbx7vqZ4Vywv8/nOum9ZpK0dT8ctmVLwxhRnQTFCqDf9bMYFHgzBMlePYejwnJq
QYfDFQw4pyr8NSlPslsk9kZy+KsnG+FMHr3UubEthsrg0gBwNg/glngzl1Ycj9T7VNVE3fFO4Ms5
QM4MZ26a0wjsQgQAhSSkPMZQU7oxBUfHQoXSfJCJ7Drx2u8Wgp5BKi/GLrKyfIzMADj1u0UB1mqo
5t0Xk+pnVHI154FWlkisCCx+5WxtUNmTRmTw8ZDFJ7bS5bj45Pc00LKeARy//I+nauADsCCxcoqx
U3yjth/90RwX6Oisz7wU7wJQQ+NobhMc8XZElTBkRWDz2/wWb0xwkaJ2PPCU0FNBTUjkAM8AELvV
phQxhlQ+/UG6W3QkJJBxUOyVRsHf5vYKYgEMhsUySzR5nHQh7HIV+iefA1V3HoaGh7BS+HaaJAz8
F6nJvF7uvSHIjN22YVqG6JbmyO/RKJmW+g10XunpzBtkjCRgVud1gH3cozyGHwZ3GMYy+DPVe286
W7WJJvNeVGcQw8wEHlTFn3JfXN/xOGCyoAUsYIYcOSLaVLnGnJDk3GGelIkFnzZ4Bdh58fhZ1LPn
iSc0jRZlT52FBGPP93EdP3a2aIdyb8EsSFRh1GlPY7LmdCN0+bvPfuvrc6bRI8eHLZKfmAhGJ/VP
aJaTmrS1YQaQLW2M7gdYf5Cjwy8gudF4GKM10vmkszd3cQxtihWHUe+jricfq2AP8Ukjg+GEfgS8
a0bFSI5F8aZiQHTbFCfae0P2mCtYOdFM/15LXaSMasAOv9USwEqT6AXVOVoeB92+heA+zbasyurA
dz8xxZhbow0gXmnuM9ef3AkM4pNB7f+oOlyyuMWkKFfO/SlQTBJkjsSWC4eW88IF9TJBVjY4zS2M
gjFXuJ39ZfCp9BnQLtwezmozdw2K9qxXzqcd1teex86V8rdNLUNkX0I6EoCogPReW81JLKehHNzf
8soozxa1xrGL5dd8POVEvrf837q6vt9h/tdoR7P8Y37t/hIu4KxYbQm5FS3Ac0CLeFb3+EuLBCB4
9m+u+1CBrlPYcOC0ROWs8DS6T9EohYh1h20Oz+4CUenWLNNTMg2Vl3GFTsSzLOPfxz3t8bpm5Rpb
w1T6DD3PWSdvJAWJsWNGmMyPngCWZLwpvAz3RS1jVIdmq0znR0L24OPo7l8fPtvLGoGmFw+eKsw4
4Z5nci7dnZ26QnrqZNY/BVRmGhDAJCbyGo4Xx7TJ78OTMlrK9pUozW7oQgG2RkPCgM3AmU0FiwIh
WRxo7qh8e3GMMJoi0UCrmkmA/JinN91ziVY4bDSj71ORvQXYT2gcpkjfLqZt8SGf00UZM6VQKory
k40VlPty9N1kVB0kZsubSwW1rSyM2gCCaQKYAZ6qhfi3I5GuEIn3v+RxS3vk0I2+nZnLrW7HYGo5
O35dB/HE2T6IyILa1JWB+2rtVT7BM+GUKhIvHfflte99m7Flz5l8GrI6Biw6LjiLEKslmjZhjfQQ
gXhMyNcD0fJcSTTfAUWIuyxMfwR3QEcP2fypaAY508UX8txSxY2wjj5mSr2gNcU4mcLarMB+qthy
EXD92DniE5N5cTbZhvl/qI+VYblGirQ/9TD0l1cXTJRX/K0z4bG3surHjDNIUu/qOS4W9VvVEjGB
6dwdRI+zuQMLWoJGm1/sQfEMS64Eum+klv+2X1UuZkRqr6swZnDWH6qsMLOnNzASS3HxaTsqHlml
dpprc3vJweMtGV6my7qnvFK7q+ONZ/U2Hrdqc9shTAcyiDGS7W+/bIdBp4rOKKzM+EhWzoqVPvn8
VM0VLE/BiA2UHQPGDojhuicjQ2rj1G0WJ3SHLRJed3MuGhFGZgoJJsCWEojVZSPFfFCXqvxH69kI
qgn3SltijldLH/1duaDUnUNc4qCEHqPhvHK9LA/zV2dVyyLslOMP1pYz+k2osd18gpseH0r71HXj
7sOyZ8TEtATPMbtYwPQW3AJPR2Ujwf6F6uFYYdRwkUegaI7pGtUgu4R5c5i3gvT6qUSd8Gb6Bhc8
IVgHxpELlQXr+fow6FsCRCL4KubKUx2u4Id6Ic1joTAIQkL2iKQgPlf00tj3ar08kAfXlgD9ckyI
uZPYZePtSlkJCd9xGbzqgY3g4yKTvfgNVD9GAo0UXduMGhGYnkmzDdQmBGYnVBtOxVvmF5Dko43a
6DU5mQq0B+20QrCS/FDlQePhVcTQKnth7UeCiK5CV7tTRwifdXDtimPDn/45MfPnQvRquaX5MHW4
y2zwfNvVleJ3sxsfS2G/RSo+6o5R69Q0kGXrG46fQxoSuZhdEkXjmCUj1AZ/1vIX5l8RDKZLp13W
1Yc2ioJToxIEZ/nEz9zmYLnzSmSdd8K84xhtmfcRUoG5w342HtedeysdMbfedhFvD3lf4GS0pfaG
GRwTEBFicJITcvYbfq2EVVmxsDlI1YedpPH1DXsjjB7Q5Yte7NDIaC2DYnUmzOeVXTUDgGtDKJjZ
8iUHqjB5KbLLXGD3pvJnhY3fU+FkoPm9GO9fbQdHxNpPM1Nj7K7OFn/F78zFwA5MO+FlpJdTzC3i
OpZ4M7l/tqYrtB7voA5/yIDvHAHdi9VJOiAbzBdYyKmdKQiRQ5NIgtsOgFwA6dyoiXaEkV5ddXFn
fxfyGpbdRkz8oFCWXBe5CTCIyp7Wb+JAEj0XYuB/YZwERZFtrb97F7XXb7Ta4+I/+Zas0249hxhH
8S2JqUbFt8VzZ8sFDQjI+lfMUJwTsQjE5jyAnGnfaTTrWKR+oRjnwBjNKCHLiy4UIZkkmS5rD+/q
XgT/G6tNwC4UdAyw/4GpuoxRmvpzsNfKtfbk1d8s/x3ueI/G2IwLtANJYSl3sp+QTebWxZ/iorzZ
54d57gCbEreOGfcNrNEASUs6kTRFA0JByo2+oXBdAS5DzCzi3FkHFkQ1JDhOqn5KSZ6HI4awcdHx
wpp4jDv9GupkZoIYRscQdrKFJj6Xl3m5PWHz9GPNqIyM8BonBEf7LOkhbnTK/CleUKNvv6fVLZCs
nZyH0epMv8ign4dBd5TsNyUt3z9nVujsrlSbWbRi555mypwRlWxlyuDnLkwGDfMeAXeO+/QPN2yV
L+fjyp8Cmouqm3p7WpzJVsglXvvPIon9OdmFnK2vz1m3nI/2bO96F89l3C6xvc5WD9SFMo4i4MXq
Dc8WpWPRJfMWiqSbHWJ27Xrr9lpM/cKypSJ+GrRhdvzIje/f/DQN4M2D6a9zq19NHD0e+UU/yPI9
jmN+5Ls99Li5XC80cTBwo59XAtdJri5ZAEHA5KC9JbIDEvwrduYxtUFceEBNw077/4P0WmrTDHYd
SHNcQIfnURmvywGJjKtMISRqYzHgi5x3gljQZ9s/WuHwdEK2+eRUOvrpPvA8xxeIoTZhOyvxHgUr
oAZFlp+UAMxxqn/GStCtm7FbZzAD5FhkXlYdThUakhKehtQgmFTHSCSA27tel1qqmoIrT9Szo5Qu
Fvc62RW6nmpI8QysvYePYQTx4SlUSUxxIP/FV9Lzg2VaHVK11XTNvTVwFGbF5gzIJcsuDU/IWWbI
OfLDAQ+q9Mtx8B0lNToDO66w9PgAcms1AT8yAxmIlfIKDgItXV5jlYzWrLYtwAR7y4kzeiLZ/Msh
mecGbz3tnLo7iMopVpezxm85I1xmdEapH67/S8pyDr6QouHvsfyIIzZhMtua1iNzqTXKXKpWbWYY
x0RbcjFnZCBbAuZVFb3m11MjIUzueKJlAeLXJCHDNnyf/V0tLHKpDDZOOntqBbaa+maKY7PRKyBT
nxCAuZ2I1tWXB9dqP9GuWSvwUtuxyVwlV+gIWqDf0bFIpfeW4BIhyQjp3y/p8x8MSppfEI4MUHts
o4rOzGGS3xdRHL3vxL/X4X70xh3EsLwlvUNY//sg0yQDXNoXd0O/PoKEhYanzD22FbWCUGn64wk4
wFCbtd3pFbtdOkHP8hyBjTyYPHHZOOBmxme4/d+ObkOAPQvwCb5pfNniMOEqjSbyinLxpLzx4GaC
DTbIdV40FnF0P6K9HffiK2stlWBg1saSvlyBp+rNyqHvQA9BAYszPz9LeFu83z90Lod7GoPjOyD1
WwlVpyMQEibFcwtlpgHcB+O7nYpyEDrmN5DFjPNhrDvIEmcbADszTay3QuaaREfj/x+IfKPSIsvJ
fi189e+Mnr+/ygSOTswrS2d3E4zf8JFU1XeyaFMGDXfebxPqi67mK+2grKMMFtBMDl5oEJxrFZLA
00SKMTUZ31X9Ig3EMCtuarSta7+0ZDC017DUyRSPHX6QbT8RmhjjDVtq7KJtu+qg8NSXplWBmQ6a
OeI6PDQ2cet4ODKciLt474HbSQkutSziijoVW+vm+WzyYIgL8g2JFicq9AeRckTEkecPCXd8QB2i
OXxi4SFE2oubDTnSrjrG08J1Z9CAlwfYWjr9dYDJ9gKtgdy/15KZpImIyPouMKECsqgSdjVVwY98
ZL6eabVDp/BHQIjnlz1IQeeVFcszILGF2ZgrjoixvEe5CjsguFuG1rPOXc3jlC6qpqwRaYR90RV1
cJRvYp1FmhPIeo1qVXZDolUmiW48KUUMaomDZJFCpN4pFAmc4NLyiNgXY2CrpwDDScIGBw4LRkTU
6Rf9Xm8rV+A1B7MEp7miVIZAZ6eZbgRINiOEptx+b5iquS//CVMSzsuWFAcPNOJJV4fYC++dXjne
adjYwhh29E8fA0os5E1q8Ehjd0eHLuYw7xWEXc2rWiRclGMm2dal7A9hQkVLAPNMteHbTRTbqwNH
j63RUgiOtMj1agdrW8PKq4ZZJNQdKlajoHd5B1/8qa5G1EBfVSd02DtxiK++i6La6uk1suO/zuyO
tQJUp2iMNV09nmHbe1fMER/SubuKkxR4JbSF9pz3Gmw6O/Jw5fgsCv6yMwlKQFWqEqlu/WFfR7vQ
pEOpimdbI1LXtstyMoCNRPTuSoz/npbSg9dSeeAGA6q0IHw9/QwnIMrkzfzppGirVZ8JsrvYEA+f
Y5NxIzCrPtE3CeWr2XxJZ2YsiRAkEFO+/nZZnzShq2A7tX2GB4otfH09mIRUQYL7t6cd2ExjTqDm
4xKLx903NLV85A76Et8AxjPe4Z+EUhwAxdmg11gMF6mUREuvJltdx0+9mbRm4MuVb/Uh6e1ycDry
iYF0IKHuDTsiIh1pvfwH81ccra1x84fSPcHSYYtMmZlrLaR2FgenYG41HcRSIe/2tFVbH90cch19
1lapmNQcw5UdFKRd9gpPaV0Rp7iwYdgNHoVp6VLgscu0vZYLpfcHmMSsh6feT6SvAUnavvUxQb+y
+jevUnwlT/TXlq6uVRMBoiMlFWdAg2QT7edSO6VcKLd42LO4w0eDxHT4+8IWkonjXRb8moz/ENiC
6e3mF0eTJ78N/Rzlv54EuWr2PubHZYGD7ABSrlIAjNhOf5Lfv2LOlJcnC1GWJQB5/D8q1Qy6TaXN
oSinjuz5t85XDZAXL/mH5dGnvszhAT5KPHUmSVagiGb8q3r2qlEWSV4ApDUdZ4NTdbJ1xTlAR7Lw
wlPmo38Zhswkt5oogVlKFprXMn8F8rD0NDQvPNuAiMawO1YWXQrhBHLBFesz5CT5SRIQNyIvUaVD
bdVqxG6kv/SrtEzNDcyltYYaLn/hPQ0PY+4vDjQioZ8sYK5HtEqI29rNpvMV2r8UySTRMGMogCFd
sVYi9nTIRV7K+hDqPq9klqyR+BXlEVTizpJ706pXdhYG+NAtSG8ibvN2V5D4Jef1Y3//mym0aHLh
V1HLnf6VtXQwOliidCzekkZVQq82e8LLqFHq88Xe3egUzg+NSXHp3YoRsxv75lPUToquQgWQNTCb
WeTAXn402Lg62AhSAWttVVACd1exNGXJkm3ADkNNsM6h+CaCRGnLtTffgGM+AwWilgHul2ojHEyi
46P3L4k0rZHVB5cB6ryNFECfuSOkPv812v9daSzVoLu/KllU/6rSpvnaHyofQmZ0dWCtuabTe9QG
Gl7ZYzv9WN2OmQKYXwGpCnqSzbmF1IOOVzGhseQFsAK3JLOSybn2DANOTUqwQ6RSaQAhqEGUKvOX
GQ5xK73WO19e07+Xy2XIVUOauAzfpUMIOwt8S7UMmnPKnMApp0Zg5YRcOFKti+g6Oy6ZLWSdz3Wq
5Vn0cggGpr6rs5u1Bn3jAq1+FWIhEAvwlQ2B0QS53LMwKtdh/5/1Ng31mJmqHVxu50R3ydoKCJIk
+1ZfD6QrQEgDQqleDXz3wrH48DPSqXKPsuOiNTT4I2rfqDzmHXrOfEzsCHlCbt0De7Ue3ZWMqnWH
EQ7oWcPL5zmV7XFhf38IKYkLpqp+SIe53TdKZx5XJuVnbKuXHj31vhIueD5lojjA6ZB7PXHl1kQI
v2LQPcSgRs0QnDUShnmvYyzwAqDD6F+3GcCO5p4GM43tpsv6H1lRs4CbdAT8cOkCrT39CmVGLFe8
y+C0AvGB1mc73KeCsLuWf/D6o5jNkZW1DitMCsOpgFRQ67gmlDh/i2KrDCxM3a+rYSUS4VGMpsr1
bPABbbrzJwcdmQ1wKMnd1PDC61CAkjlWIdP+8tYH00noVKxMz3bC3W3LfIcxS1YWHpOBf4bid94X
9MU8XT/dbSJax3LVrwHIXOB3mQxCv8D81D5h1RYzoh7x2zbAvcYZfrMcswEpdAXiJgqDPUWpAIi/
+GE2BtvS8HsI9h2S8ikf+cmL+3ZFWJEGgjsaiD+UGfALCCyEyntfXLwIZlr3x14ZS3szDxd1iZp3
PpECmppTSag5VYhN9TsAN/MEZe576fGNp2+2WSld9gRKrUvr115kQG5sIz5g8/zlenn2lnWV1vNH
7faH8u2G9TSmdA9f3VkHkmlrIXeHHteUNZwHwi6JRvpaEgpWG676HZuuuDZf7H+FeESyXxAkg/yr
e3vF1a5ytgrZi0B4llTpeLDH7s4stsMpXjrYCGhoO3v+s0WinTkXdu1UezaH7bZwOxCDWY/teKTZ
YZTILunKUAoln3wmOmLiB/2D/Dt06MYIHaQJqiEAH5+Nl9dPk91cATPw6WF2RJxfWnnMhQQM7trl
E3GIvrA8lOt/COxPFlrzeNMEJORAuGbsBT5k6iO6kOsHst+cs444jt/Dy681quLzXgBNF0GJfeuw
7SrC0H4/TpTDyxYUjeZ79i4kWQLIPYnKW9DI0JVDOY7lwMNheL5080hWniUCVBsgnbcikNB1WoZd
vYR/kBDqcVNaLcaXAsiBhOKcdfbJ33Uk2PVazyENqdbxC3agfWpwsocLAJmNmnCQN2Z4Nvx32Bhm
W2AzD+IPht29oXJm4PU30G8l1p1paGzQNfuKIr2d7g0p560UiqwdMifzggI7y/7SWLe2FkchZUQv
+szt7A0VUdcRZUo3ekZvAUEXNtI9zoMKEjkuYzA14+yFB4MU9BvD7zbfT+7qj9NwObiorWIDdLFm
VjMVkM02hIfgydVE0rrLHswtb484t/8f8aFOvl8928NojV561hbp7MO0g+p2Y+XVNn7Nf6b17v5H
UiPPjZk+HnuDrgR+lLsh9C+FQ3VYE21hHqzcGSZlAXaMsRVqxYCeLW8TUVprHsAW3nj4/JfjQYj5
CUY+SPGzkxZ9617KKF56dJv079L3VDSuzwTQZODUS4wcv5Trmx5E8iWKiIWmYRIcC+JX9fmw6lqn
s/btRhob9J8IPly1h6skB+llflVP6b2lTLR9ymzen3Iei4+H+Dr7hLXBSLscwxxKnvndkgjJNQML
1HjRMcPQC0Tsb4veLtQTpayL+o26Ckmgb0XhONnY6Gs0BQP3Gf+/YMvq3rblC0yfXz+Bsg5ddcQ/
gcd/JUxOX7PfH4KBrLJ5Sl63vhEOafO4qPgk7viF+ZdQTuXVXDXSHUsgWDht4QAzeiYMXrZk+JA8
dG3B9ZXat59LptLChZY8mZuL/mJlRXtBoWf7yj+Vt2KJZl1gAF37inRASgLfCsAC6pz01ffxSRRO
+dGs+ASmY/AqxRglpf8K5+YzShlMKB9c7N3nL1NEhDj4WNGitnPz0P0UkRCbZ0MAUXS32g9f5loD
MR85xIgH5JIZrM5orRwGSWEjydtZVLvSQatRrR37P7aBGTM1EwjJps/AZahs6AZiiugxac/qPw0J
gd+QqWQYPirnYrbFzGStD4pOWieKyUR5OwTKAILNJB/V3dfKs61yCzeXw22Ci1BCCQBi5EuFLbIq
pems/am7iiWp53SCS3bAwfo8pvc+3jkvoTHO7MuQVtUif7ibX5dWWbcqfoHQZMTIdnigRKBuWYOk
wHZKaXvjYG9ICg8CyotzBi/EO0kKaTDQPBHEyK2m3pBp1UAstcxAkQ/cQcNrWU+n4uryeX1MBnIh
kftl0JPOvVZZbCw+S04ydT+HxmP+FfOHrZrACNjHkQvZ/57p3/W6MqbOKvaJuFrT/u/JAdAGQDhN
dZOUjmXGEJ0ElIcoEyq6crHV8M0GB7OsmyGyLc7S7/zt4ExgKyyIxrBR+buuc4qqTBoCiKw70GrB
7D5sJIRF+EffmFhjNdLamL3t8Xv7bA3/n5Eft8akgSKlJvLYuzARd2TSQ6XYdsTJv6KslWUMe0wU
XlxEamStlqxumubjB+ggTGuUp3QkV3ecEtZnagiJFv7RCXE+vAvlDHcgxJAO9j89+azppmudVWCH
rjQKApOgeYdZXTanA0aq8mrrzTvas9VRYDGmGQtMf4R2maA+AFzV3QoXfu2qNTaBoC4fMMxS2v0K
PaWZYiVqL5q19a2ZQ4gk7OEQW7y+g6MrK6U9guuvZ2yUynEl5b8btF9h4sp3wgU4js0TSl8su3G2
qBhHaQjanYiGcNBh+FxdYhg0I92Tujvn74DfLGrCzCwbQ0g9WP6+w1iDF37mO8FbrMGA1YXmFAwJ
BNEmhQOJCzOMdf6ieVzLqqj18YcaYhU+4E6wZBA77+tP7p7wO2xBkFUCPHk1/fpf+HoctUOSNTqm
+uQF10UzHGA7y6DacfE8tU/Q5UkaBT8jmz2TdqMNCyatcF0iJhQ2TAMm4Wn9GE+FfyKT5rXsLhV+
WkMRlLtpyLEz/ctPIgNPm7rycfBpIFEkp5/Vnfeo634+M5X01KZdKg0tzPfeT6i6qN+NxrNReZAU
Rr53aphb/IcbKOjKYLhwpD2oI5LK0o28klIgjn2VC6GyeEtPHO2em1lwOH39SqSOubh7PPS8X/0A
hxLAGSdjbnm0vpKFLrRWQL6bB0IuGQ0HcamfUZzl6xM5k5WLCXuik45a0eT58oYhACwdAe40tkHA
1YHvy3u4SkeKwpocTbUqfDo7XfF8UYBQOKk+dHZa+/0W/tYGRUyVIiRZP+D7r4mLoWBAtUhmq2l7
B4Sn8slvVpXvKq1tPwiIkPBkmhsI3iUy06iAjJpv849FcBT/5PnINSiNKCVLgMuzVgz4+hwUaWTb
tEzIYQTBJmHr2TiXCL2qX69IcyjhiNXxCjlOvXLZJqDq/d91UYhmNwfaMVQhYoP9J6Eyaoifees7
P6ZXADHgOm6ZfRQMlq6oiJRrZb8z/WQ+dd0YxuaU6dYCJDz8dEQS+1XDV/Yn09CeAyPu957+1Bl4
p4DxbYaJKsbDmB4xBp2s6W3WgL3WkEjBDFwVtKs3ZN82NF7NtPg070WIknwFnBEF1a6pNkVg/fWv
Yw6FTHFYorTIoS5RcU8o3Qz4csgzmlsWS5w4OC0pB4BPInahjdlA65VAWmljmmnJW8GPGc104gSz
IwHFigzf0D7KRsRuSNqmPbifIL4Rf8Xq0KuzzWcRJ44gMNIFEuVqT00nzFDPy6cELw73X513ksMB
Ii8e5XQRG/rqcjc9JsOMucX7ttrubetgScuziDQjr6uGpszd2LcN65TCigvolO5NhlRpcI55xAJT
AFOThnKUkDYGVq48S7+8XIisDo7c9+/PAQ+G8+r6LhkLE/oCkfKk1oFjItZhsyODNxOCHAUfjVnV
sx31eQCqicGcXgopbyi5N9mQ51+WX0ujWQLZbDpaIGT+U5XQztHMkhfn1qvXD8F6R/qE0uJBcWlF
BUGvvQ4D7TWS4pqjRLgfnjW7fvkAGb5R6nFQ6iKJu12Se7dzqjufhs1HhC0nvCJAnap0Fdp4FTjb
z0R1w9pZ340hFW6FEJeh7Iyio7b4GKstz7JtZgUPtxDBn9+rTpKrCqqMhnEC0hUCDqwfaVGO1iiP
kSGXMW+MWM010y9HydQ17E0pWJyS5wjDsLfYjirA2Rj+Z+yF7paigtFNawEubQ0IQw7Yb2bND4mv
x6s63Ena26dBfoieyQ41B/hYfxb/O1Z7IWoemieIx9UuyEJtPAUqH70EFxtNY/Mq/7xY0qGLJJKp
fE+LmVEqOE8phn+fK8E6fIKd7klTogneBMfmL1uvkiSBKxo56cAW1pKwSK5Nm81Ga2ix0boPn0fc
QWWiHOiLKr98UBySxOdzeFzRWm8isBujKCx5A7BhtuxE0AIBa/ywUrVk2EqTz/FLK2aqjVG3ppf/
KqjbTMwYoKjmmdaNob3uwTKYMFbTlg/+4yrinrQlH4ZQW31fx1mNAQpyocr87nNAisxIt98dn57w
D8of86n9TfXvu/0Zb3Y9VXY6LXHA7/AuLTfBOsUv+LrR8+9IFDCaZ6HQ+Dl2D0ouHzRd4JeJHa9a
owAY0HZwkCOodSg/Ng1rAE0du4yroJ0/lV2RMfk+bXXmsB7Yt6kHV7hyQ4ocCHduFmNvUK1+RMaF
q0/6wD2a4UyZvVb6Fd1RTI0gW0h4hbPhwzvOU5/yS957sWoREFaHcSfV5p0oQIMLqUnCRz+TC828
q4Kc6qG1kC9GG9xJyCiohSh9zxS2QPbEFfFUp5SpRYlyCPKnp4qUt+/3JUsAUP8wVpWroIypf8ml
uwwY/vN55f0raKjVO14h5KlE1dDbM/91UmIFUKk/9qRhUhNQoyMefAEL34dXHVgacF7Re2Td9iEq
xcIa6nGq1oIfsKFx3hZvakeGriT0xucYVtfNa1vADdpw/ZZfaSmEDz0esfm2jABtvjfXzsD2R6yv
ywrrmmIeROVSMv1O4bEifFMNkmZw9onsS6pBxPNqqxg66qVwU8uB49DXboq0zk3LQm25zdCX4+M+
OdtW+DfEGNRABJ5XNs3k+U4qQ57UqR/jPJCtAvqc96GygLiUJRgpD4j3i7VOT2PqbDcWaJAm1AFC
B5dBwIg2bz8pKiH4/glj5fp8d09lXw08P3c5AL/8lGoZ4SqjZtEYcT2vNrb1Pt7sY0/pocIrOE2H
pCa2qN6fJ61ygtrthAywKXYEEmMkdbYyHC1Ve6bmDhKUjHYd/Bv5wBvpro69W+x2REcSGwx9N4BH
/pNXbzh8vZsi6a7J5WzFX83hslNikXdwYNW0JaE6FpgwpsmVO2NX6bqQJ5EIWjK69bWcxxKd/E1p
XKyGFby266TbXOX+BzPXlhM5+Un57IUiZFIC/HZE7XSARycX1ItLqBNkkBKLe4WRBUkzpFbeyxwI
MFhSnNvNbWtdMP6MsaZpgcJtg5yHQmW2kj7REYUplWDgvGBkM/gNUUh48fY2mMsjidAeJ/qRbKV1
pubdieG93CpqIDzyVmOVIUO0lmaVyHT+OsB0S+Ba5vF9L7pq9XIi7LYz0KJxSIpz+Kvu10yrVJJ+
ngczfYpUyggrEI6w9VJTlW1CAATxUEk3E8yNBi/4ScE062hRiNxZHdWiV6J16JoHJ5wgfRSU9bPL
tYoQvsitWRB6rGLHDqtGyxJDIMsD7tDJA+gExMYNyr3PfQQ6Foe/pP85Ox3JmQCGtx0dISpd2mFK
++w7/LoT6dj+kWzRimLxM+LOCj0hYR2izsaHH0/1RpmEuFdR4kohxcfUepD9uWMfV454CkPZswUp
w+RyLg/kWoCIERCLgu4QakBq0+euCi3Cit5Vd4j0ti4vf1iRTKbaS0yyRuClEsGjc5IrBgbW1UZa
0oDHFlOj6KmjTDaNU6ONs3EXqV5RqMCUSFJuLgHb/gjfKtKw2AVp8/ZgrEuIME+YxdVWluapjZXT
1eVc1c+j5l++wyUui5HkjuaTTdYsyJoKPypRGEgEkJisCxHr5xP7JHu/K0cJNktybxETnmevj8Vv
vIDpBDv5oV8OaYf2b4dQtCNDmxukhH6qP4o/P27x/lQSVQ3VGrzIoaGq4uJRHb6TU1loiGPitiZE
mler30EPYSeHQCjrRdBXBYeDzJksTnmkOTSjzrJZYSPXVdujwerx1BC9eRwTvzwonjp0SZtZjdWp
84ai3l0Zinq4MCdWwy0xCX8AyRkNTwyIqZnB1zqSJdbDRn1rg6dDVoKpVkuV/fmUHk2hiISWOOiI
Rloi0Hz2NC9BZ8wTTTELlCIF/xEAr0a9S0chKCkUepyAeRtiz1gV0JJqG3czmdUhS2rpWiVfN26+
Kg78SzW/MHsoGC+25r1k2uSAuKqE1n7eWBIxf+LBKs0zhX2n8Mpnp5q3anZ6q/LzJa9ItbKKNgii
FROtmwE+hu0Yl0dhU3seSgL6B/i9Dfoa7potyS+GfubtzIn8m12TUk0etd5VzrQmSsAHNYnRQKhO
omsIQ19MWL8S/W/MdjRP1qveVounU6tyLV/OK5wewLfHbvu53iIvfbSk/HIktnA+7ef/5F7zJiYa
hMMeT4Dt8WsU59X/zpVmj7gHbWzTDt5UWZ+Nz7M+tmhRyvwA64COunCOH0U/9KG0fRxCiNefbb0L
v3HXAjtTSZ/spaH6tww9w/0PlhMqTT9hUMQRRfnSWvExWolH+epyycy0StDQXx8PnMXPflDVshkx
NtcsDFh5Q8adWo+OaAbuR+j41H4jPk5yjxIXRm8gkKbWi7vn93j6HOFu8qMipzWAJENDovcNDbLz
Gl9FTz4aocyI1doNhn87DBtyhRDBv3uAgDsLPfLwoJ9Vl7jBL3oYrYgonyMIppnhKNJZdWOW5Vox
04VwgGKsmWl7cb3P3n2s+GcLVPl1qdseAOcbULGgKslwKIHuTuxtkgF6xwx4ZZyi6PknneahOeda
Yo/rtO825iJtwGFDAFFC3AqIkyGWgHcpQsOE9/QnT9/T9vThU+nH6yL9YS4hLiddjBomfPLiEf8w
2O5HRHXu98HwhQWVPTjXpdbMeiTWJZhO+jPICb6qc7V2nOQyKOdynBOXdVrJW3WB9u88UKhqFRKt
uB5BWkFz90Edkj6Hfj+9Hs2HNBQeYJf6cH4sO27H4NPyaG2GIxSxFY+kDRqZAIPjbjmDOV45FRI9
PKVAKRdNBdLfkqpGvB9lb1iVc7uUZRUuCoEipnGkVM9GJiFoPsOzdtVVe7FbfNYHToImEk48lRGq
P8OT90WCZqYqm56OcXDyoazw+6q6ChnFhtlWEUxAwoo56MWN/Bc6JqwQdMfjtMrp99GGtwXBo+9b
GjrmIsCcwc8NGHS80WPLOVPl+L44q5UVlqF5V2+xCBsfFiGyWhCzaGQ+e6gchaNgyUQkr3jyittP
FOjuBr/UaOzNlOj3f4ep73hoKHVM88/1/l5+ff0E+QtMEOzjA5O3/IZD/QbyiEM5Qrhydu3PLCd6
dleGr4DzpFF+I2LF36emDCFGAb09H+dwt1Jg4dxG5yNLZ9IlHsnMP/DQR7kr19HH6Tx9vxB77rJd
l4daRwZHvH8kumN5VRRYVeiarRNYAsFno4lJnCr4u+7n3TDhn9nwp1U059u5XXpTh/pjgJCM5FLk
zikcNsOqSM1phXFbXewbzzPWizvAnK2IUOuvi2m6kuAVKAUYdOVgRPsdiyjQGy6zHwOQqA5LoDqd
HV7brJGbrofwjlM+pDf+pLyEhhrkuTmb/tb7kySnFmTMDL+DpvhWmlhNa94uDOYZFJguKJ5un3zz
CdZgJpu+hzRNuDP0tMBZCn8fCmx5hBzcfYuEayoaVw2MSmh5MCkMy8COadyB86Q1jmj2Nfjr6kEK
N+4muzZ286XTEGfAUiff6OXAZTW0W8u5lq4TWOY8xMkjm1+6e4Co+R5Sa4uOB/jRJt/Kr/55XQB8
bEiCXDwK7WkduSdx1EzKLDiBBWHy+K9ulM5BGwx/p184jKGbubPmWYjOVvgqZEme7qVas0TCf0im
ay9Wx433BXMV5ZputPOEqqA1amOnCVXVCVTe00IwiCFDuo+GMuS6x16A9D7hS6ZyyYCM1MhpInGN
nWawyQnfe8mZ4qUZ0dDVS3o0Bc6QCCiO4Nf3DJiUHL1mypyhliH4SqKtVm1JIKTWBLDse8L8982k
5XawWezZyW8mqunm8B3tDy0a2MNI7Ssr2GqbBrSlE6hAwHXnt4sT7PkeryXdOT053FPseplhmtqF
MmFV88+ubi8abzlCFwxSw3LrqG3sCzWtD3//QntaX2uGeYATTNfa/SmODmsWRDl7Ll0MYvkZsZ3o
bjUzpSbIPOrVqsDtkE2cloqJVikxR1YbTvVjoxzeD0Ahq4UqkC14khQlQyoW4Au6HB2vfPULkOp8
6DEqE/XUa1sZcV6s/BJWB0G/gYefraIzLVPDmuz6lfp9ByABd/j/8TJ5UWL+98zS375uTVXVrxiH
RkteX7VTEYhZ5p8Zup8H9JrGOZ2RvwHSOtRidV5h/JZAPAhObKHgHEEJ0mvpdgVBKtpY6bfmeW7M
wALzUHBqBgQb6hMIUSH3PhH8DzrBurTHUlbLRNe7zidKnlJXGut5kebZmSWfFff5wkal4/tGNV6l
kOEXCaZFz2BT+EEaB3wD0UCMPa6sNttNjn7naEDpxaDsiKXueQ0FVP/9RmZpvXZGAm6S3kI9oTi6
WFMY7CnbzA11frSUBv7NKlX9i9zLT+heCpshbvWPeoAXYbwK/itV26HS7MZeHBaysoIzh5rHUooV
RTmDNBSRD5kDhFY1h6QBKGpbaHtJRgjt0jPUHlvLOaTRP0l516wFLdQLniJQ5EmFUZ7Cz4efP2TL
mfXG0vSOGzCfhlEbXiz0ceA8AAu+rNgF0DObXOkfpSEW0nzz/Jz5KyTVRaQx1sC4abEtZFA5pmKO
SAOMb1QNn7SvD6SZB35v8QZJe8iOsKroCLeJl50YKcxsNhyQnx+qK/AHKySAdn1IeSiCk5Dv32oM
Dq1uxMggfJbr/LHdWZ+SllEQVyhnkFV/uQEdg4pCBurC+y1R3M6pstCsGvNyZ4pdW2LdmXiLaptr
2a3YEwohK2/Bf3cJx+dQBH3p5JFapVm8pWUpnfoJMAHYUjP7OOd+K1Fx3dRmxZInp5A8fVjJL04W
kAwjkAt4Scl/3xx45AECqXbnv1Q9YBVSmB9Iw1EqVqSM2DYuQ/MGixWff0R3itPXJbRcfszjtJst
+IruXPC1m99wEQvBUBomVeeOdJj4Nyf68zRyWt4gQsfI6AfduUXwn335yOhl1WnKbYQyBpVSTAhM
06DHvLPE2ZmHZj3451xwcpbF/W34wfuKVCKCHbczswJrmKufzkT5qgSN3vMH1ObuzX0GD0et1eTE
VZUo7b+Nc//cSlDcmJbjFdDN0ZWx5d8ir1WzalnuMlTNdU+O/wzVQg+kL5soubqg4uSSJKfuzlgD
MVKUNUa5vO9ARYqkgLHKeTMao8sj6Q7hf6RutFrSbnzjRj0ORpmpcda++rqbx+s7YJRAOyn8CD9o
Q1lbaIltOczHwNXGtdIOcmzR12wUGSr+BK0+/56oR2nnYJxsSrnIwv3UJ6nTPJxE1+ZTDThLEKzm
NvKNJWUgiSyOOc10uCPqkEuQ1GxhZ1zGSyXBltEv/w1wiCTycxHUm1TsSBd4EwX7uuL5A9lDOmi2
exEvZebEP4zUB6xwBzLZ/Ez9mIFyAWYaVr4NAeeBN6B81hdQish/26Q6sXJ1GfaNSEp9NIEwzc6d
5l7bNHD6Zwxt9UxAn0Mn9o4SOJ9Hy0V+fczQGiNlWgzcdcKp2qfPLH2mXWb6qcH+jYAZjz0OB2/n
wUWDaineRUqM2EWTJ17dIEjN7o2hq2EAn5+YpNOyXzM1QvQrJwzpWwzHuIn4nUo9qfPw5CHU/eny
jzNbkDPvZ18HKmw48gvxpcq8EW/EnhpESALvez+AXcy9qXr8Vmz/iG+2AvCl3uuZbf6jghCmljaN
vMzlDXyzXjhqmcIwR/BkWslzOanJpNNje1eNa/pkXdzspD/5a2IZUYyybqmEGX5yNM8vvp9Tqq/q
xBlTvopQs0uNbG/2p/w+rpNYpU4W+QKuOqdNxUGZpUMloRmoPVR2m/u4Rzbjqcn4pzOnF9YWYNaK
vfYjJjr5Sm0X8Y5E6pW11gC9gPl9+ofzVZoXRU/jSD/49ufaRWAf6jO0UBmoVUDhZm6PcZ9vqGnv
N0dJfcXB06sdrD7PRV/0JKOzT2Dzt35gNHy6WFH/lnC5cQWyUapubLjeTPMGzEK+wEWe1tY1reer
2+dLBEc6VW9i1EWfcYx/jbtfSJmASTzKxAitiYLM1fWUkTgqP3z99WGNm+21evrww1D7QXV6ZJdI
idd7gl4ozvxb8oOr0GhfCua4IoT5Imn10WwSq6V/9ueQaIPb6WeNBnMwIqBmaa7/JUcziZReGZJa
kcuBexRYEg+K+/6zbJuvgoz6HegnKUO48Iy6W8cTomvAWAye7IfH7OWsHQ0shNfm5FuQJ2Nbp6A0
zhftpWjJYzeoTEwZcOCc8mN3pPlWsDo0hfXKqENO3uR0NGa48p/3QnV+9VPxQKR63wcDBArW3VSy
/md9dVNUYi2R3SVUJn+4f19ZcJEjeinm4nwhO1XKngDarFSuN5eEOhVgzjKmoNzVJ4eX+jQxx3Yz
gcHEWNdn4TKzu44ngh8cozBji5AKK0uDwYO6FISYJoDF3H1kHOauwFIQT+sRbDKBwb5BBosmQdrM
9Am1qxYq6/n18qQJjso4ZOSqITqrT4tNZxx+lQozDqnv1/ed4k0/DGptcItK3zvPCHRmbsN/TuJ8
T/c0xMMTyV20Yj4PHw6k6v97fR0JYK0M+PPMVdTcH2DWMDWe8wiz2Ul2ayDoQjfyUtQS2Ga8VR81
seHw+sCilXkwLjNG00PPTWquAJ19+Sduytcdglp+d6C23kT5sVsAcm8M8ph3I0EPkpRzm3qSlfyL
F3LL0G896uO7QgK80f+FEvKf6PjQGnAM9f7BZNoiYD/Ckd54V5iMLm4w+niVoZwWEcLYUoVX9XY3
cRDaCkzcFMALZJ6F8JQzk4gWBVL2Fl19+679XWx0CbEAmsRpus91bG1rOJvaBGagUoDaYJ2sLXyQ
UwlvjNQCEPUnvyI6KnPpID+lt/AZ7+pRn48IxVA0WyU3CbaxE+jeECRvRCJeWiG0zoxYjTOpEdXW
VxuiTAll6Mi227Y6nzEtDLOysVtp92iwwOgLQ7T4FSxC9OHC336ssjikt5sAoj4hPSCZUghCrvRe
pjeiyoD/dxgpKpe3FtRTf7Oq82+2UE0dSfyzF4Rp7J+1/sL95IosbJjQITtggp2glzLZdxCoVgxa
BCkNKlSiJPr5j4295470wWXg0pgo5kdOxu9vVZPexIvc+rjSp1tIrHAoDyAmXrGmng3P6RYgDV80
d1vby1XJ2Zhh2tBBeunwNOsaYVKgfASqYfluPwifJlvAsOcQG43kuGTlgISB2CGI6rg3AE8FxHUJ
+ICTKJZ2dAUyEnS+MjlJbFKgBI62Xx35te4tiEWX1OEQ7fVJ1GYJrcbIIjTAdnlXBKTXcghcLFMh
m8u+21SD9hQfBN0ocnp/jgHwKRAcbcGs5LNXYgUCXQwSS6hjy8f20WpWNUD2JBR+kckjUUYimQmD
S41o1wPJJxjDlAqQ3sxeJyQp/F6sFovo4qERJD4TuGIhMjEVAKy++FVotoRKz+eCicZynabOYh0g
OIFnu+ZmbV5j3DblvlBTynv0oVnFHgS9Rm7E7yfjGqHPJL94kNhCalcRmKRC9XAxMFP3fz7aRnRt
mIshujrGwufGManNzoFMSYwGnkkBZIf4Zp3nY3wYUAlow0pxvARVWxvXdX3uB6Mhgrz6KfmHmrWc
8Vi5VFIVAoZF4rmW6p2HSphYyzDhlQ7J27DNrtmDCWZHtBeIpiHKeHJfgKbDw1dZpE1JKG63rbTl
kShLa1qiXujGfpdNblKM9rIO/PNprrSTFE+/W5CiYOK1ssb/GyYdFs2KfN6UV4e63iYJCSR8Dzwy
9lt+EufJa8EbquD2FnINc+KXhTwGRkDXxrRrd77d/a29UH7/UlVBDNNxLpTOWViaEba+ONCIQaHe
L3Y06Myk+PtV1hy/foijyTaksgr50aZkM9MX6c688qdtAC03ZW7n+BT4Z6eWDq72YaFg48IkyaFu
92lt/KTYu0mw0HJRbmOvPOkcQzowdLkDaFARgt2Ny2N+aZHh7l7W8TR5MSIPZwHY8kBQxXOqKRyA
JU5mZO7bskKKl6qAbvVhsDzV6nlCsZDeUHXYvPmzbn8YpwNGh3+HJ/LyB4RJf1ao5c/J2PRYd6dp
nY6TTBA+g5g5110m/b7PX6IWcBjFvaEpOPMjhigNWKZlAhEszq+8XdFi90+/g6UN0qyMHFIpx/FO
APeH9aXjfP+n/lSPFB+o8dtJnYBS9n+bKX+uVZLHnWUSE4xODXgL3u5OrnjQTT8ZDu+FK0eU556H
p4C9i7nU2fdcyRTrpD94JmURN1jPh3pYcM26O1Mig44+OIt/Yp2D3DVceA6oKD51WqK6B66L4fZ/
BdcA4OiH730KBM1M+wUbM4lAYix4lPRnnDw06OnJSH01XppKFyh7495+ZhmIhkHF+4qUv3OlReYm
CqiKqGff29+NFQfS80RoM/LQ3gWwu0oBtYafUMc6IQRrHs0JCa8aRtYXGwe10Vpqj8xMJFA+ip2R
AFv7TWKaJAqH/mToGRjmtfkbb7YIZ3KoFP+TQeMKFiXDo9JyT/OwALcU8Dgj4eFbUSzMC+lggibF
h+47t/YSeAx4dfcSs0UUz6KNxCtpHZxzCitCXQIYp7HgxPX4VPJJdMltpQcJu7m3HRLcxpLmcky3
Jhv8rLsxGG2DxEF/DRJDq47fvf0UA3rfqM6hfPbHIri9LR3R+8ypFjNAv/6MVkxbur5SdTvVEgRZ
BRPvtTIEhCJVDz4BlxN/UslDLOz0aD76Khn5OsiLm0+B3nJX9dqfxrCEzlNgKW0WmhUFX77oRQv+
wzVRAd06bK/DjrgxLTXwiBh+kXRa4kulIDEkxGy2608cj/maANffDq0yD/O6GsveFwL/DT/3NhJ+
ARLTZi0vFNUtBWvdyqrLzc9uprINBSIVHNfCE4GE1A1N59UuHFZDS5tpkjqdWhNLeAMuqaJcBNGu
HHFFNQtTK6uyI0Vh6daYTWuih9/i1cYctP404qIYFYz9J/DshaPhsBoLURUMvVNiQsg1lwUDy5fh
lww1hgwU18si7j6dd8F0U2sq/JVTf+GdNH9FvzVt+Fe8k/0noExvpRpU4/SQHue9jQoZnVgRUxpt
ygFS064Hge4k7QKbKGmyMUGDGIuh10TMfaMo5PUPsacHQ9WeN1/GcLsHN7cU4xuffFVABKCUycgZ
swvVdBOsHCdSmAAVKE/ZA7b4BrUzAtrzIsNaro02UulsplQzdnN9XOd8loMv6Mcheu2dNWvicM0o
fxoMAwdhcw/nRkQQWA7paZCte/SOcYlqGuNZ1PqT2G1Zim1r5erT9lKbRH6YxwsV9tSXoF8xKDLN
LlfmvjqA/I0daS9KgrbfvXeBmBkE5yxz3lt91GwGpkuTwMx1aravOqF3s8C9cxaS5tqcM08Q4x7h
jsXyKjuT63A74IojtIlffq97GPKO59mkHSsYOl2c0+5jc5aUvVzdK8bS/CeicrYy0GHnDteUjnBm
qgeEFA0zCOiXse0PCXH4OBcp28UpWQC0hAmi0/ObzAu1QL0W/7qXC548CnCrO15yt+Yk82QGQvf5
GvB22uG23ybo/TFX4C1qrzMFAV+o5JSKSMO3TM/EiLHdD5T+nlKt+0gkAGnLWaHXzldF5m/tXIaP
dhywU4qGhZ5bsh5i1OP8VEJ2q6+B7rDjyNviyHnp1PP63ucVRqIhyDcyOnZkOddkpTK3+1ze1sR7
G1dHegrfkFX5Ql3QJHPvFEqluStpNhorcp8M0RUeJWcrD4lp2EK3KUp/Xy/pbJa3a1WupYycywft
AwuVtNsPhaCshlx83PBWes0/81pqtMkFAPzis1O1KjxKJPqojor3Na4+S5zVvu+GpGxiXpAkW8uK
H4DrbUeh5d3FcRXds3MbJT9hobP4U6WlhFny0wZ3CJyZZwCZKiscsZpzpWbiqDqVg6Nhi25fnq8J
P/EDNlKFPsKLnlTzAJCbKwO1ZATG8S8fI8tsbh8DRtG8lDC4rcuYJMABC7doE/Fsj+bZHTWV/6ii
y4lMKo1KEuFTnRd3lYOrIW3pa2nJtFaQ35Lcg0iD+7ENVRdshbk2mMq4fPl5pk5Jlxr6obLjXbKB
kYMDyaOi2T4wD8vjyDA8RfnkRyre252jAlu8dndqwQR7Dwi4w15nJgZZu+/uBsUiNuO2FzkdWdFr
GCe2HBRIgEOatbk7zgE8AMC0AnqlUn7HY63/ULfvNlWmQcnhecwbbF3XfuBBNeEuXw7Ts2RmmKK5
diVED4/wR3UjIyPoUvwVd6f8UCpjGtRT9802xEFL+/Sg45jEPt04QIZgWXkVI/s1oC5ajhejR7k3
Tnhp4Mzmv1gqlzxbKQS0mdNGq+fCq9mH7+O/kQhcVgAgnugrugLhYb3FyTrvlMD90BVmo8auK7WO
XdjItsSDwln2t8xG4sk3nMXyxg+wyFsagcEAAUsT18QprXSnKzKflUi/aDw/rbdG/hoidvASVlVg
TkVTsQZnxip9d94IA/Wwoiyc0uHD8BE6PIaUdJd8Ok1QSuBV5N2sI3MrVlFLVwfZxC196AZbfAdR
+DyOwzupzO16JN/TAFYeQK2JrA2UZnCi9pOGOEL1QiGAtSF1+os+0p7nSeNyr+E65cuJpob/WWLX
fS1hSzl77x1wFTQRbdjckbCiCWg7gtiKBo9a7bV8Fbh4++zqPt3TdWnOf+Cf0SlPYE00Mq8eLwmR
qBf6rnanDzV2NKxbBc+WrnPd/WmCJeaZKimWEBL5QY8REfCYgt6LDC8Zd9voT8BI0zuabo93F6n9
7RMPrA6agjv5DVMyEqTvwL0Ezch6QQBfSuXIJws4dsWVNKVACglSj5xIRfbV8QV2IGBrhhzeB+88
mOgud6//05TdFT4HverHxwQr0QbauOQH2qPjMBTmVvAOwJH1lvMfMnz6cqLuuFPYqCMmQ2Re3gUN
cgFtZs9tZ8fwTyiRaok1ex3rx11awNzVCZqZVKVXKRy2rz05laY5XCXjQQHDS+OPurmNqU+Vne3k
68lFKga8vptU4Lj4mbSY7mg/xZ/8zfm5o5sdOGY9v6rTYII1WjMatvHcJMEdbzdaZ+8pkjzPSxRf
H8Vgs01iJGmEFaBAyyc0tw98iFq+ZyiQ24u4QX+Fs5o3kolosTzZ9LzjdHRzhYw3J6q8BXtEsKi+
jxlWK4Zm6WXAIdwOTTWbDVYbLrDRPJvX6MR5Xi+2jlneNT/4570crJrFmBq+ismKR0nt5TdckqkC
+Zw15wieJgiuhMsYUIXI+PB4CpyHpyWYlM3GN+BQoL4WhCLozarosnl/nlBlHtRPlH9Oci2CIeIw
OAaPURQgmqtPw/GSlT1S3R/uLJxMl8s12ROOadQUVGP7XuSY/ajPuywl/bc2Hp2oajvA/QPATDPZ
5CjecW2R38agmS7wpWHHYjpQUJl/nATU+7UQyghAQukeaHyCIlK1NTtRbMLov6uBHWrYigxP90X7
KcUwGyAJmRNLF8aXbP5CY3iPVNy6saPPMP8SDFr/m7yI8Fmi52uRwVjC7Rn7YUjPJc+og0E4oQKB
7uadvBg/911yiOLI7FjiscZQpZHyxc2wzBkqkBbTah98wMPCQhNzj0lI9nu5k6txwWqxVlsfxfBR
w8IhsYKSpB5/o6FJlJOEFxTeraIeOWfs1+XeqBm/2dXxPLUddTJ1bXdbNu8WMIS1qd1aQx+DBFTJ
eucfy7moTkuoKgqhA+z6hoKOtiRsg/ckojvaR2MthyNYcmPrl983bMXUcFUbYoPiFc7GhgpuJ7zA
esYEgwiTTBxdAlHbk9giv7yu9YQyWZ/OpzqOqmjQCdHL9aVpy2FBirpWskL8VBsxymhRz7VX3Z5e
puCgzhe7GZ8et/JC/9VLjjm26ImkETPBZ5nom0y5+7BHBNdSc4IMmfHWWC0cRRBTTQlLQbP9uKMA
UzrMKcUvyToDVcFyCLO7RmCj6hHA9wXDK3NHvnNMZwHk+UuYbe7FnDXMjB/SCOahDmHdjr+8g6/b
G1Ro82P89mXZDcDoov1q53OShahPVqTPiBn9UIp7YPnPR9LEq6wFLc63nYI+Krb9FVL9hlmFEOnH
+YLHViqAKHPEoWam1s33qxOcL3rlrB6UmuVxQ92axZ9wHMBhjnetnRM0oAVxCfM2MxJqXZzpW0tT
Gp5Z9xdidTISkDA/LQuhhojtfq7biC/k+Y+NlWdIUUX5Iqymes69JlTDRhU55SNv/c5muuSJsAlV
PkwBHINP5e+3kzA1fBgsMk0r7Q24IyELvKrX+CDDaOzBUUdanHDpv4k4D1Yx+VqpHcBtO9x2nRiG
r89BUX0/feurYdwAfUvxQHtVGpgey67Cz0twKZSI5M3dK2UxamvsRoWw0KLorNCWB5UN7dn1cGiE
aJiRRJpoz1rApGezmpVBtnyQIu9I5KeeLCIyFmQjYST608z4is3lsJi3WtJdbJmUK/YNTfHGnEZp
mWl4NTaAHvQ/WMXXkKfZnZiOZcP5Wo5h51JO5vihVRoenthBwBUPtfR+hgMft/LFb3cBEfcvFnDN
unN2EHRv9X0lTD3wp6zfCbBvoNSeyQTk8WOhK28i0dZQWye6DaFCmqzKYB86BP2Vws0hmUipfW5k
25dwoNAiP6asqclHgIpiyzG7k/tLtWUtSe6v73TajcJFjiD/25oo/iBGxhivukPcet3ECpixHkAf
C39LfyLBWF2QIBFeqY06VJkbp/an2gFumeizLWBEOJWH173TyqrCWKA8TrCwnAOSB2aYY9VopTRt
KExuBWpkYcODp5cXpbnvyw0dc2CRrLZ+YiboXdAsWfKSEMU9GV1Zy7a8jFwXAh31oDNdF9Dgi3aF
2Ed6B2QdLtRKhTdX7i0pr0dGrbj3v8bXN9UfitCxy9gLwi31Jg+2/3nUGGa6Iwz2j9yaHBx7nUTk
PNPT7Pnkwy2tWtIjy12UIYUw/UhA4gn+d2v4T+zh68OQ7k1ps8mRmxeNoS85Eb7UHN5777dDW6Um
TGssdhAzF9OFakmBldWXeXpnBKcADkY5mA2S9sSFSFzVnkfAW8GvhfGxC6jqcVpup7xIeQa9JygP
4M6FMRc6IXZ4ZDzx1eat3IwkIpg/dCX80cQNcT4aQ0rJmGYDSqVtDX6EnbvHuxQFDLFbxtQP4ulG
GfJWMCWTIW+0cNiCXOvsT0F6zjgA/nmhSa/4xpoUq1P6YZVLRncsKECdVJTqRXPzqcDRF6/rGhlt
fFQnPAESrnzqW0d157WAFfQrlliJIpkorb9Sfuh0r14uAIsKZqbTumT5DvyVmuyP3UuKryIamRYh
41AEHM2R/Lq56bpM9VYFNEsb4B1RuV9GRdRs83AYAgJ+J+oK3WygmHRsHSNYnDv4DysowBZImP6j
1cRCKMJ6Vhy3CkP/hsVhx6kWzXm+ekXyy3jEB7AV7inPssCxzgs4Ua3S/obj+5QiwrNSgRDVjzII
moF0kPdEn3kXNQWa1VIzGAPE6eWViKDDA3VoRdZlJTx/sJLNY4gJXDEfxWH6zS9wR8BNtacvq7R9
yvZgpDop1YqVIE2mLL0pJ1o40NyoZkNc803zYkvV9/SdD6VJ/+T+fM08bm17rIWE8eX7ifFtO98B
9mRkFIQd3JqoTA5jaBmUyKrsExY8xBGvy+MkCmcsKacheITC52e2tUcEdyDVWdpUXK9/SIhojl5e
wyc9Tm5jWzSZmTb3BhMjZGiwEzLCfucC6sI8N2EtF8yk3C56Fv6JHOc7ZxwIDpWVqZEv1MRIPRla
FZ4UGGxOJ/3VZ4Fx/y71iZ1nSSFOehFRMwySmhtvCqYCgiSvihfQguWTcYK+zIlHjN6bh+JCS/tS
TPnnCAxsMEaYZUuAqVhTMIuFNZUD2DGK8eR421bTnEBWk3OiAqyjTQ/GjbaweD+izjtlI5rqrIFl
+CkTSVb0OxVpJzJsQh0UufvSyz57TJTipq2tEG29WxmFlqb1ImBocWwzK0rtWZ6OB19oWcWRwUqI
0V7fPJ0vbw54Mekp1PDV9AI5MtsBaR/sNyZAQTKQ/ZM81gDQTKDUnYstxib/dvIjPJ7FMA886l7o
QszQQa4GE5nkK5GctrOgdoGsIFpjl0e4mGaIdWhzN6QLQs+Qc29TZLfRwEj/oZ/FA0m/STR8APjP
ohowhLb9C0+e4hpwdbsj+dzzWsYrtNzUcG9iNr83BZGpL5ftV+ZrDv6XFgdZc9QjZc8UkVI+E1xZ
lFAY/K2tsfu7SOJRotuHJtoQ2prIVVSmur7+qNhVsDaj0JYo52oRss75FHOOiAdXUHnGt+xysDO6
pz3tFNV/bOKgqqmpXusHABu0zleZZspr7dzsA3s4Z3P/9xiGwJWqZV8Cznd09q0INM963d+281VJ
PqXJwhcGDAx0OkXVBFv4L071laBgF1OaecXUeHVSTmb5DLB3oplLrY1uId+JyuFUEj+cenbF0CpF
ER9VaPbK/pbWLnNrGPQqFVYjWVbhF1RfkH/2fC/ZMRbZVGQWQsiIkWQ2R8llbfLRyxMN+pPQwLzm
2GSuBXvZEk2ckdoLuP9rVlknMhmg93E3HqfC90IwFidFF1oMo0FeddHAcNg+2XApNwMBT56ApYXb
GUoG0vxR/wnR7BKxrx7nyCvXozR5KGTFgo1xZhiHmvz24Swa+pRoaJSxN0Lp16eXpOsZ9pzO88ad
pE34wsh3BgQ/pJ8PBV7mPmh5jEJ8xunGXEY8/Q3s55Zf/bG24F7W4BjSz0FFWCIYHGWVtnQMO5D5
7XaxZzUFfGObP4r2kEvyk4z5VML+NJVNnY4ZP+r5BjYtwWFTTjWnad21gXYv0VgKHc1EkSw/TrfW
AeIhu/ux1GIVJ6BIpkbgqnQnlh5c985yxLdnCP4Q6QuObFM94rIzb4ijGbAc/loJoNEPGvtOkdHK
NNFuMjkh2uMQtT9+dYiG7ols+3nf7hgYZv2Je60HrU/5klLRAlxLGsSS47mKSprWb1IKuon6TN5z
VVsoE51yjkqo7u/J94z1BhmTs1URnU9spuFcf9cTDJuakXatBFaJSstuitUUjYg94e6O9vVh8y5L
TP9+GrOWafk1eMWcQ7hZFIUW/emZSOYktG8AJTwLIR9w+vkpEnLi4tgq0hviLYkGRDSoMOXLUXhe
QUQTjBS1FHLzhi7Vmd69Y49z2IgJfkJMsTZgQ8JyThpTdcmzP+9UW74hb3W9foLScYT7vXZ20OX5
TDz9CXANLulWq9Ee1IcukmvbzOYr1/e3nMQgdFyspTqIfpGbJeSYBjiC2uYNnGhV2AzKwerTiHa/
r4w+eiDZoRJobskHalUmxR0xugdLpBQ4xVTmdPGiqi1xvz9KHIu+Yk15jfgFGBdbc5X4/Rr1uUsr
uZEX7NStq7qOnw45EHa6I6OJD9CnrF76TgPY5CBLcrJeXd/t4rc+wC2X7UaaJ60TjR85zX33sB4j
NRvIjaL8PJVUS4aNhur4grwUXCWw5yYaALq1FbJyfo1OXrnIwr3ooueR8/+2F7pjRrgYfdg91he5
RkhWbfb2Lwl3qEpyXl6H484usov/RUFVxnAdsCkHgVf1g3WG4NVToWBYCtJ7bjORRRuI8/v1+DNX
OYkWRphRfgaxmYLacC2T7r3M+hLdH6LqZG/SdXFvP3jkMQY7GdVuUjsyz29Ioc6dVtXQf8xA6M1d
CT0CwwDRw+jtdIzKhRINzKsyS8xbL5iGLKq3zR/5Fvxc7h08lRhRBNicY7NXD0/dpUXDui41X8UO
m0up9x4MtZlW/oHThofLn1GGrIAUgCk4Ug92hqJn4xMpnvPEk/1/JycKkrfO6BbQitg4DDjdz2nx
mhLFdUrlsejr3oCxYBN5A9M7JHqJnB0EXi1FUuGITotPvpN641IolfKUCAJjcZURPuCQj0bnNgx7
quDLl1T6grP5X/ZSQ3UzUu7OIDnJj2eSl2HcBrINr6s460mEeD/qQee3ueMEnxgIOZnlLO35Fsin
dqs6ZG+yKuuIfma8T34QPUrBIV8UumbLCSBGscUNp+ZbqR2PjjPhE5Zjijt0MEzqgywVsHm1PqRl
S7qhwQB+AjJqJDIU9AFmSIcxSDVlg1L9apVHJ/xZV61WaKQL+UD8qtS8xHzGBC94idQ/ZjrvQ0LN
I+n7E9WhS26CcrA0SX9v96fAh4fi0TyifBW2GwbG4c/ujcHQ7XgNDGygzNeNipaw3H8hU89vXvee
1eHHj14PiYTQQ/jYjak1wGquVw7z5ouUDoIIVCXjhKUGVVFhQ+2CHlsMXxJQfAfTSixDpztmqHTe
1LYJS8hmdoO4JT9ydwDhkUZXx4h4dqg2NLIfja/UMflxFHxVyhxz2kZCHptL/KtipGuui/KpDvQM
FaBnma4sHmrf1DeWMGJ+SDmHEjGsL2AsNwF+q99w/NAm+S6epoimrsDQckFw0NRBWtObYFpDSNJm
tGuIy/bMxu9ZLpEc379XLjaFeRq3YDR+ZgrhxunLunvtsUt0/qVc9G0Qvnq4h33FNXhAqrH8TUVs
5JMGmQCRcgWYTdZSArPmq7Zez4BML4zSurPro38ZFMRLO/uNgp8wedcSSNAz8xuctCrVsnn7NVK3
l2FaVk6VD5phpQkGgaDn0zmMiCXtNhH2JC23Fqivtwh5mt20vwemFkhCMH6qpngJ4RYNnF7cb8sg
Za4pZZYPN1WpkCZLsbRDIWjINNsgZCYhi8dW4wmIOD7FZ8/z7NhjrLyoIYV9X2W7C0saSWUBfKCg
cgh9qGCBs7mToshKmOhNfOxQA291JDYHZn3ARxP1Y1/dJ3RzhrE1ep9Nx0XpNXcHWA+6xfKw0lCn
toZo/dilLUi+Lqkap/OtjWSzKLEiiZRmZhcqhFOtaVBeXgmCT5NkISEe6fdIWxBJ2yMOXu4pavfV
FARhhd2xQcmXO0XHfwoRpfKyD0AVRR/taqN5/5Mdi6fSvQP6w65ceyLR/CjgLVT0YPWywBH0ePF3
aU7/QE2HD9L7vXP+5cpR+QgybZc+AblcJZq5oOejLSQqCGnI5Im1KAV8rxMfApHcM4TYgXonvxnj
/2FAd/jPB8wCDppJdBt9vwwTwQRZNh1WvFUxbWfXgq1mC+L1+o5zYlpNtACtdYH+LPmU/+41BgY6
c/0Urg3RbCOI0nk911D2hl1TuoEXdA1cFzPfk5pZ+ZFbm4mFIALcFFlfLp6sMasVo3JwMT/BF3oS
F7jgKKroz1tW+N/vnlMUpW7dtRUuQqcwfSpPwTW267/8nev215N2LQPtLKdtT5/DkD29diRJ9aVb
9NkctlaS39amoxrubydoEcWfwDL/tdS76kc9b4seIDe+QChD0r+epkuDdy7kxE7JtjIOJ2TQ2y7x
i+t8LJ4z19Gi4dQ9/8kW3GEqAzhjpb4NWJV0uhx30dnOgxzlwUYQ+yWvM2flDTBEZn3NOylAC3hu
ZutW7Qsj/Wu9CrgVP89dUnOBdbpQ3o+YjOD9DhKx/BOztgQHHJvRKp+0k+ScirCGgV2RcpVAmgVd
5xJhHVxViyJA9X56Ml7mYEvf0Ax4ZMBO9GLnaOFtvKNwaxCzvdP0mrvyzFHTS24NR2ngN3mXomXj
6qsRKzvgk0BN1V5M0pm9F0efN2zkz+uBJNfQlgA4PiJOPHLsPVX+Cb5HEA61nslZZwJH5R0lgIRp
oKxAvSs5sYnOKfvOagGwT3zEza2TofiPB1BcgB4di6KLh+8bahz0/ur9fqKMD+JGY4GdZXej+08g
fORyoTyyJoXRs1e69tMCVvXZEBanvZJiEq+BwITSQrJnJUXuMqngOi6XPufBG1+IdAhT46KWxB8T
1vRJ5GseXFAnQSj5mq+CwdqXeRhXjKsj76S+GRCfbmdb+VTbtwqMQLwy3WaOM8CAMBzYAns+X4AA
MpSFdSGdDgmqfRta1OwgDBESWOz1VEPK9L+O1uyA49ZgL5OidNZ7jx1nv6oOyXXFUC9/Hs7NlLXx
F4F9FO+gxxRUWfToWy42k4qBJLj5QWSwGOoA9jRh+iJIksmqn3XvGfJJ0Dgy6NVm1t7aOwIQUrq/
U/LPKHqyvKKRvga36hu8EV0nOCCQ+F8dfaB5gJzFWZuSM5amt44z5JYNNNeOaNiUGp/RJmROExk7
cL1UOAJFOFPCKJZnp+lzqBwVU7yGBD2XJULba/5Leb5Io8Dfg0RWCs6eHnI/AX1/xdWLRApdPyTq
+/NB1ewkieb2VxHmvfw8zCkRkSQu30DPy4zCyd6xcjD6TJXJK1rMYZuluZpQNbxqBwOLtPUnmAJE
BMgAybeJxtTHMUInmRn+RBsP39kLVosmjtZHET6EuCemc5U2dd5vjiDxmVY/ST1/KMWziWzDJyWp
etTs/oraAh3RVb3WwZ5P5p7giH90o1kg3H0i+kod9XemfHSkikIF4aOCq1Ip05D0VazME8zY2/K+
NSq17hvQR4m5yXvja+Gfl+z+VPs3o63tgX8uzLwYjiRHbmHYFXAyI4PthyRC6aWOM/XrfrdfzeGa
/BwPE+jpQvsG+sr5m8VkeTVQji5wfqxN2PrSJfX5P2vYw+ARrUp+ZIK/ONrzZ7BN3wZwCPDJnH8G
Kq0NH4aCTApUoR16ZOCmYUhT6QlJCnjupr4aoR+3QUEL6pS8rjbdkfBIoNHBhBms9De06up8zeY+
6RIrGmX+eOD3JK66vND2rBwOoqSGpJliJVc8J7DvZc9EVS4fwzWsdlJTcfAOg4NMShWL21ZIliG7
1lE90qXoQKMHTuzqA6YUmHgtxsM0KrgzfSBuCYrChb3G9ODv9Eb+zASdtfqgkWmBMrUO4pkbYv7Z
+X3dlxSolAvhhET3LlWTQRv3TBUV1ovPuJLbNNfjpOkcS1PANtQDNQN6FEVvpL+SrHIv7hDIoP5T
sEWyFCW7sRpcfj/zHu5PpvrgCehXG352AYC+l7CDb3escm5d06O4AJeeccPGnpsjyZfwiXhCP1KZ
HcY/DKaByr8OHM8z08Ofl2w2gCkRKorsS/TIGPFhx+bAbBmXoRrI6Ae+xpwc1WjYh46PtuVAed7y
il/5HGzsMfWK1OTNCGMXax0ZMKQXUK4V0Lte+O905y+Zvq1GRa0IxxY5EkGK2KANQJ/dLp7CMKxv
HEpyHY5YfuD6N9Qg/+jSLOU3XHwnP04eX/e26D34FsHFPhFOnvluHVM5Sa/Yvvrx4jwkcS3wjr+H
1bUYyhYwFPx1+yAjOw+8h+hmnri977/XQzxbEXw+uIBJnw4N4iA2tFxrkqMFvmabLJ41lymmhZEd
EibsVhG4b5vXXKmgik0TuSYpc52vh9H6kdpICGTTm1BeO+9UqymFDIer4wtukT+v5iGckNtYabvK
wM+/YZKxSxW36hPsDoFufOB2Zr+2kRK5V+acVivfpEUZaWOVnOvf6xtJoAppf/Wr/aCecE+CoT89
CY/mPdSnQZbJZEzrQYFojPBlj0PowNe84adCD5hFuxZB+b7MQQE5tHxcjys4w/7EbhQka1YiLiHi
wJZaGFbS7yYDeTiBHTQbCt2poYxSp2d6dZsAuy4rs77AHz1AtXYHVO7Kf14tcTaNTWXo5woYmw0F
Aq6yV4sUNk+EdvRgRvvHY5jaXJpF6R6kAVoYuYpnTKJjbIrrv3nkqOT6VtR5Au29mH/kzBitChUr
l4K6HIo/pReYVFR2CZOuozrTmh6bKLNZ72tRMrrrp5DbBNAlO7myOxfdPYWiwM0YiaRX0mcn3U3J
PcMRnlCVzUlMlcMR2T8D38IC/4luGXsyc4Eqvap3pT+CDGPvfdd/d/l1XQofxHSJtv01HtmkZC/9
P9CFcxqx3nwoo0fQsiD4P6ZbrY2Db2g2WUT/Cb8DtowThu5snXrIBiW5IKGaXd2cwu6AItuHFzVi
+IKQQ58HbatPvsm7YnBFGigXLiOBaAfIhGwFoxzkHmNvYa74FE/mPLR4RmBbiMj/SKLoVw49LtA5
iF2xDCjbMUjNUQOHvNif0koodogz63Ncj1q72xNHeqb4L2SP53+PBiZA40DRJSdlyX6CXsEUqI9N
KpCPFYD6nb8RhcP0Q4y4QLpMcjUcc0sfB2WkY3P6tMQu/CbQcffFivYO+m3Fe7oF7dydpX15FDup
YvGVS+Ynqg7aQbOFakUzTwOTusAtMd+oqGiH3m5IvP/8pv6zvoDloIaPwrjNYtw2iFvrQOa+Ap2G
8ugFNVyFk+vVNSX6jIoKTTP1zPjhak4/1ZHxzxDUUmFNt4bH7BzrWZwlB7PBJ9pYu2X+i1BztHX1
PtkuOG9QWdmwnSu3ctTTc9AfuYVDMnknkmANQZG+eUroN+Wephp3hiposyuIDOINtV5vPAuXehpv
N+yNrFqFBzhQwj86jmlvXtKgCuRaXMk9yLe47aX3sNnvCWBhXK9QD1mVpwBAQ8wq5keNnH90vnos
RDdNeAWairQ1kC+tDvQQBuIKwLmfB9IZQlQ/f4buZYUyULUO9WbGN1AEDZ9wWN04MB8E503nBu3j
DnGsmU/CnLVqE4kAVVVjme/IW2Io1j3hrriaIeeP7B0lwLMPTek8vZH7c4RMLu0wIwUOkpYf9FOw
cpeHvECIBSVQy64gEjoPbSt/U/GTjou8petexFXTvMlv8FSRpIKmJK/a6QrG7hJvXlF+ZptRgAXu
MnpwJNtQd/v7fIjw+04Apob8eaBnRsxR7p92biAlYD3BeCce483q9evXuxWG/u2BuFr3SMw9R4NO
HcuH81l0bSSV7/Q2JNTgcgIWiTg1Qfwku5kcOk8cTa6Cr5bF9eID0Ldy4JUPCnfatUYCGXzWhieW
flc+/+O1X9/J6aYS/DHLbiK7sxPggqwD7Izt/21IK4NEatqgeYKAdeN3rU1f69B8I02dRAN0MqgE
wg2hitx8vJJdoc8mLCz11wsWnHZk8/t2MyI7Kczf4e3CHJn7Xy1R5Z5gWmfl6VEefvAFzA5PkxuA
0zWGJDVK1VF8j20o9x427vOoYUhu2LLCC0SoDuWy/iHImcc2DAzeD4m96N8PyLwUsoqnDB0kLTex
x4yFfWcV5CPZalRX/ejN11wxlsCjmraeeDlNjHKepl9tu5ziL+0qiUniNPDYh9YdlaHG+J0Rvhkc
DEkxhKkf90lxSk7Y5HaE56zeulDgojxvCGCbW2SOBb9lBcXcpbahRcZoTvUzaUXDPBWFPcy2Sqtl
N54tYYoynk6D6r87IfK/Pxg2JsIf1z/1PoQrMnHbTSNy/CzLwONWpjKypxWwuGxNJ0ALvLahHYnb
gGnno+QLUhCiA2O4YT9KMb1iZxsY0uoqsFdDSYo5+H1KFCRBb7FwUcmnENds6YXuKL+SKEWg5FE0
UAtBhQHAHfzfTprL/Fo+leldvFmW9hrDOCC3l+fxYAS2ph0XgTxuXp07k3hS2f9tWzc4VTErcW3h
ULLhVHXg7+kNyUmGwtNl/3UtYlhrJn4jmcDBPDqU/OLiPRUj7sd8IRY23FA0h1dNbyBJXaadlGF8
3QGDP+hQsSHeVl/YCTKFQKaolY+sJQ4fdn+vQ7NJsYfZLGQCwCsuf/Fh+uuFATOJKASgPezUi7ob
kvMoa3KA13V5T/7i1WOO1/Qs7Avr8ghZA/FkKRNA+UdmW3PetBlyKtDnBEjEMW9/MidYWI2UPf8U
uPnNj030/ALE210c3IX04VEeadXZ5Vh2Gy37XVzqv1sgQa4E3exnnSt8w79zb3C7BwIKbtNrc9Dk
I81CQbBrIQXSoGWZL/gn++PYEm6GO44HSpOf+o7y+QAdUdFW5uDBUQlamG1Cb9f6QXd+1vdaGySn
Talcoi1rxTdEjYeWCuEeJYXYXgoAL85tgSQ1Rc6FSLij8/piwIINZ3BdxPQ68ZaF8+bFlvxiEy6Y
pLXRB1CzcCAlpB8EvwNUE61vRdHyL3WzwEXahmVZYp0hUi4TrV4xzVV8eoFU6i+n8BrAQfRZsMPU
hj+yEcmGK5KpQPlL+Dp9qVgWlSPU2eeLqp1fyPythFx6Xd3dv7f2HeaPdY29szYJ4naFY3lYs9WP
YLLMUhwe8CAWVu8Yi37cnGMGCR3p8UxDg9cIqjUj5n6N6rc7sx8pCgsfuNooKDn+yoVCKezq2NcW
xvid0E8dOqrIrxaw+YG3mf3jhv2TpQQ3tyg7YfYLxzMCDkVreILe0t8rmNN0GeVWhF8M7/DcHChT
AqAE0WU5JWU+lmfU9Yo2mhpp8+/gpsuaNruZRz1QILPdgDui7ibU+lDdG21Ff1nPyjo0oA9zCDds
RTmqD3ojkTY5D3wPVpTEGnEHhzml0W3mIqas/qhcMC3RbIZ65CA1zopqXT955SktZCaG5f9cGg5u
4jSRoxrYnmE40jS3wuA3fwy4uyMLYAXkAcxLUiuAHqwgpG1kXY3sAJ4qoGeuDxzJBAwUlhBXTtTP
tmELrSe5EwRyM405v56ME+gf3MgmnUY1K0sxVNq4y1waVbgEltZdpKVUt4gvxtDYOxb9in+X6BW7
OUB/wsOnlhRsYDjAEUaICLhQJZcffnQvw4xukZkpWbFjL/a4WfsQ8KJ8zVmut0xRCyr2AvBrUkaX
7pE+HupVI6W7VCdsOhoaU5H6QoBE03HUbl7UfWHlqpFKqFcs2F617zz0ryIO5jHHdzc80cuz6jWy
f5HvU4GuplnPtZieF/j4b+qYfOyQ9N8+mx0gmiw31hE9Qi5B/KyTB/3A0TB9uVQAsQS9eXrt85Wx
zyoD1YqRBilA+7EFofQuEg0AZ5/VsWn+H7F+jihER/XSyX5PlnbOdBTAUoDLPe/fRM3Hr+2Wx9s9
YlbOv3Jp+9Za1IAS2EbvY9s0TTvYt5sm2CiZpujMBgWDb9UZLC+kGytFdgCAtXJxmv2vg9+sae7L
LPTcCbG+eHIxGCBGHvHO7+Ua+dFjakaeILZRZaSny4YEPil9PuPX3kt4qhtUoQKbepfVkf3X8AmD
Q31B/KtS0uFhDoBIjEfLXPqIjCLUyXLrGtgYzbQA0WopNWfgU2MwOFq2jBC0p94OYAhse0tomIpD
thxnf0pxt5jYw85y2cfGAee+nXHN3hW24EuPar+T49VZev0aKwi76P6BJy/BvZ7TVY/Vh0hzTQHQ
zX5AdWAUyMrlaDGHx6xoqWdU6PYVC4X9XXd3GdmBOTylPJx49HOVvWO9y1QoIWSv7OdcCWvoE3Zj
/PE3C/qZD6HvP7UsOSdjcGoi9NwycTDvLLoLhrrS+1rDPZmL0X2JHQ3eJ8klUsOxphGq4gb2M45e
kXI3RKW4AH7YCf8bxHygzShJkhzGsz6ArZiEd00/l0kezkB0SuUwD5hhcIuxZQtObeQ6sZT5eRHx
RZAph/+ZWk3fuP4fcI21C0V6pW8l6myK+2QjfRE54GlCKmeuJjVTdrPlW7f7ilD8iXLkThZ8ddF8
iKdUumYhJPdwZFMRaGqku7smXciLrL//Rjscl1d+p6sL/ZrbM+NiCN0xPeWN3MXIga0N4qK35kTv
A2eUUk30PxOpYQaT7xqfh0sydT5+3vOHPdpfi72VqrzfA6SL1rmuWThNrICjEzr8L/Yal2Ny4YKO
wz2NNs7wCfVXMl2CmaK4u2joRdqurKu+zHAptErDfy1M3nKdfA5pVqrNbLm53iiddLDCOcg6RN7M
WPzBIgkzEu7hiyakTaX7gsKjU0XA0qwnmVNy9CKmNmZOBLuLksIRJw5NCQlSs5R1eU2nVOEGrj+4
zcsp+Eo23kgLmwrbHUgQspWgMZl/Qceh0nxTU8SfI2iCeE7ROITAM2KGXZbwM92MkVS+tzB1AF9V
tuIgJpzPO2Bi7cWlpE30ABTTfcc1OQq8AAtvs/Opkw8KMdA1fl1cshWs3b+4lFnhcH/m97b6nhUN
vOwJOAwM+MLhLmbhuYEVkcdC55VCQGWR7N1FT1vIsUHSXZcQIHymryYduZ7rsmIhgo+xs7NHmgdJ
psX/4qZPw0rWjEi7ciEK/3yupEg08O7RmY2QY9pYeX0lTU74fkhFQiGzbEqO6mu3rte0srwKs+lp
fWq+BiP3/mkXGy7TVpGWJnch/tI/dvjrGZv3n62zmbBIM3HxDWZIxBVVZ4QsLsA7onxnpRbhTzl4
+MdGpUOmOB2QiDOqiHtHMIUFHRK62bTL+W03XzWEoDhJK8krShOmk6gRr0+TuzBRyng2XorbYAMj
nI+iU5x1LTGOhQLguGn+6V2v82FA2zDvopVa0N9ZIxFtmwiAnugFLnEhQM8+qmG7ATP6oeqWpAk/
zRVYYbd7PoWWYmWHGRhHn1PARw6gU246ygEGOz25Du7SQHYX2rHsk79Hi9CuQXWxz0z1b/HiRofK
acLWMiWfZyzBN2jslUYO5ax8691eJumisWJkRn82oXmSO+ZIxRNjpWcw9HQK8oj3Ylv897ie9qb0
0wOh0yNU10bJeybwx1uQzwwvXylkee04tUgCZe52wPk3kntEwoMlJFk8l/62qiV96j7aRTPsyiC5
JBjeLA5beappL9ao4i+0HwA/3hpxYIiQVTtgNJJdk/4tRzLh+EZoQ4HvlmDfa5hQadXp9PKjaomc
5+jCzVFUzI2JYdyl+5YaJFztRMsmYFsxjh3X1jdeVwnqrjO4DXKY888psg6XIxsKskmCqudNmr5J
5fsnCSyND6BUD5ghCqzva8NAXRb6LKoEpPClMAovyKhmjke8HEHqSd4xPQxaoKjL7SjqHXprC57J
JF5/LCMty2IIjpe7Ub1y40GnRUB3AbDdeAu3Tkf4q8gxHU6uBxH+h5U0nbwHMFgaKVuHURkatYqc
25XVAPxWMNBNWiT2MGeUSCE844HGsXiHRtxySeZhdVtcHAPNwhL3gspCrb9EYNDgqS6kIjHaym9c
uqvxTjMCKHCwvt147SAMOSFEu7KPcbitu9Cen2mZ4t3fFTCQ/0MAnLJ/ti41Sm+RyaQPqaWgOOwx
6QmNZtEIITEG0URFs1JUfvZuQLoPuVz75LbiFRTgSvA5q0ZzeufUI3akkkKcjYgcZo776WlDIPHA
4Xo9oZy0iIMmQnqEi6Fx9JGV61mELHnnKVkmYfegXKdQRls60mh61dM6X01CQqQoCSGcwXB53Mwk
cOizC1Mk+ehxk31uWfNprQb4fgH1x/1w+BD6smTq1SZLvHjDGsJoO9JaA6QjabYweEOVkF2iPw6O
Mzhsm99ThQ0EDIDlcJEuZlgoQ+u8Cy8ynKnYYg5ayDBpn6wW559HX3Szpo8hPu9WJROb4vpl8Z29
Uy5GgiyuzzYsrT6jOubc++7ZPBBtAsG8d1+KnVGW1sFn4s6SJLG6G2nEV1bHW+bJoEvPDzg7SqXu
m7NQKixhTBwTFVh/jJNJLrWeU0/HdMy5Z4HmiSqGoC2JVzBkm7fjBG6KX9YLcDBHgFcCyGN3UYHr
Jmad2qm+7dixovIwqw5cl0P8lFONedWbxToLk8b4edauQxwz+uxr9N1KEqxWqLld3oNnQeNLlkyK
3J7NhqktDrSBUi6orW5MxiF+B1U5Gf9I7BMw5S7IwvRZLJJYCw9CAiF4T6iOv9NIHgd3zTMXNqIB
N9Mp3Hbk8l1J56L0t9IWnC57fF5ertMO8wd0V2URHGHCdO0NFvzB8hfM46Fb/uC+Mvq3xyahONvz
7ElnnONZsyUOri3XkU8fLsouWd5zFTBCWP6YMUNAtswBuvdmLjb5B4zVSe+oYQwxVqFMRrUqqbtz
tK/mf1YC2b750+RymWrdhDug3QQZgbLr5UFylKACoLYT0dCx+8zLxVglu79hg+b/RNzDS/J7Cz2A
6is4jI0c2NFk9kOEJf6yWCYbLFIQy3oqrWzqXX4BOaRMACo8KxXer/pzmWGyAm0efuKOgyuXMRab
NFsCRiCq2zQyGQfE4kW9pM0jPGQvUisFbuWCkhK10dB9OjhcaGbFepduIka2cy53zGXr6/oHGUPi
wnqoeoNuTEbvPxEzh/zO7fP0HkI6K1HekA6TkMRmXmLiwPtKdSfsJeClEdwlsBLEU/N5/i0Rmo6b
pnt8NZTUYb/KyvC37aWuh9ThBZLLNh1Yo7Qx3GQeG7LECl4SJw2CQGg3In0vMSRAKJzrR2IQLQPD
OwcxWWr0bIwe1HiqP5Uo8JDShAXqLDriBcJzxrDSDtnrJk9+mUxdJ2o0Rhn7LS2Sida97L8vScBa
RGC3t5Fi4iFjNbjdq0y5Gn7viZkZOymQrCNFsB4azHpSpgr3BANfsmdcLJSwbhqnHU/kglpQGIJ3
f1vJXTSu1Wt1x6rqGOlO7seeAWk6o3XK+iec5n2KESfUqLcVeb1QTh9P9GWu0yR8Aiv37ENh7wkx
dj1sXHJLuAnZZRw18+ifONB38ZAGEf1TLb4Ikce6FVHwDbBo+md1X99SrDYjHyOB5UrdyfL6wpf2
LkeUdLqABOmVh8DY4W81e+vMChwH8pwTHWhhDAG1pSts51bXOPDAF8Ad4wTPt5IdHlisd7ERutAn
j8/4m3pJq8Ynpeg/0YQTOd9aK0Ggiwiy32bF0XJIydlcEdGZMksph7UqC83C9r5SGmPgjh2Vlb/I
Hw9MOJQ2ukli8wKqgw3tFaEhGVSiRByG0q6dvlUeoLHxHE4rYjuPd8b1ZB1C8FnGSrds1LSIyWDa
9qyChEoE3tQNQmgt1KJKUnKaI61mbng96mwYqp/5xP9FkL7lt34J3COtTHTSnNyUYPQ40jU8SX9u
YUgyHwuNHQO6vf2sjAb51CEveCyaeEJZQtFx2iw8sbjhOo9H4ikmaZOGk0o3I5c5tUZoWDK58Ck4
4XJs2Ms7DGuKEIJS4U6Hh/BvRjWWMtes2BYcnfgb1mi9JVdjREe2Zm+o8As8PS626LfkkDSEJamr
AOpLhxd+Hob7CIPdNyEzmAcFyHopu/q2R1J8dSrrJwAPu1Rj72kQdefOyaqYjv3Lc15xu+YtmaFx
e3fAD2os8pas+DV7KIiso856gFAoZ6xmVkaYGEqQB37iTZlz9wQit5a2NTjz2LXGF98XM6BcnbgI
8Be3BvPxg9J/eS+HLX/uA0uucYmZmkkYFsmJNAB/M/jaysZCzcAuCmmxn1c6NU7ML9Jj/yp0cfCv
7CdOLzntdMmfElbiQi9eOw+r/fetcuhfPtJGZH73efT51Px55omHk8I1Yg5/Fbf+7/ilmhgcOYUR
i+GH6NJHKmA0Q+peEm0/Tli3AigqlMw5hxCyuyzodUX0ehDJmOixxeEzcRfM99C7UISRut7xiUau
JE5RSLf31EC4wmIRvq28JnmduEPA2MURPXydgU6pIMqwVcGjr+fy09Ksv32iI7/O5ZDPA3HVBD1Y
tqqu0YoHkBEs+tBfIRv3Fp9SIzrIwp5W1KExI0nAJEY9oZ5LKYH3a4FiM0SxPt+ZMMKHCxqBmWoJ
idzPJFKa+oS6lpWdKhxNNf2repnJdTFJuO2ybziXAnWF80BtJ6ApO8Nzayjd41JSQ0kNKiQEqfAJ
zR9Lsr/OsN8krBGFLauiLFDY5CMJC+Kbb9QsjpahOZEd0B88iqtGTs2ajasffeadbUF9UlAuiCkd
A6QxKw83rWZ1ku6LbAh9iv83SFrsaX74alWe6zLwRazWNo4RqlAKFcbCjztpnwBx//1rSYPd+5Ox
z2GeewhI/xsXq8gGJ08VvLF4Tb0cgYNqSrbFrQD40Zj5nS0TxyjRjv7OGBo3XtJgVXtZPHkSVLJS
wzLg/YuKOUwnQkAXHKtsyKjLzS0DpAaJi/YJuI4YVbrySsGHFEiAncrnG5VRhACmg2Eo7qNNQvPm
siihB6CIQ1dXLuET0owtTZ7SVyUTBrpc6RdDr8rKNIYcDvToWpugqz2466Vi/dcs0s5L0sNDEufN
eZ7Ce0te1mHx7YzNJNgxuJ5sK56PRv721fTm/JcgMhts24Lh4a+BIpyWPf47JokCtKLc1lzpZj/q
8hGDBeROn1T71H7MBhkhjRrv2GRMQPF7Y2Qz7o7V0/kxcFcQ+7+C1He9HuE8abdvm9SIZes5a/zg
XdpfgTttNkEhjhsa80RlUiM843F8wZiNjUAVFe2GcMFe/gqzFQ56scwUFXV/J/ujB3ZiTDM5tvzp
Q+MAMeSIRPoZ/STANywLq63OfuJbHoxLR+x0ju6oBut9c5vvXgtsgsad0i4iZUDlD8qD9oSc3CWY
crP3YoIRYhKU4Pw/2F0jkxDUrOQbSJjXmJsE/GDwkuWPpy4VmymBftNNIHhKd7Vvx6iXBq2Ysdtt
zpd6iZW7nKjsRj8wMTG4J4wePNdWHO1JufhQdRBEt8ZcWoKrRLDFZs9l/BCe+36h15S8g0SR0J3J
X0HGp/sFgbiWNRWByLO1o38ycGEYbzDRPNUvaTOSAMRHt4YBXKIDMpl/lqcMMNvVvThSnAp8oDSF
ElVC5HIXbHPAlun+9bkHqJHnH/S8lau+i0bkvgg+CWe8xtZ7FEfiitKA7GOXLwyFNt5NwKiv8jFO
sjGmxgNFFFOLTohul+PMfzl3tFQvbYWYN4GaBNslhLsv/Do6s17Q9QiaFa7+KZykTrLZBK7cUFMo
A6wbnS68cqTKSJI7XDCcO9YfRa4wzjOPZLfwRUko9pTkeD1AvQVPV39QR9zgazmzTZqnEfSVUg3q
q2vmEpTt0Sdfi9vAKhbEUXTwCZLv3R5G67El4AabPm8BSULEUOO4gouVmc5VXuB3601Pah2+sOz3
10pWTNDHrj5OezH+rsS0Nic3hWp9xuyeziv6RKk1tBwIyV4LGfZnctNWjop58ASiKfen9ArDplhJ
a1bVoOC+vR+YlrDdR66/VplWphq52sezAlacmNLFj4UKseI9fvPZMp+In/2hwEM5KJeko1pID/ez
v0F+8Qcxi/S+W7AMv7hwPOkoc4glz4HJMQ6sJWQBacIaKBVCLPD53YxrgUbMec8kwlY/etP02Hbe
yAHErsk+5eL4aNg6fwVnyRtJ5ZJ8lDW7JJNHOusQs7sMpnRZnRP3wY7otPir/ArpRdHXkoXui2v4
BNWAHPLr5gOlYVOYeqxJRd6HzY39J92cFc4/knzstvWoccSXNFHfU7UTxoSOTVcg8JyrtMLGRmUs
FW8vr1xF0qTXuPWcGCcV+zp+LAwyfOHc8yw7otH9ORbuw1edgtu3zOwYnXCm8ab5O8v1QuTPEgRp
t+jeBPOwhYD1bWsc+7CJZaZ3LRLNO/ZfZg75XERsfmNgjpLJeiM9mir4lDLwQAroEipmPA3QO6tN
rRvRr9z512z1U20FUcF90ngreAU/ItyWJcKPuq3FKetnEezIjwFeZbriH8YDOIHSYRf9idS8N0PF
lmc1geM7oNaigeRIXQzpOEhVoJWNGZ/869t1SN+NVLDpy6r5mSJOKuIlbMQd6gQdvkDzAvg11TTj
qQUfpX0JMooNhhPxK6zfU1lUU+LTEienE/eGwibhEAovevfydB6/0LAf2JNLkPAxVCr/ov4yV/9a
XSSn+0WBzt0DsAcdJ22U5ifVaPaNEKHXlD3pM34T5uJ9ou1PprEjjIWINcETCdca1QSv3jobJ/xM
d/gTdkIhMri4lzgC7zmUAmXDFVY5Mcaz3fs8lMPgkxohSb9kxV1VTo7R3x2PHaAG5NQL+k8BBKek
cJ9yLb1LH030y7sflwu1c0HnAwWvVtYPeTuK45kiQWn3QVziawRRzNRFcJ1Be1PTmUdZzi+x2isZ
Xa/6Uev+Z4+SmhP0dHIIDIQ+4wvO3I1BwILKPiPdGR3eQPetCUyhZ4lCryUQOR1pAUXY/GKhn+Hk
z/FOF3RCaOSGg/sW2gY4CJ6QTWJOYEddXu+Zebzi5BwCQP2K2EZnZsvc3LsKizBJO7Uf4E+p1TUW
hb78vlR+x6SGSBkcCwg7pP1sE8pvAVMU18LXamSFFXqxI4lduE4uixxAwya1AQd70O15p3J1K0AH
gBFSU3UKe4whWU2EUQ4Rh3rg5/p/Vdau3rfZOU/IRGeVYzKS8DPDHLWSpiUPUJTSwtf80u1O0h1u
XLT9DlmFYD+1VFU3wTz/DhIeZaGsOc5yXeOnNu6ef1Johcv1Y+W5BhPF2gVRgzUsP/XFLWbBaRm3
hBqj4HSgE/IvnLKVI4ns5RXfqOejUJ9ZQ/qEFm9xeN8JWKCBVkWQrGiZory1Xtj7m8/qxuzOHZMN
MXKG8+rvs3alKYnZ7r2amo5n0W6w9m7cxiw4n45e/BTRW7SJOHzbEquaD//UIW90nlM/iAYpcSGL
EoLryUOR25RQlVyIk/BdWEpUkL2qTa/eTj7VUZlpKEf6qCxDtzgBq0mBXQRoPyk+0pwrqZg1l+3I
BlVDeSWVnQEUwRFVWe2+8rLFkk/I6fzyt+4GbhBoTKHo6bFSli1g0H97LW4kfg7+ZKt/IG9xeDhQ
YiYZIivPPKfO01+0O4kwaaNfYkFvPPJixnQ3sgxX5MmIjhYd4emnUD9r/D4qVDNAGThpaAriWwbz
6BObIO8K8F40fnILT/tqQu8ymkPktAzqcKUyA+RIzyTtz6rCCoQy5f4qHngnLZabI5Zhh4rLKDTb
ntFHM/eFWkrKw2sC2PPBNuJVsO/3unvdceh3S86XirGBbEem8xwIjnbhP/w7H0/MbGsTPrpaStHv
fdecYukRKjpWWPpbGjWUqY/gggDX0ADxVaXxsGbgR66HD2sF9wr6S5VyHcwKYebXEHrrOSYkBkko
nxRsB+CwWPuRGFFCVrcfO2UXzRw3bc7sTkOBNSeGLrCbL0PIPrPIYHpM4KdoZ8i5nB0ctMhQ0ScZ
AcjzWlQ3+J/p/ZbZMUtjYFjUc6HK/1db99GSfRpTTKbFYzKeN94L/ecSv7QsrXZ2NCzNrzQ1X3gb
mliGt7T3GcH/JfN9XNBUqAaS5aqC+1L6Bn++LvSuFxSRGnMy1fpdpqEMmZ6VrrAvSTLrFxE8VLU6
D6Yf8wCD8jbxWIidgPpzbems4ztS5SL61vDizpf3HL52O9s44U8oNItXY2tNTm4DKZAwpDUbOO2i
RmIXm2lmKfc1Ihh1woxc3wL+TGEs75knXIzs9L8dNjP8ZcPmPsNdTLkzFuUs47LLgvjTYqwicdNX
HD7mZSiGVyt/SBoA98eCd4d0rdFZ4B/GhsPNoNNk2eVv4ZQwp++F/ETdStFHi4DsBS8u7iusBiod
LcfMU6oclIVU7mezc0u/KlGgXp+oDm9SsEcaT8MbkQ0/MbIjn8M8I93/26UbbYGAAIVCW7mr+794
DwXcN9nMn0hlpceSEyKwECfRmxBJM7kIhbyKBUKg4Qs+Fpm7MKOXTG4qMemyXThDYF55C4gruEuL
nFmPNcZdkRWyjrba6ahNn1oRnZ5qNZmjqxRa2cfCXDUgxbUwliVSHYPkCpZqa1qwNVVp0ilhqGXD
zRWtDWF06OGoXT6K6168arX/gTiHClhI+k8h8sX89jSjxspF4alewuTXGyFNjxmF2tOG+z31pTcm
6loPx7Z2KUT8i/4zv99ZSMPdqWn2VpAOHAzmuAsSEW1eayKZ9YmFIx2UrQXjYoPF5QKf5eZxKnlX
B5lSn1VewFBt0OSv5/lB/6q+sPSuTJpq3t+GIpErdXWa0Wi+Wi43W1STHVMtz1PEBLWhAkY6xYOf
7WKRlJtGerWTftW2nrR0Zh3dyKGr8sKTgKglXekcB5R3QMWwTmGd1qaBCkfS2n91DSvqjs9eNGZE
go6ZKEknqWq7Qr1UBDqjSLsYrNTOg97Rl5+FpbpGIXB/dTW9Uzhe/vOgxS72QPeSiiOLpcAUKvIR
Y0ANNXzqmepzZKdpB2nDnuiFqZfmWPgQ0P/r96NfnfDUli1DtuRWOCinuIOjHSBLnrn0/TXrOzha
LDRKnyAa9iW3Jx6vaMHYMkbCwmX/Xwv4LN2KJ6thXNHKZPUWyPcIe0RcLPXHkaxgUJ9UXu/LwF3v
1155UZagEBKK78o5WdSCenkOcFu9Szg5njx3tSo7xxJi2ue9aZwX5s6kWEv0C/LiMSBHZGVMG46Y
XFwk2jt4Ow84Ec2rBAySqGV4wULLbjwBYIY+i8x6AC+Ie1Q2/mohtG2N2zjHzgjHCOWYehAq73qI
2PNsXatfWlm3cf5eJf1L7uWXJVVQVywpKN33LZvnSh2pzWxXCI/jxyTV2emNt807nyks41NWP5nf
F5oBWJaiHrNmYxTrD8RfTF4yD8AmGC9S+fd6TUT7J2MZ76Ei07MAsUCPF3BfnIA+BcPB1pWu7j1d
sv9lWLifSv58b1l/kyX0PBC8pQ2OoW0HcmiwKmbrMrOi2ftwvHHFK7cgerG5k7Th7Sy0ZklUd4Lh
0Tp0PnZIZJSDx4mgOOb3ZQT4XqG3b4VtT0HB7eJOha/Hnmd/xN51KnIM7F6e68cDlVSI+dfTG1QG
A/5MJpJNg63QIG4cXwuVMRTegs8optlg2mUm48CrFJz02UpWgoh9LlYn0W+mHicRzEY9DspZnM/a
i7qLusKr+Wu7tFdLoCnabG4XiisOw5KPrUFLipkbw0n/p5TwMHdMU0OefVcbVGZ0XY0Tk8wQUmgb
1N2rz0TcZfITrGN0BkMZcRkRv+/sd+53ZBjqOZuzP1Fq+akWdZVLXL+JWcZsy8QZN8XyaY0zvQtp
P34qkxvUT8bWi4bhBhy4sfa/XtM06S8bbCGC2HGhPlzEIviwad+pbEp6Al7kVnLP0onRSza7YD1d
6mUtnwywxBST14HJQ/2ZSOj2XQ5vP1Eify/bMyBddto1Lw5YIL/EB6grFGYnJBAmOSIC9dnGHUWB
igf3B5FUDHNUFSlaSGt2gfkQ5jrjwH2r0qJDyC6XyXUKJGdxBKoYWF7bbbh5N1KQuQJKfs6v1isA
pSWcctcztaScXY3VomSsOflxCu4tFhu2vRi7PM0nVLn+pqs/WdVBJ8iXAE9a9t/ash5h3X7Nj5TA
btzYD5+BIe7/YuMRtqxU4DtCgCpeI6dkSRu9xQcMVCWhR0G3jSTOzB+fz5DxS/hKS8qDpBqyNmYy
CUvG7+doQkk2c/Myv1yhrVs8ztdJuxZ7q0U5jkpIqXKmIkz5T/1fSOO7zak8tYw8WHh47oLhxJkO
BJRPWaOd60Ic72OXcK1kdvi2HXl2HEYpXuZeCEQkniQvIIb+4TX1CyP2uGxXjM5ulqlSfaSHE87p
ADl9cSi1QRHBz4vMBs9GLokaHvmNy+ZYZ8j3JWGjideMX6AxTuw6fPSC0Q7W0ZD9Lp38xoXs+28t
fkNwmFCyaaFTRTAskigED+1ykqG/eNInwWZVkek6LS0RZ1jM29FpSHBYwegjFQlcZ4urwnB+TdyZ
1/2NpcmQJIaLYkxy4x/X3Vw9OR7Y4kNgM0R5qh0aNRyw49I6R/7YZzs/Hu+bB8Jk31iOnZG+FXpD
4QLr57knBg/zYzguPgawL6TqahOTpqnea7F0FqYzyJ2j9HLbe11Pwju5i5jp7CmzRViwHjtcA53v
ojftgi4W2Et4HENENQb37rnFAU3V7ZPDGbnMFwMCwsdkp4TYFsu7jLjJO6r2J5EV6otiW1G9i3pX
DNdFONy/D5LHWYQmQ0+50282cqGVLJCHP9RfqA0FSLECqUdjNN9TwbwFWHGTN3RL2AWDrZJ2pnaN
60+zqKB5P3dRmfJBoYtPQe+nKTbZ4SmFxbuIAcXsy5+AKC4duTxv3eVmUWtNr7LLwFeSsxYAbJDI
Ev+elQtZTTVMBHQo7elx5epOV5dL7bP8Kjqnjvb8w9diD6a7n/4qMHKSy3d9vTQcTGK3sYRBkTYx
3Za2rwZUzt5M61HjSfhDqCPpyb4jc1HuoywD2SrDd8omz+It1X82YGkZsmoU3OuZ6ktYmICd7/SV
7djKdeANBPjm5m/2qGf+DLOqkoxd4NTB5mJRG/erKbSB2n3+xby+eu1D8RpSwIQUhqjhF8dlrHsF
lr6Y4jBXd6mCeZY1dY7kaxyJu1im2LiRf8+BeLMfF+QjoBk0ynCaD0zlC0FaigHpFfLK6lkg/Nqw
FeHpGwkAGbaZtSglbaGkRDicZcp1MMMx+2rsYSzzSqk6Ey7PJ9qIfSWQMnEPeQbI/dLYlCHVXBUL
eysjig+zQUvZ7bAi0QEskKQIHYozBimceRAda2G0ctEddW5i/nLN2XaA/ulqpBRRXLfSwlPK5BqP
NBOaUjLdW9edYCoUwltQpjvuTfW106iJ/fMwpfd56WDWIwUYHXmgk1dEHkdyfa1sbpnk+Z/b83cP
PRkGnX0nzhzPfq4CY49OKYTOIrZ33MlKre3JuFV7ozYk40F3vVNiCtUidfpZH8UOlTC4NEMdfu9l
IZ4qq+F4ZTOLJnCYC5vkAFtvL6ntrdzq+4e7fSyXfZVwQZP6hHEn3ZSmNjXhHQwU62ml68cAYZaF
6oHDVTdC5KxwTZEUBPeTCY4V35Da0IshFOQCDkucinrxrCIaGMV7sWyCzX2oW0z1t9qlohOkpx62
IDlVXoO7slkVbPBjq5r4r0L2msojzZOhzOmVFaaIqW2eun/rzqHGhsAs5S7YyOb/q9Jt9W1ifdGa
z1Txd3UxJBHlGcLsfe5PnsNF9ZKTGHXPHBAVU1Enyil4BYWQ1WA69VnBD7FaAYz//s8fg21XkfAE
F+atTwiIHBMl4+V2cUjonu/IbLuaCbGYpVau/v+98npaVpVhWRd3Jjd0PUN4m7OurI0PC1g9xo0a
GdxQ46lJcl3w+y2glgqihYoribvzOkKUqua2ZtkMSs1+nh0OyRbSNd+PCNAhbCWDThvE3ZjYUUJU
YeQ62W8ObdfbEz8mUylvEoD8MMt+qH9BQbt79PD5DKAMwIzTXevoCMDyhpptkaGPYXAcBuXrelVB
A+rZB7h5Vvw3pm1+MvPry8XCwjcifEVOPm4IzpwoTlph7q2vT+bfDtW49e+/07z0daO34C+0BkVt
fwCfO5NPBhZB9e3A9tThjqR0AVU8dUGvQ9orZ6YMw3JEdY67ggxQIcE2JpcRKJdbazX27uz1YvVZ
kCW50BYFBNzRHnisk1pg5J54ZBnnlh/++1b3PwBFTFDM7ETW/JeyNsYd5pJKl8Y/yKcDJZvz9lqI
Mn6C8BkBYJvNtFE2nt8chdg3qq2pdHPOzn/5F2he14hm/iJ8EoFUXPVEG1P4R2XS9Yqfbi3rHGTA
twlwklX/0tlScmEdv3zHPcpAr/to4SqbGzx4Pi+b38SLF71cJTAolrLgF8JvD5T5/YZ2A6o21OrD
mYWeSTxpDgqxK3Jc2wVbKLlUYFRSTZoxxkw61J3b/6GYGdBcYl0kwukqJpoHlyUhG+dMdiKo/0LC
bXu5WD9oDapcDEBlvdGm8JhTwTfQLaskrPd6C1KnoucBOZpLKWtgEOoh+1TuKsRXHZ+kiXCmOMqF
Z1AhKwUutqVLWUGFv4D4JYlLTXo6xnHivKtTGEZklU0EwBQg9Im8+jQ6EgxgdfJVlMDJdgkzI0SA
v5L8RaxnWau1goRCE5BTWlvsaDzVQ/OPrOnNBCC+EkusphjrPwgecy7wzq3Fn6N965ihTg03K9Bz
kZ14yjWjv23WthPvJVzuijoVDgJAQ7hqW0qVL3IBzMzb+yyWDCLcaBF6/lc91dyci5sxXAqI4S9l
uMRQkUXH1oiQQ8anMunL5pyL+uM6UNNIIr/b1pgEH6+1Hbr+w1ywoaEskENi3oi3gjx+C+OJsrVj
hZmmjWqDvJvUlZPUpHsRBWh2wjcqcY3ct8HYyzB8v+tnCvZvrtYPB7GV+9DnSpeIl7bR0gTuLXQT
5+vbK3VYWyTvt6P9/J1Q15R69ruVvhulQuD5ZRrVYzTloKOmhI21wFkaDVD9GeZU8pTxhazgX/b6
u5nZv/n6jg30we4z0DI3liaLSvP1cQOpdCMzkO36AxUkwUfjTuUd4jHA5slOhxLODY4zaG2SNVPq
6stz8Zei8vj0lfNWwXc00kqicsq5JCa00/2nciW/N9hbF8rj6HS61AdhUmtB81QYeOYTOK1uBkjM
8Pi5kfVgs0JZznnkN8zUyBltymQ00zpzKt5HU5kOKoKKt4EO59Iu10qp2Da2dIfZQlUMqEonhQhq
nSIK2Hszf1qdcvO6Bgt1XzTXO4HpBkolhlor4ttoHvz417FzAdC8+/3YrYqm2Dm0f9xR33zFMuVi
XUI4/CKJRnB4/LRALlZY++5GgU7jEby3xnUsbkHCTbDtMt8QFetKrhYTYhgeg28t4pHzyfaNook9
tvoOfegdd6LcAd4T7YZYQEJk9V1IcdrI11pgtFayrS8+Uf5ZmcSu8M+VDS3g7YH7hxu+VUn/HBnx
zvA+uB2kCI8zZ+IjYSLDGFqnojqh44+eHksdtPVzptxqcfxshzzJE432TBhfAtaevk5zp8gJfzF3
OeNn7lftOHu6J8wrbgck2ngsMXi30+IZxi+MsW79wunDhJ8xWqbEkXzndxTYp8jTVbfGoA208HET
5nk1PsqDoxYZ+SyjNPK4EM0Dw7LhvjACR9EfD8sf5c9LZWLNACHW6vJQ3KFqGG2PZ6VeSoM4LJJj
TP8aCTOD0Ujb6YRD5XyPKAo90VCVctCV9Ip8pQGki2JR+WPtCmTdopuwjSjnDSm3VO3nIqOkas9z
GcLBBS7z4PSu7w9q+ddHYoDpqyZcMulg5+AWtO83TFLa0xCa3nI57F8m61ZuPxySuUz7EUPaGfZF
bh9Fm6f59ChrNv39qbq56Z22XQH5ivl38HAHVCPnI3MVkFcUK6aAuvYgHOWFz2PXtIYfU/+RZTik
jmkBc/kIDoW4IPuYR1rN7Mg5OuCK70ycRMEQo9PDa3B/hR3zQZlRdkkhdGu/QA9LJBEu2FNFvPGC
ndpRad59ZPKL0oouzOC2r/r1eHo95JofWr91Hl5yEo5nrhDqgDnLTJaRei9oY4Mtt5owJGfzr25l
7itFne8+lyaPIBmuBpRevlR60lfixAT1ondsIA+0/7NMafaaLRfCpIRAj2ipRZ/QQvnSpZVYD5i+
vjbE6zAu28clcT7FV7Sko5BXzzZ7o7IZKlCjDO59HtDD/G7n8TaH4oshyyrW/tba1L+yxrXzcs8R
6DA/PrZRnRLz5/wlZwXJ874jPD6mO9FZUxjwdlmKb00+H0qcKpeqsfsVGthWhsue1EZg+o0q8Rwl
adsm8wv7IERUHX8tyCue20jZastD8AQRlyhtOgmRCDokGwNyJGzdwqWijw4z0BEgobZKmUTqcHvX
fGCBsUdg+NncHTzTQ+f/yJd8oXEMPwv9CHZRMjVSWLL701stzpkwR0BPIkBaAppIm4QNBCwewTP/
Ci0TZxN5BVTEEehMdcUZxjZ9PQ4UwYInDbCSIGzsco34DNNAA7fQYHxhIBq54DqIGNxTzqUM+JHB
6vReymYR/OO4Ye4scMPSednOECdGYxE6mYPUzWFPHPl7LGvp6ia5VRSXhyTNpbQSLpttjZQV5Rvr
YrfdI1Wcg5/0HnpX+RTlDstMLyFgQch81J6e5w+NoPzYTjTOsUXhitq1bOArK69uPoFJNFJScz6K
8jYqi0rdSMexphggcgNfZUwCBO5irAKz5B97gdaJb8LdjS2udpxwHIAWHP2s0rxaPkG9aSvtq47T
2Yi0MSrsRDJrqTA40Sik14p1oRkgo6/22juEB4ZYe0JekDeFkgiuTGVZS3BEvgr0iHWnqTas+QQT
HdiJDhI4gzrFJnOaZa5S0KnPWWQGfWIMlkX0MSRw6ssdNVkaeFUp/hFnM6PDwEY+UoEYiH9IgYwp
k/zIsC9EibiGr+HSDPyO0pnLOAr2WKydZApWjpuyUnqB6zZJSJD9Xp7JHnqepYD1zVawUFFjnS7c
ro7SIOyEQg5DKElBFHVItBkZiItpLNh7OQBacikNfqs/UwcXeqTKlRyDroMfk2Jf2c343w+PIjbM
tX9TjtMSz2RNmgvXolPmAiLvygZ+bIkbgwR63lCshODS7qOP15qiAqJ/j3frPdrHCk1C/5epyBEh
MPhgsTkPMVUXOa4IeMAMKT5+homEbJg0c+MtUaZ0sdmuGasCnfpZtATjQvpoaZhaRTG1ETO8lEcz
KXooLSc8M5O3PqknronfhgoXBb18T1i9mFJSOwlQLldQB9aiEbxTJIltX6lt+T9hjsvnc432djhi
dt0xoGRBoojAwQUvgY14Fh+Y9t7jADnwHt7W/k9HaVgdL57OcHMQ+5p2M2hhYP44UV2lqm/DmK/3
lj//EB/ZVQXvk5sDOlzz4HSxZWhata+7r6E1BPD6bNQvQGsbjsx3ehGd9G3hqUsB+s4pqjW0Y79a
EQ9q6izo8z/7LGzajvXrIm9apETayknRTpEQnxR2duTP1omF6E5A0JKz9m02EU4HWI0e+a2P7qoc
wKy5wNrOqpSU+9W18F2q3Pw+YEtRjhQ4gjF/XSwFl9XWOAdGQymUcx65Tg255XjjVcSTy397rNvI
vZdm/b6uxjWdNKPtPDVRmkeL1NcdDBpnX7l6lzsJCIUGlNsys2ld+RxDXpkZpJgJ38sujDaigJ08
NC6KpiIeYOfc1ytRfkYqQRPxOkkrZ5AlsusyLyRSb1dW9Nhx2vXYX7bUlh1xyseotWGquzuEi8p0
P7z+5odYLq9l5HHEZNzujKs9/6hekTTRgnD8qws8zugp+sYL1F5aZ+tMQjKdvMf0MlCvkVvlTx7R
Mlj3Pw0S/zDvWYp9o+e9Q4GzQJ3yBBIms7DxtkZZXrROzY1pZkaGP62InhQiQ/YUUfdLHamI9rST
pvWyKkJD7zdarscMz2nOwA+fsQ2+297M2J7Iosv2MC40dJZuiwwOBKc/QYD9sWcy0a1jVzHyo4v1
O2GNk7po55Gq7lhZJnVMn2r3o9zT1+YX3tit/WewVVJqCawnKti7vZbq0DwEtWC9AzEFTi00G6GQ
geK7ddoXfvGw2tVU7ysuoIbxtb5j+SIvL7aPJSsP7WXsMrpbf9o9UmtoELIVdysAOdQVu/lwBRCq
uJS6JDG7yhBVVWUNiZEYkHAXSV6HhnhovMgTGkHid9gR9U96nL+XT9VLdQFjKny8g0G7dixkwIEl
YByG6KFsg9664qrOkrPQVNRmRUl7PKMivFkYuNWlGIr0kMq7PKeja7CJ4TDoc3NE9e06ci8s05ru
NByQVNEk4EewrX6bnwN5/6rIwsvWu5p1PnnWz1Lwg84w5niQDsSzLFdY0ZlAN3eAPDUft4QAWS5/
+bTLHua08rdomNfLP+nyUv0ehdBENJCeOk7tILtyRTSUKwGL3xVG2LBxga6F3N2mVuBbf7RZkj2+
x9k1MIt1fjuObKlYMD46Un4+g7GgPEtEs1OCYFjZZybGxtBWQl4v41K3iMhJ3jzJoyaOFtEHrwMu
hHuHBD9dNu5fe1oK0PAaLK3LLseXL4jKvD74/f2SHy0K/Q15rotjER3GKWOCTh8TC2vbSBvgDCd8
Cv4S1lqUJb3zbo73jAYDFM3kKIcJ603b+VGJn9Kntea77yP20vZTt5Q3dc6rFtWP8KRFSP2y4oHw
OAeEb8eqnCALsyLzDRonLd26s+hdgkEx/QPYpc337LSLUid2MDFiWbZfvqjAXh2gbelQpF8UaAe/
Sg9yY2/aV/4QFO0VZSP0AIOxIZMU02Yf4GFA/l13aoXpzhHFsRIvqpEtTXoEu2NtmM9BdKkE/6w4
+DCJdmi3dON89unsjm/1jNBr1+BCWOMXAWVBPEtxYfw4THz4EH5i8gFNqsZxyIY/qy+gQw1Fj8qH
QlzUbxiOYCZbtnk4ZnbfUY5FtLDpj0fPMBRMi6iSWGOwjoxU5Ebry1xRkXo1Ss++zNUStmrw2mwY
mAjd51ogJLGzvRw/VVQfb316A/d5/Aky+YWBYUKc7+KUo9kps46lrJH7AkxtDgHf0BMyZDt3gDtT
GXyWBZ9kb+Z7mdRDYVUBHpTLvMcIJkZpjoNdNMoxLQ2izhvycvjYB3L9AqaMr7UrdSC2G4VprUOr
14STinInF0mUlxX8Lar6BiSFhadGvZX5bopsnHYibSJtiLoigW3AiySVAkQG9D0L3/hBkwq37dzz
ecDZbXpkuF4/ISwD8+9o3eByJ+TkF6GOhRF4C3/PhcGSYmEJKDaBeG9rb9p3iSZXqM8kKxsyHqun
a+9pGfk4HmbjaBQBTHKdPAUYDVqRO4c3WKYFDpBIJg9fl1TzMxoSDNBtun3pGxJVlfdNZAAuap0D
qrrckOJQXHbFRVpSgtgdMN5dulhwOOc45XwutFL+lSBouHDnpWNVL13faorj65qE4f36jN2z9GBH
00ghVmaJ6kahWCOsjJyzSxmOnD1D91CdFIuBGd06jzSmWkWX33bCkBsnnHlq/AIiQkglTRuSMqMN
6SYAAH52qzxRW7TLWkKGheJCy3EqC+yn4z3IyxvCIZOUWvVysD9Ea7ExNAAd5bPMef4KtvSiiOi1
220wKoEgADvnc10PVmmIHYerDvujcCdiLFeicXkudG0NTulE/5h0qm+OYulxq5vZEWIKRy0rOJA5
fKdAtPLfMj+UdP8zsiyZQ1m/xjtnju3Dg7gDDsCBeveT2n7dfqw1cpxmvWV8yxCqbi892HpoNpi8
hcOwqEh3tm5cuzPETwNZm67DKshZWfzHaah4eAKQ43XyX8dPrY5MwBQ93C4pjAC5MrE2nr6jfPK1
hrBFdBJF3eOsjVg1b+cbpoEb9deL/19LrizFmPQwIu1uN5VJPJ16BWlsR+LdJeX8jTUUXdQU3i+d
q16rcf+IpZ+E0wx+4/bggc2xsY4GovgFopghsJ48wceBnqAsSeASwlT8Ua8NqjsIEtLoYPEgaDX+
c3DDYFi8W+WEnw0ZvCjekn8SrK+FC0tHDShB7apz6D1Bl8uvQMtsoWYVxEI+QYyxGxCAnYwBfL1i
XZtzKs9DSOTuMcWPDWEMspRPXTAkYVV58o71GPE3Zu6ZehUfDtjV6xPeW/IIQlovU9BAPAFg49g9
w0mkTXGf3XbsVUMyKOJ9ms5MhMBsVsCXYIdJ24QHvc8DSsPQ7tQyeDUZhGp3YnhZjMfMF4ampSf6
K5ebU79ompCgSYcwOnaCT7jsmjdU9xtveVwBokJEdLkvWZNAyjml1Fn1W4kn55dDk71m/PGs4Qzl
hWmHZqwtzE58Yt6PJWvlnRBfMedOdYvz/ltLTJMik8jutI0+jbI4pISMTlqgCHnWHGsZHs5MUJeF
8ScGYrTkKrauGd1Ltut/pUuhMa1BDmUj+f7ibbAnuVAvn6UcYRLS1iDXVKBM7Z/4BGiDP6ttVN9e
La46sEF65Xqp3Ef1qGFeYTF1YUpK2n6vNt5aoV1rjyAYkqX5mB6E6RYz4R+bHqMoEowi8Y34D0gZ
GLMPYMUxNvl98Rl7YB5B2ESK7I5GtThn3i+5Y46snieyWf8thAsbS69HwO2UBLrKFB6AEdZBfQcX
XNlC9KOHqYyBxv/8VFufpmTUUaeZ70ugUX6N6qss4tHIQ9IQ0PBPdvC2IoLofk0/GvG8muvRuWqT
Ft+K+r0QO9jZq7PIf+db/duzv3LoimRcq0gG//A/TeycBv6JDKnX0T6Od6WuYHSg71qfEZbvqlJV
gWciiq5OWr3kJjwG0RjYy0I37REAI/9GnvsmCZ4QGSIGax+BF8atL8punXDrSan18R29HOFYut3Z
uYibrLf8/MX5uY6H9BNQ3DM7S/KH1HffMzhGiPayAek09RBdx9twuZORNpYRI/es3uiFzDXpXyvq
X7knpoIfe1u7RKyHlvRE6cyxJY0kRF4O7uE7EzpzfS16XDXF9qFMH4BOvYwHk2/LZQtjgbvncuPP
JcBSZK0Xw67Sv1EHfIcQJhiRtxMDgGg/A/rWFzFQit18fwH6gIeUx49Z9G5CTAUAqADHkkg0D4w3
sTIr0n/HWK8mcA5WaVWDb5HFtE7aSa4Vqnb3vm84RsalJjYyL9raDVg641VCw+lDZuEdnJ7sHWC8
vFwQcD3Czxn9tNvODNTGEsd1S0W6l/1DSAhr/1zqIzCAPw+r+Z6hI3NURdnRzrI5r2N75GcGjiOF
y0Vu2ahopBcYCMkkTbOXUfNe0KfVGbyqU4ZxSqgxpezTjSHvt0kCw5Ip7rQFzM2Y18+ziMyKYqys
csS0nZgtmjPtKTWMjAfYWI0ptSpqxJhSrQltPKxRTGQtamRvmkurPp4SAXpGbGOOx/Lvva8jAJet
LEEaRT0A1wT/i8GOd/9pqX+p91/djaYNDCGk/MES/A08Lox0+oIGUbX9XBUEJIr1LwomwwI1BuJI
GERrSBikP9L0THj0Fw8muaUW2RkgSR8GseWFDbwc3mlljrbhQ1u0f21F0B3WO0KcW6nee5Psurc+
Yr9INueYvE3XNEs1PK7fnn1X4pZ5yYz2mEc8Jjg9qgNXa/3kYGArzb2+MLwAZPdeBMFCW3ZnDxn+
kGRVvH/ylKbk18fJxvqWZBp9QAyixniCAdSB5pYKY07EFbtpRk8vCGy34YDrJQLCorysuJ0SBwtg
R4mgaMZ0JX91LveG7O32jBnYjkCAsyw5bhy3BkYv8bQmPcwgf8X7yO7JeSLKpe4W6GOr26epRlX+
RcmGSk0pPayYnYMtWzBFvTiqPMtaggzaoLOOmDqkC1dHEKrrc8EPOy6B5nSuaj7D3fiai/bkElun
QE97kl0KGRWO9Ql9Mi6TiRLTj9utvuhI79VJbMjDvzcSB35Vw3z8WwpxS3e2lG7Kg5RZ4pq+rGcW
OdmOBN3z5u0vooxjAs2EjneSo9v8XMa9XTsbj4W/RaHWrRkZSkmBT5gOzfIUS+3vwSGo7TkMSxIb
PEqXSI3Z0vBqBip9xka/qTOAYVLxk6bGCuNJYAlU5vVBG7dBeQ31wMMWoZ1rIug3l2qJgy3L+bpt
MSsh8Eu1Ye2SF+AKNAT/JBeigF5dLb3hlUdRm916YG9EievD5shWie7xr0NA7tIkxWDlpm6Xxi6f
on6m7zdFTxugii59S7nC6LUlNjtKBcFIb4h4aT7d8pKoweAA59jD80TyxTgL2uUZDCmN1ewrH1Tc
rgmyCxGyAgqCwsKJVW0GLfLmwnew3l6nrWDuM9S71zaARXr39tqEsN1gi7YBXjbweqPtysXBMx7Y
nvacrABzsObVN5+2oc8FESzQA8aqi6oTk5LDAryplwcOjgZY/FrXZIzZPSRqevy5VySO5BOVP1rR
usWCaiNDBI7L9otKFMVnOqpzd+C8kYmuNH3xTE86Gu3jpPm8e/PjPxOKT+V/M6n+phVo/C8Tv8qN
D0ujtw8Hqj/S9eJ0rSagomYHN6rnlHw+AMeWEooDe7a/aHEpK5STFJiSjW5DE+aYPaKU7snZF0w9
yd03Wv4cyvSxh2IjEfnarZqPWf2FllnigOmTxhekt/3u8BI1IwzXkTLriFV1EppvNtcWi0bSYACz
Dl4lvLqvHtlv+2CNV2SHFKn+10HBnBv6Zbgo08YNNNwPQZIq6VaMdEovR2KXSYzoPIfu4nJOzKtj
B2lis15ql2JPVgSrKDKFshJ9ReQ/QM1AWA/hS6iwNaW7ZAQ/FleXhXpgHbIEKWcLb7pHL2eebNre
wwH1XOwOKMkoW+xgqWARmcOvqsDDk0Ohi98fkI48PLbCymYOZoC2LFwKgzg+mOcdmFV7pViwZvs2
urpRpKHGm8jaGzKCxKSlLSO2VCCT0DgLAg+V/hNTttCw2/eTXpSDSs+K2SlCCfcuPVqrfwm5V7C/
EhT5lmNAkv5VD0BCQizg9PjlzpyLs6Us3klnb4juGYPL1Sfu8r8mPQ8HeAN3KmZNVFazn0qaH6u1
ibjVXYvSfv5cEGPZgRakPEN0uJhL3pMFwIb3/UxEMPpAiWP2l/C1BxVe+Nmqiv21LQrNLuxIxJq/
STkN9c7kynOBdJzE9fIXoFo3bc7foD4Crwz/26GEwZfMcItch6kcnFJm5q+RBvjfFb7PGu25Ms8t
fxUCbPNcDdVFgAuz4Sx/tA+Ge2RvE25/FtGoWVQmMj0Swx0PzO+ywdCqsGMDZjFCRARnA665EcPN
Wx6iSF/b7Gyl8AkZP1lRETg2aGvaKSnGfPYQ2SB3y5yG6fhSFvoIS3fu7VaTJpTxoAvy+rSNqxvO
X7AikzLyJX0XnhQPX/EKCXpd9ZDY7xgwuTosjsWsMjFcAFoZFaLQ21E+9Ch35yDAXBQO0VK7raZR
9ssizPzvIOWFZucYY+mSbh/iua49NxE0bpGBjZZRoRTL0enLiU5mEY50KpgSYWrTe/CfrWWsNZ8q
HBib79O6kxIXVmYvdpUg9ZECZXYNGxm8vxv62zF+5YuzLxG7zIx+8X1BZjb97oBUVHywIhVaBHYp
LjOIdcwPvyeh66KL2baQSREd9MayMlY+x1Re/XEPwYEEqNiX6ySkaIEpihXUJDYWBrafhkkDbJzQ
TiMBBp+2G/r9QT1g/N6AxgCH3rAFenwgGv6MJINnUDV+PNckB2eDNT/Cbj4V+oCeH5KHWCxtx0Ts
ro19NQdxIqHehZ4oWOm0nhUYZPaZ57fjoXlcvWSIAuD9GFdpYzltdR/HzYHUrx7agVKNsO4rjNwM
x4kvEIlIo1Oc54GDIo3TGAheryIvo5wJutkPmdZ9JIS/a2EoQsfcTTedD3ChGHM8HDFZHtZy8toh
96aI39yD0wGOd4nWjlCAQxI0cp7XK6oRAb8sV5Cy04R2OG8/51kUMX3KGkM/cUYWF1QmczAE92oH
/UmHdp17ALU5V+d8fJm+VvWBEwEe6L7aT+TzlpmHznRThg41p4FSRhUvM/G48SRC4sGKi0ggXLzj
DQ+11BZg6THEsV8Q5LX9ZR8KX/59ksA50WiADkqQ0nHXtGGUC1ierb8l4puhKBbX3i0fbPKmfYLP
FEL9zmpq1Q42Ayvt3XOJEkOlOOHiBv00fzdp6ggA+SLq3B3o2gEhcxSSsysZc6oSFO3XlugHBKIx
m3gjcScohBZXBl4WdqU/OToXs0Yyf0WP0HEmkAldCSBLGQUj8RtpU37zD4O9GlRA8qMnbtdb6C5Y
z/sCJyIMdQCDDNamDxZIpqTL4/6Gpj1Z0pCscvdBRmfOl4UWJvQYhjEx1wlaBq4ouY+zJ/yoL2Ml
RcJrJDanx+bCbrHGdDdop/Yc1/9sq7Kr6+SBETVoKkPw46ptvu5WsZBKw93SXjt4iuErIoSR6IeZ
umQ8Klyy1sZsRhJktr+8MHP1MpMbTa6khSHIkZZikrxLWPo8aeEmKxRdTSZjrxxCSZwcAVQ6W4+r
OsfjasiABg20oSp2Rc4f2puvJFpYKFRd6PBGqgQcMWiLJiVqCpQ2uzgnycQ+qBdC9bWLJWwBbER6
CHw4YgUVr6XSSjTVArdsJ12Hnl+HmJTI7eCfZ7/9GxbJCy20lLhjs/9xOqOmsE6ZLdR1T8Ld4AOw
Djoz9+ZVTBAlzI3MIEC/fNQ3eD/duTB92exNqUUl+unlKL6ZFJeYlbdMzCm5R92auF+a6KwskuT0
EE99pACt7DoM4zr6e3navHuWqz9A7O4kXkAwD2T24XH5x7w3b8oJWpdq4FbW5shuzhQA1oRAR6KQ
Pz8QfTUEMHaK+CHG6xByADX0njpD+NE9pp1073tR5/jq7l6dWqP8p/+enjsU2QDJtWMHqNibHxmL
TRRR94a1GOHvUENJAl2QSAIjDLzxhWfvRo/HZK96QlpXBz4DAbS0NJNzOZIdF3hwWrXzDg6ZjBJT
ZdueY3AId/4tAircTiU7rXPzZHH9bZBW74dZB+WSTaQj0yyT8OnoED1hU8NkmOtmRv2+D1uNP1FJ
2UtDNi6cWLbcOqewUn1FmjOxB26PhoCrPAQEgqAzA5xP2+LCh1RDiLhFk76xLFI2idMgE6pY0447
0xdvLJzdxAL+0NfUCkcFHMcgaDjML6XhwTxiF81BU3lxDoik3il8mjOYYXbpwNK/0Axx/BGRyePn
OLCRT1USllwhbQQi6F1B8E7crfYhcAdsZiKTn8UwGjgczaTKGCFxtlpoqdK6GxCiKD+VhMKl1/gt
zCCQECvihhwhoDLUCPezxl5s2oX1N/7j2sJvyJqtEf5mu4Uj0kFNfXX91KirBLWW+Kem8rV0TUgQ
2WwtckvMvIrx6kxAs5A26njpIrX3u1xbiZMcNgyug5KNNwXbVU+pPS//nBJj7GLP4lyStNKBXmP+
PoxqTeJumBiCivbDISZ9CIJhQznEjzC1QuiocTEZjObOCcyiOjdkIHasUv43JeS9xNWt9letN6Am
L+2bcv5ZBkkZBDOkGruLCDlFyv6BC1c+Bf/5JnTfqh9zd5lYcEp2vdC01tMAHJL8MJsP2aeuXiDs
d9P2JGFqMl7d0S6Idp00IEMadfkfFjMBpHn5vC3zVhUNuwBZodVITLgIO8eNzwNd83cVrB1qkAYr
mfu7hCZvXzqXoFBVtDAQNsHleqYIlvDLSUs8nVnqZqVfhhmroNePEkHOX6OMj19DPQD4xEElHWp5
9O6w/ReT9LAYy2QAe3cVgAnzZT0nmGQrS3aHjeHqr+GgePEwANidH5mLbJcybc36nG7MqufChj4M
MGDqzn8J11BK6EXl99IdSKxbSw44q5+kCOX6e3KXIpyTqv2QnVR0vvpyU+Wxk6wRlIftk5O2N+wV
2NcNsKTIUSq3UliBHy6rBciC5XWiTGkXT5i/EfVUwShrbEwdlnYNyyukWcIvPl2/y38Lf9Y/M7k3
IxnxJ73txuKdDKceyYRf5JPgk0r/5FgTPh3FxRdCTeECi9IXLOqKzY1NIUf4lelht9UXUIEy/pH+
QKt7XMpQ17pWtH6kXT6/0viV1KpWynICo9KGwk++JRXS5C+j1hSlKTqipvj5dagFLOkiNOlGGNH+
KDCnssptKT7jVKPEdNkyHqS30ThgFV75iUIGKC8rr97k7PZdvTQpRLSAuymRXuO9S0nLK3fmO9Z3
riNrTCJfjWUMv0c3GVWyl5P5NE81O5Fw947Ei/qvY2+iqyoi0cl7ISZUieWaPfNbr+nQTJaJ2rcA
0d7Kt8x2YagNQl8/xEWmoDh84rTlcWxWy5yLfQnGuLcz7xO2saKi2q0Mcp9pCj99tBDdnEJ0bLS2
na3dnCvJzy7TRSO++V2b0XgZ+ufyrJvXjYxgrmJ7msQ6fNXqSLhFwhPc2tQDhunFf7Gl14+00dER
XvQmWn5qWxwk0JZZCCk7eYWgWLUriEYMr9w3+f9xvGGPRDFFDVasOf8q09qSJQN4SwlGKWV4AEdt
RJoobiVfx0tZD8U9oHB+ABQJqT1Hws3A+NyCFBNPHs6pUVN9VG0HC3t6e5fjgXyXZUT/gXe26FR+
9Szh+EjptV6ax01iPbzrkzm7CV3HzAWRpG3zHGTQ/dTyrEOxycaYS45ZpKGWkGUnKKb1bHRaW1oH
eW+aGgj1xNu/aMQQBrODd+exiRiWOU+/MuT/eFGkaSFtyph7C6cza3d44KW0LJNxmQNz/m5f/IPu
XZYPcXt10jOy0s9Rzyn09BcNZ1UvvCMn/IxVwXE8N6wStQMEnebiqHKSxoV7//jZOvDD6YEPbJHH
XCrpgCLfi2Nnqmhkg68dHrZdUg82AxgiI133zbZSXAGiXtHolvU8qEAWZxUypxVzw+8oMyTS+rGB
MdlAoIvXLHsJJ6w70uciN9R3RqU+lqtHzg6zbBxhmXgVSDc7joFWQzPse62ByhH0i7psjQXJp+5X
0UvyRWCUUSfZ1fQwfYSLe/JgWPSugPwn6p57oSB7QGrPQaeYtj0WMUlipJaKIeofxrkakrnrZ4E3
EM0udVokA+e455tRRVYWIBBGxjC3mPIOfus5Ye+8WpKQAjk7d28AZLVwxV2sYCeq13VXLNCknfxE
7wFSiSVTFAYjP9pg5wzys1Z5fe+h8HFTM44IXQ8meSBI+TSohC2g9b1qPYFETsUaNKC2Wa21VYr2
s3HohS7Gn2KDFlHkfPZIs9XGoZrWV9LpeOM9BaqQsR1Ha/FINF8YxMiy7Sx4Qeu5rGQJ2/Ntdbz2
i4Pkq6HiYy2WrNM3/LKsdbwTW0y8lcYypTGbfvPeSlvCCfkPV5j5/D915uAotRdPQoqJhFtLs80n
IhCrorR0XxQC1snQr6UExEo7GV65MCO1b+m+DKHG66qe97WyL6rl9fRmUwE15N9myNv5VNmZwj8S
dGKlT45I3ylkVDuYtrlGsImbe+qbcVjX4UA7XH+OIoHj4jFviHVNX/IpQuABX14V8h/oJrbDfb9a
E6YXAT7hp/1jHJu4oUBiUR7yxYEp7t3C8VXmBAjkchTCfzxXZiXMx3vt52AE1ta8VhdB9BFKI21U
oPw5t6eJvQHI+NKskbWZvrK42fZS8R7lmDVPxcgL+AgLOpAFAH113+4yhg2HYZ7a1cGMjY30r0Nc
ijkrYfSffz4ZrwV6Z2E4VGSY89KlhRTYfy6dsyb9BFv90XnLfoemycPFXyd1IO3fNlIRiiLdJNd/
yfZlFN7D2Ak2oHpWzHZOVytrs0g4lKIh8bFd4LUk/btiExJ5YZx5m/dJlbfb62oe6w6Pbo4/q5J+
75awQymk8iq2/Fc5HM96DZZiMvEBI5SWfTjnjAVoK0mHu0MUahN5i/+aVaLXNjWNNOp7BWANiBII
7fElcLy4j4ydzbBrM7MhuC0HRUCD0qhdAOAC8Mw+0gMua1+UJrEuCXNcpVFfOsHDVttdVC0OUzcy
WKWyDGDRg2ShHBqU/BZXqUWzCXpMga4QXPBKtqSpCljkIgF130tyRRDeZmN5LLW++dw/uCNf1GPl
7bV41MAfS3su4wQyDlpskdu8Lsc3tCtYck3sAx2MDR9Wtc7PUy3uVwfJg9FtCpo3yb0QRHFQGT5z
RMovxm6dcix8v6wpnmBHYNdJ4GW8P63MjCgZiPOvElZEosQQhrmM0f1XaZZhHtPvIOKzmMvcHGUm
AZzz7C8q8ctNJvoJFamu9QkKTaYC726BRFtykHElVgCbLXTRruYj0PwqmpcsmaFu+B5w/qeiqo1l
eT5hkWHpgNKzmeecrPL/JoaCHOqvgicw6Xkl+ejMqLfrzYFfQZ/PktlmcwalQ5nZ/G2BrNwoE8Ef
BFNsUIv0wi6cSZD9zgJgWls9C03RipAWMAPppNjkmwY0LVDX9I0AE1iS6GihKLCvt4UJXIjaEfOH
dZfkpDIJequhKZGYSr57OH1vU7Xr6blLIyPhrutMv4sQrmKbSzozoZf581DSbVycpYzyrI0BkM8V
RcLiOwPb10zrh9IRjr+yvCUmOW4IJy4pH9kzgV3Kvk2gTFGmYCx5MT49DYGXaiQRXwh5ACAhgH+D
rWDEqI5sZFP+9IN9QYZryJcelmMIbGTBGAfVpxJQFXwVF6hriX7tFIBAQpS/+vXZiDyiVaFFGobL
zSiFx+DDC3Iztb420Yw1/AKZ7wsJ1Zd4eqG5M50oBTdO7wHUTVKfK4EPlSEh8zdmRr4PyPFMUuyB
DWZOsW5bdFozviBykTV4e1fAI0ITULzTlkdEVkdVcyigKUasKMvURx9vBlYxlshjoRFpSWxeFP9v
9WLoLOhMSL0uoC1uQ1mIKcG3TF3BbYJn6DNZo4Lqf/8pAl+j35kp5Lb9N2AFJ7qxfuqyxaG6xlUM
c0j2LMliJwN6hwZ4YR/Afu7RBVaHv6oEr720IEoj5Xx+PlSp4B2CN9xt3LgUiCW3KMC+lFzamwL3
QX4NtU60J5cWDW3xmXCEC+VPtVR19HIIEwNugQqrB3JUKnOSua6CH7QZa+Hc7G4x6gs6YfT8Ywi3
j892ouwjxw/psWgBzuOE9uZKn6aTpSsgomYamJlNtScP5hgkcfjCi4BIVg/CmkgWKoNF05Nv/9BU
Hn8+LmjhHaZLjgBbj8QP3qwLO2+U/pkb4DcoJQnqY9D4djFt3uAzVZUBJfq61sGcY6Q7qyHzv1Uj
Qpt0/gbNNYeBEIjBeisn5g3hrR1Hpkx3GP7I39vLckPKxe+9Nd85yV2cKnjo+hwVwk17DwP5XRpW
9VqHn9xZCYeKbuVU5V5rXv2PcWqHOr/sLv4S24MPHykDCDzZxreTc6gui81BYYy2TPdRPq7o6RVQ
sd4ew7BgCkEe4oxTCXKBfBprziBlSKdFVVOwThsu3qaQRnzUPYFcST3lwrvQg3eCMTSh2k9g22gZ
3conrOv9uOa35GHfhXKDad7n7b9fKo2UzCFWhvtR+WFO4nacF+qDyThhAwCnJdQOh7kHzwxr3VRI
CQYlSOYr7+CuGr0AMunjkHVkIjQl/g6lVefLk8wjsdf4kfPqU4EXpuhnYyB1LKZGxgR8iZOAmof1
CYZEihC8Y9VDWPwps/YYwGnaEJWVCvDvLIGEEupdAxLgOHTo/239Pi0FX3OkWen7KWZqb0TbejNJ
MHkHb/uKRtYISGmUZ2hpkfhvOwtbRymWoRkM5U0EAq2GyoZ3zxZUvpPB/GFYJaerxkWm6yQa8Df+
IBkxrm5ZjZhdkH+VSlhCOWiN5PfPS9v7YdlWvpadyzqmG7Nn/+WLmY3u5iOi3CPRxq5PBU9piH9u
LlxeVDQvPGOpIe9PWBBW89VP5iovjmxUo+nj2rQG9FQbqN6m/5QMEsVcAaE0Qzl7calSIRBgaNaK
UjY3Yy99JRBYFEQpgAvH4hdbijarEccwW12YIUASEshIm5DblFAaTzcvYRt4NhuxVDJYTM2Py1mh
2JZPN6BQXfHSNz3QFdzwzFhu415SmmAqUttBuTKd0TIVklKm2bA+pk9Cf55CFzfn1Q25rBYfrSxj
G+q3XoOZxQ55eUIVGwXVyYsS67ejDp1+jEDDG1q3t8SKJHTVkbxTTjTK9+iqMUCbDtfKlVR1DSez
96ls6VCHMfBSrTeEbqqWFAhjKb5FDBnyaEQ2Z6QUgIZ1LC2RwVKeVrZsB2K23CgoBh9Az57Jo5hF
A/eF7/ZX5qmfcChFQGDjZIHoSKCpYaa2OfOsCsxgyEzRTsNM+nZZ+Q+TYr3Bu0TIbC5ggJ6veWa0
y1ksxlerh1T8m9iOCM5fjwcim7YXvcNAA/ZqHz/W+suAJdqv2dO9zH2YFtyuLjzepWHgMOlX2gJ8
koX/Q5fkftbmA8xmokuKf2OQKMp20RHe3axbAE+AJzhI1QM1tYi+aJlCeM1dMf8fJmODECK57FtE
SYxYpaO/8Yi+woZX0Fq065CMvgsX2ozbKNuJy8LTh89ICDHZy/tmRgecKPHa3e5fdZyGge9dVYs6
6th+U7cOAEH6vshdYdPxoH1R9klEA6iFBda1RiNBrzmRL2V1M9EEagQ4qQydOyD5C4sDnKSBP7GN
cpt/ztLBE/z40+AUjQkOlccKIIapmzJXKBLnCdlcXGNm2SKD3zK4fiiACVsVznIBPaMsjf+0eky0
PLOkbgYCJZVgHlAXzuiT+VKm97hBEOHn8vi7X/K21td1/o3NBcDt5t78LfDhyR+Edk3dZa/VxXop
xCZ1h987TLNulTkW8PU9sCpHl6kfLouMJ5rpaxa54DOPyT0HHv7ldehVXxZ87Oi4XfZQckgGqw8c
70allHqGmT2Mv19N6xoZ+L/Me1rV/qYAoh8UdPJZG88SlrwngalrSbJRKuLIDIAj2IV9/z/CO2gH
hrvNBZ1yPbngKuBbXci1tMRKZ5q+7MBgJbH8y5KdE3W9jA7bwGdnhF+wdEiNfvBPGFZo2QKiEfPJ
aKBLUUuIKWVx0O3MjrgARgm1Tpm/pdA2xr4O6tv7ffMcX0kepsgw8WTSON7kgKEDldhU8RW7+iS5
VggdY2igwUknqyvJsAsGvOAYc9GQtu0GACAFbhk1sARLi4RkriHymO44M0fjPR0El0AlNz0xVaMI
uoix7YCLN0M2jArbKxFiSd+NOlnU4MuaBr+MvIt2ujj18GduhRGrFbIeJAErbcNzSnObhfiO2ZIK
B2/ETmZkJGPPo8saP9UUnuVgu0CGi0MJ1N0u3LP/Y4SkLzLTpc4cp+ZMaZC7/RfIsC95ZpVbiTGW
T1JZ86ypoc0N3XeRIi61UcJOYuuhxCwpNCug4MeZn4mOjRP+Trt/vIp7Cs1eOXS7WQgscOD3sVhf
hH2NyXsJuU8hHCP2NXK+hlmgM2yapeI8ZUO+EoVge5p1PvE/6Lb5y3/AFX5YSGF6lXIn/YvVjor5
szbbbjIeySySAL2jrGqbt6uV7YuD7p6eXnsDurQTElHHAGO963iGhICZ/roFa/w7an+hvMMr8G8G
tc1EV0EJQf0A5ObMBnWDyhj+Rn9TPHc88ZbqfBPn+TmlP1REJgGU3eAMD43skAYnViU8cNaieK+r
WG9HHN8vClDkpTYRpNA0ChNu+KFSaVbrX8C69ouSI3lRjmFnwoLo21NhnabAYqF8GQDad6rMOVYu
vXGsJDa7P3R/o12lPYEyQ7A4eYCAzypEYz36B7Zu0iFNBI36/xwVzalRnWFlzeWur/MSUQoUoy/T
UZNZXITI5YERtThbWIn2VKF9TuydNvqHmKPArO6EYjhfuPf08pXEYkzLZ8/JoKVi5y5AFx96j4Wd
5jnp3T49tuE2oBbFsPvq9UVk5wtUXvvfb8ElNLDnE2XKbhvlP923YbGsJXEUzR1CfwXL00P34l/E
JwJpKTogI/t6Oh0L9FLTFjGDjLU86RlinJINQtvAnAc842ld85pqqMqnPVScwwvWA1eEXo+KkD5z
ld5F02Or2NgjoeUF3wHdQhsyBLuZsJwv0dmQGnlLSInLXeSSxrceAT2eOzGo8ABU9M8XGHSd91PH
Ts6SI1ksBNPUGw31FiTl4Q13pZIlZS/tZIxaMjmtYU3+ll40efD1vS5Wtt67mZuK18oeslNCvPtr
TGQAwS6Ngg90hoOAPU5dVE8IeXnqgWchL9k5D7N7htcLmdph/LuXnXHwBvh70xMZ7pW0Rgv0JEYQ
VqA7M4aqi/1+5Fivy8yCf3PmIjPmkvRTX/QwHy361ejxaStkCKqopqr3o3dfav/Jd5jNd36RdN4r
AR0eO5UDCf6oWICEsZpGRJA7pmNp3S/GnrVXxBZqbizBpjcdKWR+dN0tZh59z+XFDepRupBIsr2Q
YpxzmweeHr6sTXnDJW0pN6p/Mbf8aFKQpt+aDPe34DXWi4xrT5zZ6APj6WSuK7pglQVgf2z30Ico
y7KpGT/cK/60775+7bVg09d21BOB7fQC0Qx/MRM0NRRROPurHDBwynBm7B/pzsuvx0wwicgBDH1T
98QVRtBlQQspJZyDYvsIPWmCji1J+Li0JKySWi6Vs2IR278aMHd5JiEiwuXnCcNWdJOGtDRrnkLp
aebj3w74ST0DRd9fP0KXnKBDa1XJj8+ABx1VJZFv/Po+8wXqxemM5D4NXR3Bglx9yQ2+RzKwY8/f
wjdnQSQmpY1zVYqe3xnXn+8DlVG8Z0mNFQEAYTQxKu3emiM+4KKqt2jevQqHOK3pVIOtOieSJc8I
QnSlHIK3khMZzjQ2XY0JF9G6cZDknOyq+LhVi3Tf2Nr/F806+l2ANLHfjNDxfLKkCavMANpN4F17
8hb1F/bstCqdjv6v5oZb4fm9zgKtkC8T4KDeGQdXE6hTj9+NLpiXEnKuy4pzRs/k9e6N6Vc52C/B
Vhf8XhyFAUossc180O4U/068Z5gng64bRspl3MfMEz2Vv9FLpGCDKc8UcV5xzcIVsDKSH7Aowjn2
cWXqMWb5tremKOI2Mobk84OpWJbeOi+80XwEmSwFgez1BFWaohV2vXWxaloPAkh25sq1Tkw/k1Tf
HOz92aoxawZo1XhcNFeSpm3JY749QRM2tfAFkpoUZNz0peHNh1e/lPAIuxnB3cqSqyK6c5oAXbGR
uZCRs+ssjXGUSWPy+RE8J/DCHuQckLKPOyHl4cI22qHL/PRbBfKsISYcoE1Ta73tOdHeILYgAMbf
tbX4157fyY8BcY3H9rpgEnEPD+gUgcmUpHXE+Hq34B17suTqP14UWL8k2d7mMsSSh3MgA3XmM3LE
EgXmEWgEE5iSnp8nOze/OpOq8xgKLn58tR8kopGRt/BLqFPwVdnrSj1GFPJDuF7zODSFJr3lbXui
PayBN7kc7ce0T+D+L3FBq5ZNtmUHHC8A/ASy+GnYawjjgnO81IknAg6oG1v5wuYpLBvfrVGn3YP4
K9A/4xMgEC27W5Hd+Kce6kY5BfgLzZ1LGUzA1g/5PpUIj7kfyj2vTOz+qescPEk7XcQMIxJPj9i+
RBLcrEtLBEiftVsHYaGKx0aabnv3hR4MOtbyD0mUZN5fgtc/b5IH+6Dc0zSwy5EcenEKwTZ7wr6h
JqSzr6IMFtlj4KSR/qQ2+3S6iBbYBwm2fcSzDaZNzyhQecXCiYDZsseZPPSFZNGWmp4jHdLdpXBR
iazAHl9+SI6FO9F/3CqEcpu6oJcr2gQ4AVTcy/KAB4EVjFYbmu3zmgi8Pr2acNSklXQ7YWAYQzjn
9oNXkPT70vwDl2ZIvoEeP4VaxPX6vvLnLk5tCHRMX3j8U2NkGBRT/5NO5oeitl6Iay1FG3d6BG1o
ldnVHpXj4rcnSOsiz54738rZbCaU05mRc12meCt3cP3w/SSkDNa04AWGa8JdzUpTblTRA5yJYj6+
DzaGyyz5XbmilM+a2QX8DtziI7UvYxx2dJSHbQqQx2AvSa/Y68WrehJGK4UTAkxH2Sm+a9pyPH1a
qnuTcSyu1KMKLXVZPJnp64/cvKsAM3RKwUaiAbe++zHrJvgTOFrHsGhhYUnS83/YYDxwqixcq/Ze
/ZfVsgLo00ml6C2BBKVLq59ASZYWMfHpzp4Ti38YzEr84sO5+O3xL4tcPXyAtWLL7IPSuRqUwpUF
+HGZXtAU0dnYGnQeO6X578ycAJRmKJI4VG+8GE9aW8/CFkfihPG25OpINa5aM9lAoBO0ryGO7H/0
kb3ERKZTkxEszWM2BvKxtjzpqgAC+0D0LQ7Y0eyOgsroS03ui/fhUjRglkie2RBikZo8o/GaHwIt
Q85iCwstMHL17opm4PDPazgfB6WbT7Xe0Hlc4C+wLM5h9qB1lS8Y9t2ySfgJD8Cgq4rSav1l8Q76
MVDbKqtQLJcQXERqu8xmP9LZbq2zy+heF8uZy5JJA+SZZFAD9gzpk4CN0SOD9dURoF3cOH4GF9+h
5m3X/bKocq3SGFDI2xlkOceXEXkL59Ugs+D/hjPr7L0ZOeKWiQEb5EMjEafh5s5Dk22wAwgEjNhN
qnkR/PjX2zjZtE77MzEwx8caaAwimVAVxnHOs+GW8n8nzPUorslt1iqsZ9p9j40kY+RCBE1uRmps
7eFUMIIDFaHxzmY9cPxGnnEDJlTbdRL9TgyNT7beONmWksTX8Tvhsqn2eBMfhCRpuGLD38JxQ7lL
f9fM6b/cG5srwicOqePgo8dX5qvH47Qt/1Fc5Sf60rpfkJe8WEpUJ3YhtOT3DcGTvUVwD6t2xf9P
3WZmqkRHLJFWIbExPyEt4Ib+LL40uAeBAuix6RzRhoNQ36K+IUGlHUGFWrJLJvclihm3fA8EQMpa
5VvBiC0dEdf7KsbjZxKj0xRcOVoEl6Rw1jN+dFaT8hgA8jFQUld64RD6SejVsLvHNbvsQwO1nBGt
hyM2YQpMXTTgtMsVSIr2FtiumaxLX2Nit36GcNMDBcuvPpGc9gxMSFW2jpod667P2E98g0GZ47wb
2Ebj/Q2zw6vaYoQvBISGEswBw5fC6VnsCoPSBnfTr+ZNZpJh/S0QGSPlbkjge92hdkFroAWk2N3n
/QikVxQhUOlSI7PgnTO/TtnvJTzIhOINdf3da0MNSyuQkpbhhEO8ApRAKcdzANhJRvAxT5kDs6zK
qVwfQDRnl4FX5roqNPFRfNqy2SSqyaCDkl6bdIhDMsoFxIeah74hppuVXyLL66xEuutLsN3KQL5p
lMvSVwhdCeOKTYB1dNNC9WW7foEUDo57CR3pPIEYDY+mfyU4q8MKqU+Wn5St9Ok6IqNkKZalu6tE
ihdwHzgJodNS96eBOpeIxhdMG8aGaxYSeYWPNlvHa4u5CSHKGBmZcwXrRlleM8cNlL7ZV5nSnVS7
xe+QlK3SezzuC67b3fMk1R99jqntXHkE9WThpOebDqrg/b283c5KSllrYSoFeWGBgbev2OAV8bEf
K3s9Bom89J8Q+482dz45e2byVt/mHPHUpprniZ8RIOFsFgCgLD0V7gKqKE9N45L3Rh1mkMsNLjFe
xOSfDFfNOLR3aXgYkCUU1lbHk/1SNHfyyoad8yi4w3HV9Rhk0/D36HfAQxysadD49pDqaWmIoTtJ
HTpx6rRQqnu4/M4lSTbPngnJuJ6CFytlUWwUdsPJlu1G5VsOySR7IUCVtZFBC2nZ6cRMGUVD3Vo0
05qOt83ecnvpmxuNgzLnTwo0IIKsGayClgm9yXKGy2H0k2P9D6ctr0sMejNzeNnH0gYR42LTHg2Y
JrjfEh7fFsgPC2ETB+lbpKoMPnHSL0TwvPh0HbBTYoyP5XTTqJ8NEqXClCU34ojtoDnBJnVTCqSk
oIp0UyIzq7kASJ17kYwFmjs2IPDWYs5e+O3Mf/65QFC0XbkmGejfiMLL1Q7NZYznX6DKwmTGWEul
++UA71GV6nu88Ry0iO2MNQzrNq+ro45v+jrzCmL2AA0Kl4wf7LwKW9M9D8+LNfcVwk1rcHUfaZLz
magd+20OoHKJUuLC2CebvLCLrkLbaHU532Cabj8IQegfyP4J5Wf/I32lqmQgG4If2n4rgEcMHzki
iMzOX3SUqkZW9KaU76yZVoGrlx0kz7OysYK5Bfjeuom/7ViGqd5cjYUceC0VyyTyEGIpGRhB3UWJ
zP7m9mylljAljlB8ZTKexJIOVMwg9FyCrLgYncHRXgV6KEKqcvUTUUSKDDhwt49M2In+2WQiPoqn
jI8SvIUVbSm6s5vmo5DwyhCPtR3pPw8iMYjEBhAqbVI+appNc1snkVDdoUAvOfqm4Liyx1QpUBzn
fQ8wmYqF4qs+gyzuwupFuDFC0nH/u7nRm9gV5kALBXC3mADId7rDWrlO4iWhfdAde0LptnZoH4uD
dkEIjIjk2EKzVbJtD2nqaTs+2KdI0EUoQoZtIyYSvrFETudBx+x3buPBunvkNpF79q+Y0S/jRAT5
Bz+ZRSPN99U00EjeGevq4zmHkeis5DezQ93hJvQtdmBvGjUhPCrTFwEt78h9ovjzsFfkKyM8HzYx
qyxYFMrjGgGniHsJ2cpQSA46mfH2kb2vwVZeYEM5hlzQO+HNlG7xpnFdOxFLwB5d8NH8vjCE2G+q
oeWmZjpj1s1BJh04oWEpZljGqpc6jUT3BzsS3IPIZ84R3+rY+Wxrlg++fLasjCwCBoK2wh3/m6uo
vRLXDnwabAyOX3CZuOTGA6DJma8qJs05aBgcIpp04rKG49BF9UvD59bcxCTE60LQ2sx8OAyvP7m+
D95qjzNoshBSCv0Kv4kxVtsREd49oyYrdqfEBNoCZ7wAN0XwUAin94sNJKDWiyvlU9d8rs9kuqJq
kkXxh3sxPIqPj3fES1a2wXDoCEaJPiCUqpaT1zsFbNcXcrFD9SizmgGchkoSmJeGGymbeBtO0+yE
Mmtn7Hw7Tsa+KzH3/Vq9ZL+vNbMmRnlSS4phN2UJgnWfZO9314k6HYYU10bPkOfCLfDLta1J1l7I
7Na4sYbz2doghYob4LKNF4oPcx1Vr0JJcFyABGIT2qBVyT0t156EIdDpyyI5Voe99qFzlNme03Tx
vTajLucT8WcQnnp6WsuXQNdA+mH9N6Foau8pNtWgowH8SfgcnftGBcuceAk2v/uLmm95GVMgj33+
A9iQE0+Ltov7F8rH5sCh5aquovEhjuKFJdykZEAs26XPeK7XNriEeaSUoUtOhvcUtOACUOETbtpu
qgWZ+6q1NMFDXNFe9d2+obrHlV+HU2ic2fJwW8H/I1TjcN7yrj5R8Jfnz8ohcEF91FHy0dsQ8kYy
PS6nylcsULkRzjuEIIgxLvoI+YWY0Z4AJ7PphAZERQncRv+WUNDPLVexqo8bP/A+k+kelvmz+a92
yv7kgseLmU1EN5N3AOwC/E8Ney0/NoKQoFc6Xr9w4xI5hAS2Rvu7NVfkbMf8wLvNXbEU5fO16QHp
pm8jw51rhfVXdti8O5j32aC7dVL89930BguW9OkJd3fOyPicwDH+URm3IIgWbW/+xXEPu0503jWF
L0qPWd9QKglRqY4kYiliki8J7NN6J0BOBPCibCmCNkevQ0CJAWbUxDUwR/bBYiwH0xbOfbWFWGuS
cMjUg6D9shc7mUkLHEG42KQ+PFO0hDlSNnI9vY515C5O23j88B16ov+5tMWo5JSIJKGCDaPRbl2w
O9fpq+X2OazT3VP6AeJblpM2kJpnreVpCwIvbADCjenSbgxRwc9+kDrvkwb0yvZiumZcyBwX/baJ
d9jOvqjwYmyAhrM8YpyShQJVzl0UpTsm+4G1J9QkJES2x6YYrukVMK6xMiBr0h1TUnE41scNDzUj
heWorzeVqKy58dcUPMpMEVT2feedWiFQZW3hk8k+Xkmg9T9ewOd5+VqvgeatZ0iwKFXt4xgcUuXD
mEn4gCkw1I1uo+wUGDINCflMVI5ALlbzeAubRkazBoz3c74q/Al5Co6/FVjndEJ09sGrkG0B0xAP
6WrC8000wayP3BOlVDIksbS8nSiHKbZWVjMeUx51FRsE+ln3dK4mEUKElVPs/Qbykwzw0K3K0/7f
d4rTXmSAucYX907ZA+fS/3Buy/r8mZm2asi9zSfQAsq2wOpCc1ZrP+Hg+nQAmgWeKwFxbel2LtwE
lT2zvvLDKsPMSYTkKq7tvFzYSp09+ZuO1dRnVxiIh9iro53iSh2JgIslN02Y9kMIMNABwV4J3fs+
hTofuI7cJbWG4uaiPCMC8+PA0Dm7QHZwYoRhoATnZgpgc/cN9LLKejnt6A0sGrNMZxHqGF2Qw+LZ
jvjByjxVl9HCWTKnJszSYNoHY6IJ093Ulb7TcnHgCzG5YofLfPELqLvXYrQ+J9LlLmJmPwYSfNN4
xVaffUKFC03Puuj7J5XJCK4+vvyZyfFLm4Kxxru6afZlQ26mkeXH+0dTcDzqkhCNMQ526d2MTJ2t
iJEyisiZ12kfIE5ML3LiqIf02ov5IeeDy42vJ/pdSeOE5R7PM9SmBbZeSeg1DiSW6KuCxWaiqEJL
K3xGntRjlIav+aQhtVMgHFDYVMwQVcJhmCcYooszvbYaZIb9PXCjZ/4i+BPi+yhjnEV5/cz3P7Bb
gfFn6rwKugQJTvjZKr3f2GGT903bYbLUmruHDT+A+NNcbDHT3sE6W7B/uDarDn06YGZomDwdyb1O
6RFpvzhgzmBjlvgFkt0qjodx7C24XrzZIqwUhTlyPNQjjjK/PXMQg7Dta1Ye1VUmwj/UY7m5SZqi
1VTyamb49BdjIFgRBxC4DDw+vqqTGBRoZ1lmoHnLtv99nAW9qKvakCYddKFG9G0/XwouRqZ7g9d7
2Wp0i7XTYEO2dtMsdxtDjM2qWYzGGllQahjeMWRInxLyslqmoKVAcDZwA7xINnsQUegKjsmW9RgF
1vAUJ6RUSydoeSL8EperLUzeQP++Kf4YacxiRd0VDZdZmzjr5DDK+p4wVge8evb3VdCEnkfWOZHd
lQxO85CVLR1IxmmdW7dPtJQkZTv5Q3cR7Wn+MaJHTAoqEYnZ15PSrXESxMyIsh6hNVe2YVVN5gLr
x1Eufzo14LHudcpRNYsrOwnZZecM1McC6oYM6+LS/fhM4nqLNFTVErmBwXmrh+WaXg6bRqv1bvPu
94+f+UD22PPfIGdB3FgIES7JD/Me+F2ski+a/vkFjvGNa1Ev+tEHRlTIIF5XBYRJcl3CR5elBgdT
xRDo/FjAvUHEZkQOUIVLa6n0dBUDw+MEaGP2Obaqzb0aGdE0bsI8RJQHGElmUa6lGjMu1rm7NZtY
0dZuFaDTerJM9kYIqSP6NPl3ZpYHFG2TQTW4YUZp5MeLy1CevX52+2T+a7CTcHM3UTfDY3vMjQvK
inqW6MfYXeDMIov/rI/5CeXKorAWKat1WLHaFvhJnGiLrS3U6Mw8ZYk5hwyQHmk1vpnno8gikeos
YH0nTku/dw9Fj1qwTc/ec4+kYFnBJH5ALJPO+xJL/0kTaJZlLQybeJyhauIDI+qC7DiEBrhQUP6Z
qUmk+s997jIZBRu8wyER8dghJydSGD96PwszsmFKIZuLcnDA0qaJ6SA+4LWFuCqUlIJ/NHb50sXx
Aizcq/e1U2BKGkD2HbJ4sWRJUMCw3UK4Ij83igdEh/PdCxP0k5anpPBHVQ9ihctzlJbpYhLfueF/
IuVJe4Ih6R44faFWluw8u5iJfhzHdW9e2iG610QBp62IiMc+/nqWGX2O4hKX3YBSPNKzDuB7lTnj
EFzulLlWrQxlQeSGHXAaZqmzFS543f3la9WiEHJ3ac6e1JnRsqZahaKZ6giCkXrn/dIvc9Lb0GX8
KsyHu1GIHvBLy2/n34N6rBRMA11SRgiuG0rwQXbJd4XSm/gFMyAeaccA6SEdMQp0Ri0IG9/hqSR5
fKvp3rjzy0xuBI22SZetaTvj44SUh8NQXlcAQCkYAjKCgt5aQSXrxz6xfsXpOj/HdzRJ8iwdEAOU
faVJ6++jS5ROGDomtMUJN+/jSb2nxGmKikXOHXEJW3rsi7idUgffvmF0K3wbggmK3t5QTv65juq5
W/qv63vmnQPAsOxd7t7CcdGBA30BML4556UklxbnlKNebVD1sOysGMGQ3PufF5Xriapcm0RcfpOR
QkIRl+hU1S8tWX/wOwTKN8cwYzjeILaoQWo8TFNO8RypsUKbZQ75wrrLV/PFwig6vSqk1F3wH85y
CJzVt9drySgTSZ+vykYhd6GwgAcvSEmJfdHI8I7BhuL5fP6C5gv1bFuHPEVP6nfCNYjJnCneXImR
ExkhiFXZm2FCJ+dRbomxMBcGCk4DQPbVSyIA+XZmgnMFt7FWajsnI3Tr8Q6O0wcE0Y7Ly32/+0/o
xVVkv+rBZ+u0fUoid6+cGyMG0fwmPVW5c7wImxeB2k4z340Epw3ekI+7hT4y2bWxvyRXOpHyYO2W
qAzpisouGQhs10W4KQLG0RKeIwdmfVP4ShtumzENq3F2xMywEMOJUX30voaGEnvXcd7vmIW1g9g7
A4Jh4uMhbiJaGeLGU8fRcd43FDasVBVZE/cM/xwWv9PvwwwXLUL1JhaRkSl+4dfrhbE2HGmuiTUW
wxT7I8ZAmE9wI6abSe3Ywt6zTqPFyLLxez6zc0tT3ZldIThLaJXgoD5e/FurYcxWyNb7GCc2kv1Z
c68QAgQ7XSDwvhWpDG1+2ugPglJKJC6IjWiEjd8jUwn0RCrNBD7eqHVEcBQ7Pb2zm0pRRzhlQMKG
z6UQHTdTgK7UWwtlQ0bWmmqiO220g3vGbtJXAHL6mi07s7Q8NbIqQzIOnzEUQRMqThX9AFayY29K
GXD9RP2yZ1yTPaNHZsLeO6HRn22GmtA0BHqpoFviUAF8BOcC8mAFIFdLvoZnJiBbTC2eWKY7xNz4
cwDV5E6EWaCQo4DX+OqGoG2R3SqbmfQoTsB/D/c+etA7EYT0/TS+NBejV5k7zagbnbaGVnVzSUyv
O7BxQguKowxo8zRyAuxlNbD1hlWpqEwc2m2omB1/qpHqF9abDxLUoKjec1lbTi+irK9FxG96pMn6
dedoae6cZZNFO9MwRr8E4uxHyJktEa4LuyUiG1m7ZJrOy80dtJPhthqmhDEJN43gn+lqxYkMFcP1
e7LKtZeUFeAoeLjkt+ZftV2crBaF/eM2RciXP6Gq42WQ3OCnWAc5Q3BO/BjlYUzv4GWzs3BenHPg
qHTY5AdXdpyCKjawaQH6IBHZsZH/jIHo3+i2baHXI6IAib2tbtlEtsGu1M4IoCZwRrYFYs/MysIe
opKbIBIwLIKDw8rr6tSIL7oQWmLgATZh8PkF3ytumKZr68t0CcmkSNO0Mwo+Zl4ZTMmHnpDNaXOv
Hkj1D7aqgB2TL5WtGmkKmfrAMipWpoYxnwlYGxEWLaqQ2dCGpYDo4AVkbKVsZqHxBwhigOwv5T0s
BDPP3rIHz3knRo7HI2FOxmsm629YJBRK9evrpmmgCvr7NzDTNtvQehHV/6Yb4o+6DG+p5oCyD3BN
LFCY+beRPx9Z5tjMgAz669B9o6u9Hga3mNkTJ9ivRWwYNWElLp5Nrd9Nt3lSVAOK56gdZ9C9j0Wg
HM5X2Lz9/sTdvQTvecBVHIF04aqMg1Vb/iyaEbusgAA1blowxHIFhjuzlE3UBc+/S/uDRN4rFjfk
ZdLbRCCPhpHLdgKxOs4crk0S+8+nsvWNSDPISL/ZX84+pc7OTFfG081kb5ZGdez+KLBHfS29hmgY
pF6EhOsudd1LXVF2gb7z/190G/8kTYJn7BaLkBMeQISryexzeNhzmhqOWdmrUdN8EfTNrWCSgwX3
aa9rebT1KuJ2FTqIhukEAWSTU60iyaX/CyBeQEUpcBgZDT9+tJmDC/SrbzO/G2RnHc1YxgsSuVv3
dwi7DaTVeJwtH/nSZBAjEW4EpSl8j0y/bxCbMwQpj58uRJZJ+G2e7TwukGawOEWCdowldboWB3Qo
oo35BuGnfd7k+PUgXRTcO1MqJ8Rc3Opr3VfFI6OZKeCJepDPNPy3ArLXFPUnUkwY13wC+kpkv+ca
31vedIzjwUPkac/J4/JSE8dfEyg4zIfsO/q1TOj66NKMai3hv6LXaxVlaSdUJSdoecyZzu7CsbRj
CL+lFz1K3g8sGob2Hktny4cFMnUFWDEg7EsKGEIZ/QdorsB4sMGEmdEf8MR2H47RDaOpIGyDI6M3
3GGyV1kKmAs6Cm98yF7AZwBZfaypW7lBXiKe150c7C8x55gtL9FpqtVKKMkEhVFvgCutGLm1qG6k
82fGqiST08F6ZyYb9SRgnW1o/5ggiuywHQsSeD/+tCKfiIMxTSA5U+r6HSo//O/zDOI5NlUE/m7n
xtTF+0VhYg55X6DnkaDX6KZeXKW5jMsCVf+HMMDJo2Unfs6H7Ft5XflPdLR51Au++ap0qIIp1LYE
3wZKw1eJf6LcfnAP/+nLaW7iuZSx8ZcxNxNf1Y8D2XH1YZhAplOF4Le1iq9MGVIfxQX2QFhwWFkM
wISycPcGOjBlowhhdLLN6KWhf72OKIivbRRIQ6nLegtAUqo9VC7zxwZY7F/iAgeiZmUX5iBr7PiH
yMTNJ09agpTCR77qiaMhr089l2fEBjzTTfCwVzI30TH5Mve1ulN3wo1LqL5Qc7GAeVfGUwQxCess
AOGEF8vVyafmiPneSu1Toj/2wDRo8IzZ2PL+npmR6mhsm1LnRFM5E6+ImuBeBIYONwrdzWNFub8V
I3lD18+0M7kTxldQMd1vSZHYzG3Q+MEMr0E4eaicO1CoHWPx1hhobpgRju92lAanDbhQ37oBTg6Z
dyCWlx7IrRXw7s6uPd5NmJyBWw6Vcbsxy9lMi2nh7r8YU5NOv9d0aGiO9s+A8cv8xFZsMYEGZyYo
cuQOi80f3lDzBxRV2HkcSyqfzswbqRf64Eh4NyakfznseDeO0eH6G72TBBV6fAfSGuU63hZcuaGJ
aeDMh5FDOCU54WwRv840fkpmkta2Rp79OAlajo3DdbEF75cAZyaBO7gLvg7eO+2WzP5DkW/sRBmW
4BRf1dDyPOnCLBU2XblJTz18kuB7WHzoZaf/u+D6Otq0oOHY6tbLngFQHsupIg2suFdKJjSZp7W0
6Gbx79XpYA9EYk0sJNGjf8OugzYn+GD8tE0o4iYYgFbbHNmQGxXGnHumKetnBUREQGyYQM12aZO8
/ziFpSjJBx3ghAIkrn/hIjMDsl1nzNBarQAlwONQzD9SnlSzmtiTX6WCv0U0uwij4ar6TC1xghuF
VvGTxWw6HNIjHzqHr3niGZgnvo8BnDsZqSrnScGZNJulAwyYwTdEth8cP05/EW60avFm5ruTLguP
FHv+T+/u2Djjt8iHBfXwr69WBKqaP+mjgpBi/MYvCtdCJCJgbx0y9bwHLEEUpPhknBRNgaHNC1Q/
xp3ijMzgKRSOs2UB8v03VJbywvBb6Uj+f2+B0h/L82kJi18CZnOZ493oJCpza8h6JGJgjqQOIZ60
sQsi5R2r7ka44lP60VYJwUo8L5robDfZk1MsuYngkGdpgYg9Idf094LtcZUryjLph1RHHs5GBIRt
VYHxwuRefU7tU63Tn03gwNw3Y36Gj3/ONaU/YhTnlHjzfcHm0NFizcr+xwAhmKuJd4rhsa8Cg00+
/xuJE7czfMrJvABZWsQkd58PTVBnIdIPIPh4YjGp/c+bVoHoY7VJWYGmC0BBqvDOS0dUBFhKBiHx
EO6ZiJpLSdz6xluXQlIfYPSxoKOVUmd9j8NISLcpx2FzlKzSDxLaSlaW5XhBErNWddB8W7Kc8qz0
zqOdRRPgyhGG7tcguNKe76zlgqF8UJmgIZdDWGuWpnR8MDe0qnIUDbUE5IG2LCivyV+axDBev5HH
n0MmzbJpfXF5zedWqOEXcKavBXTy1W9h7zX2qx90lWR/2CDTH3IFRAFmIEmqGLNpxgJBZd6pQPlw
PC3ttsDPUyAqssDRFYLL61p3mnBiGX5T1qFenTWKNi+ZVHmz/MkaYU7FcOZaSEenCxgOAtRF+CzQ
9G7nNTAvZqdP2WQVPsMXzPi15C6WOjhFfPhzDo0ybS20JGLRKwolddYjn9R5s3SZ4xojNlYvn5yZ
xaC0Eqv5XQO9ayib3BbydWZlcpz2jJ1scYD0ZEac3sLrEL1wgWSJGv9Sy6TICXu6tJTwX+/BahR9
E68ti2SLGSb+cLyzYGXtGl6wCDS+talBRysIvNHT2+zmzkDl2wjnFmoOyHGtlwCPKcyxDiqhRPlQ
506dsuY0cFMolr5QHraNrglVwbc3ijBtvdrGn9spbq+sjgLNyftImlAxjWJ945ZBF7QNHI6d0dqW
76b2ZCTdoBvkrzCuoijUMbRf1jZZkNVMVuL6x7+ZRHEJtEtlkdclcx93rTWCUwGIyyQVSJOyepV8
yS8yIvrdpX4oY1hYgT5px6cC1NlupA7/cLl2KqdAB8+fXsxjiphT2ETQC65PVocF8wm7+ubuar11
vz6m/X2k1E4mCOx6jVYAd+bclFXlnhihdSar5mrHNs1pXOrbgysdwcq1jujqHOiadTZga/qWtAYQ
wekLHMRL1ivzCIWslRnCofkm7e6anxstSN6zlv4wna62xqOW0+QJ/9B3CsxkQq1ucJY3QQjBl46f
yic+9loh6QYpWc/jC2oy4tNq/qC8LtbdGnW8PctnExEbVVV/9iGxiOxkwAu/g6NAZIausrKO/vMG
28400H4kcGm3mPUySqP8kAeWV9GLYXsxy9WnKBtGlgRmsnHZmCoUvLVRswtQsLlJ/ylpzNBZqtWB
MM8NfbE+oTkxW6JoSXwfclkGDPk1nmTG1oRaIeG+0IO0+KbESS1gWPL8pdAAwDD5mrSF6V+nzZkh
XkPclvaA6UT+DMT31fSv7CfzIL29TZ83xZoO0dNglwcI+7QwvCy5B2NAWG2kCcu7LmCXhg+ZQmPv
mKgwWVAa4Jvgu6RoETa/f9nuC5z40RH7t7Z9aOI63btAEPf4XinYg77cfQf/8EK1VStrHRfphgck
kiv5P6JfeigxrwpfymlGPk3xA1YReXRpp8RjIUehUYdsF8MejbMt8KAbcE8vKWhiHit/ydWFI44n
z6pNpvT5PU08vQVjqOOt55IQslP0OfKW43Nwv9/bhzdbiPlnZrbb3PQWxVvUh9HBJBiY0tOHxDKG
K3vpjsj9Ya4YV5u6vrVvOJITdiE6J86LJAdk29CdEMx7uiPgDF/xDz3J1TB54nb3cDlU9LP/BoPS
oDeJ6O0h3/ksE7MvafA3jMDoGX5pioeTS9aQ4E9cW5+WfcOhsxg/ShvvUtQSh2iaN+nzw+OZcPR9
YC4fdvNRC4Fut0P5rwb2cFU7IOZSbrhgE9cJHv2tEP5ns+LqXoKH/kL4N39lhJNrrsjvkxRTtcmq
hBqfxVzvOVEaXjSoQzIAlDBhtVyNa4C00j0Mqlp9PTX0mxxuqNpd4kXFq2KJSCj+snQZCgTAelPl
vi1b7yq3Ld0IJDlRZozwtBzoOht8nY8n5J2ggC8o5h50tOgSdEqwlERULYDYEogJPztZG6HMZUcI
YWwiT8pYLq9hARQ5V+M+rNFlpam02q9UWN6R706iojLlDoe8YuLELnydkySB76n/5S7M8gKjfeAz
OULeFmeCLJOxQkSvLAorz9rRV6L4eYkE27Fe7iPnRa6BpK1eCJgnek/1oQSIxw2tZsZVbRWwts3S
H6a8WOxNyJF6rciDf9E4SUPx7uhJqiEVoPxr10D94C4hYiNhd9HeHajOWm+rRdUTyaDsQgsf98Rv
dMAlLS37FTP9QrEc3Z2TLLpar9Ml68zqdWj2p3P+IqeGUlzo1LIyBrha6kxzShgG3CAYLvtu0Kml
hwkv8sVNazgdo9wZYuSnCrtME2kI0LG4gJ1mMOON3ugv/U4ioXH5734mMNoC86c6VUllEV5GokCl
hQJaxa1zlJp2yE43k4Y9bfjXRIZwagbyctXiZgYCuZZIRrSfm6ry8u/lURz+l5aEU1iuI/SOAl8I
G9q4pJaKM0li7WJaWu+7ZMuBgKTVDRhdF98YnE+7swFWs5Z6VWa1XPtz8YrRj/OecJl4sWmRyhIX
yYhgNW9kXJ2ZdrZb14XexDrXH1yT/C6twi90QnU11s9j7jzXgdPs2Mg00y6updQlssN9ObfvWriw
tMpZi0vW2wdu/daAS1y1+u0sAFB2JtP87yfr7o/+GlHKU9cG8NHBEFZvz6rP/2vr6NLL9Gj/ZPAt
CpKqFwTKjoce6L1b5qDb6dshOaFZ9hYJVdA0VfTdxIF/F2DWBFpTiFdaXJ4d4RaZfAFSIoZ7BcNP
heL+QLBl8AU5o922YYGIcHhPZ2FcNELrdCu7DnSUWY5fK+mF5zZXGQ0q1wc9hS1mAt67NBKHyyhy
Fi57OrFGoYDZncryWxb2p099N2Yy03HxJKrt+AenT/vzDq0F17Rxo/2Vt8QX0OmwrGqf3E0qMVWX
08FjXgHZSrQ43yhzDUoSxhs+TQIiBaFIqmCmguQ/rtfT79MOwCkhxgXDJ4KOrDAUtBOHQLJ25hR5
0dZuyIe+eOBKD+D8GGcg506DAk1OLKXIJdjTyFIkNfZAuLME60SI3ADoQR2kgMeR0CbpwKP4MWoi
0M6gykJYQZVb0dWSWSq1vF9DKvmVpu+JWulXUtX/Jd4Op6xtKFapwPpB96PHRMe2QZ0ybSwDiASd
7iMmjs1GepKfX3//gj1UWda25yCOYnlaRdccNuDyPYOFbfNgjKinEbD2GZIu0GAJ/Fuvwj1x/24A
LG9hBzG4CdZ7H/575KEmvu3x3715naMVf5X/L7e2BYCuknGZvtc5B3ODxYdjpgzgByBQk5L0cBq+
B9XhgSVdPg6Gdb6FTCJeDQw2RQzjgIn31dPXh2DictxBYaEXRV9wgTSjhkQpUEa+B7Duiq6Eqrsg
4AwcZlKMowmgJ+jjSr6uzXyvA9UZggLqUL+JdcgFCGMTA7tm1+mMqGUEhProLPesDYRdFXF2caew
IoRHria9YvTSKnOBQ4QRyMAycYnPkhiiZrQxcgVDGk66ljKzp82KfmQycu4iA28Y0vc0WddAPgEU
R0GY7kVWStxreLDUOYrwfhDP9zWnBQn/i4MlNl0HVSNKKvqpBaNLjfU94Jx1upanuiDY4oBSYquL
7/vM+xPTJ8TiJoLo+HzPibm1HNoCwWlqc8ZH6uwC3t3qKw9OWfWXBcg+BIB+kCa4JWNWEXH5IZW7
KfyujXdkLwRV2iNrkV9mYmS6iRrdf/4oJweuUaNHYp6ca+z7n+LHyyBN5W7Jc4YS0f2KlZjUit5h
Tvsq8FXEFbaiUac/J+Ifak+1bxaAQ575jX+Qnq+LQvO82P3fxBa6KZ7uwpwcQ5UBgjRB3VB+r6IR
LOr38VK6N0pY8be9PUzm9OBpPIexh3KOs6LeSHPxWo0MCXxt/g5sBbPXyzOIWPO2UvFmHBQ9JxYH
9wD9hh4oV/miZLxjL41/0NbONO12TACBTs6mtRQGkaVOiAGHGs1dUa7Ow+5XGTD1Uuhm7qF7NjPt
N8M56i9tTXpRElw8EQY67T/XtgqmP9swza4Ay4NQcu0eZW0J5Gz+gMwZdfPsl0uI297FUQMzOBBW
UOncq+KEXmoHkeDFkTB51Otfva8+LlzIriXfYT3Uy9ucn16eM0WRJZFgG20HGdimXkGIWCrhKddm
/mp6AdqO6rx3A33XMUAobkfdrd9FB2gVKt5QA6hAoHli+TnW0X8SR6t1kCYJRlEFdrl4BlbXEKVy
thzdw4d6cTnPWtu5JSPT5gyaZehnAK9emjodAx6oZO//uNIBu5RrgbFzoramDpcGWZaNCQLBPgx5
LQON+95LypPCuxkXXYzpbs7Y66tDPS8xEUFF7QFomzLW0manIK+mevjKJ5BjXHWYB4qmXdG1WNAO
U3SBnyPYx+jQ34wJ3Rnq2C0ED+ldHjGYd1JuX2iRiZteVIa22gRtjTbDysW85yxNi/jp7LS0WQX+
bt5hX2SlzhN8knIvC/WrMsNdsqCbj7l7z0n9IfdYXeRATDQlRGFwpo13ysJXEXp2FaJe35oxDBoF
nwi/4B6Nlpxz6t/typLGnQNWNZ5CBOR7UCkIShqwisTD8+INMK0kcE2uWce8JwrIQ71Qpz/6kHbb
hoCqWF8CWd2+3iveODFrVaA9zqBZJ0rzOxpl3kEzb4aNZHEvXL42+3RI2mLaMJL1pdum8R7w/xTd
TugPu8CSIsts38I406aIqZLDb9EFmULr+eoCQbXDDDk+kRivq60VxzJGk3xNrsHD+NHjb9HsxcjM
gr0yelKO0QrhW0N9ZH1ZKYIO85mn1KY5+/xxlIB8OdCkIbYp9Yu8LmPLocR8ZuPZNtMkfY+XXOwi
ia6/NwaMnWdgCHReE4mvabYzvlh1VMi45YygexMZrKRHXo6HzmPDLKJvXXNFH53KOimPKRM6Ar2w
jYmzZoOd7Jcex33JyZuU63AQmywuOrlbR5iWNXdYZjgHwQIVux7xCO4asf/0xPHbod4mvz4/7pa/
Z58PGf4JafIJ080ipEV0nJEwIJa8gQMoxKREE4Bwb2yXaArKg6npHaEhWdS9iH+vXtqePtg5yyjs
mkOvvkmaN967y+wblYMWhO54h/h40NnyBT+tucmE4+/Ak4GLz2jkIYuE0t3EsODDObb4tUIt08sT
eJuYjikk/RqXxubDDrifcIu7zo/I+gzV7OhqxE9LKWQreV1oGZ6h5omYP69QE03ZwHtXEC0k3QtP
QuyVRQAwvHmYqMak7hKrihhegkCL0UXWJEXqig5ZEX1sQ+MRLH48RzObtBulwm/uozm/jEQy5nOU
vunx4cpORM6al37bp0nGt81yP1r+MuX6mfEUsMADrj+o+UQ40boG0qsVFXHB5ci9dLnw3d8Yc6hq
Qt6p6o6rrVsQEpCZi+G0j9yKm8bDn/N3f53s4tMaFYMz7wqrFb0T6Kx8P6uPrlj+WEIhBN+c9B36
gucQfOZf57sXoB0jqUoDx4HsXkDl5akpVZ+/Fgn0+j2sAuleb00t42Ro0tGhu5nyKOMuqGD+va1H
6BKerX2OXypGe5H+VS3+Hdvp885lh8T6ekW0MeB0sxhA8UZKe2eH3xW+bBhMKufb/z3vthULKUi5
UTFiIk4VuldnwIVEvjA3/IKV4RtHfDPqq0l4XmyCJ5peX8OIjkbITb5jF7nyNOzJt4JKsakLOEwO
s96Cu78L5ONm2zBI11lBD9Sw1BuG9Z/flocyqOBGVG+eUkwYEj3kzvxBtgMroilFS5bUyUtKRSn8
Qfe+Depzvf1Jho2TsgywbDXz/oSFa+jkUnW1isyVLePm/34jobdhEav7wzuIgzr0iJB2qKdAW3n7
KrsFd4ISkquBh+vh358Ik+zi2ZR/BiSydPvnm9dSm6+RaQlrlLSSSj5Yzf/nSbcMWfGW7KpAnxKT
JrNcuOW8SZUF1QP3boIoKvp40mBvvH1gM6Gf+xbLKMpIGwIUUaSKg/DtQ2QxIoLfWU+qRR/VUCS8
bs5YzaTyPaPpO0Hrzyz3YkYLhVzlFhgqBEKVX/wnpUDWsyvhK2E6pcOGdIJABnd/kwGc9s+LaTYE
/Fb9AJkQdqJCApj2Fodx3tnFTTkbUSWTMEQhw4nWChfL4K0mNG+YAuPyWpyta3AwACzIxMaXlUbM
4PJmanBC8PYTtezpcqxQeE6prG4mttQR4C8v1nZTxl3P9QehDpxbC6xxiF6lijXb3hMYkqmvplWF
nY0v9Adepdbm9WH27X5amh8cmOhVpnQkAN/nm5fTVS79BbZZwKjNeltx/jyTQuZEdz4dO1W38eAa
Zx0fDMMSekj5jcFViLMgFH4FRvae+S4COCDTFiJI8tvTP3pg/DPKtUoH/i+FyWa2ztx91eWWHVv3
SirvyRC6N7pl0eDkB/Ee17vat2AIgNGxYkB9DyfDSpizyQYNk25MWP2UfVbEsp0MpkMUgZfM0ov1
0x6KfLhp/Mbm5ParuR4xBWVX+dRMi5J1HHPTIs2AQBi1gRSR2WZfWtV1XBngyRiAdpDzZY4KmGaW
5Piy7BHrGB8O0usB80Onls7xabEZXcBTCqqoiplgu7GbiSn5FSFVvLS/klrvDraunLNo3C6Mo/Xn
L5iSPAXAhSzxMu9TUZS5xIoxVIQseAfQ5ChQaytyIRiMNgSL5PbnJWBzEgpekE8C8ldzimInHkza
D30y8mSgWWFLMJ1S+zKWIoTHy26tmgQ7vJoqEBjWNv+Blhfnj6IjjKxm4B7NABCW8c/lUGBPQl1x
bDUkYkrbyExDxBX6yfhcb9HeUxUVmQoogGmUhC+uI7vXDZqSKBpTVmRfxTK6oyFWxKNb1rZ0feXU
qGcjjF7N8PLrD7NnGPMTjvd4zmM3eaVims91TxpckVgjnGdSsXC0cDE2/LiA44IdUiBMp2LqVG81
jN2/dwnUtw7StQpMWAbiF5BgOy8v8xDq7PNQKxshvffQAOk2/0ysqVrY+vAZR5YknGA4jDKXeKJI
TqUQoCIgOQRF/F/mHrQjZAMOSelHYbUC1OhbAjH2CXelqiYSg9RotcKm474QdP/AnIwYkqQjZ0A/
aKuWU9lj2u5dcicSGp66jX9FFBcdOEwD9aSMT5s1yigLE1QVYuKm0GXui+22fqnUlzwao1fpzt8z
ffSEgYNQRLrGdIUUPiOsZ6UYCq/pGAltPK8qCjNUdFA9GRz/wF0LpeotTXD2gLlFW5h/e/f6Pz/r
BpwKISi0iDdAu9iUQpxu1pLxY9UGNJGOvhQaa3RkxODsD6v7bZT2EMyXJ+Kwb7LzS9VMNUGii5Og
X9eIrVGkiTCakbHIBUNW8zzBn67K5w/V7cEOcQG42OkiaGmdlvJye2IFBh+XN7dgW1J1rlAZ9Unh
Q/Z2qlP8MEOmbyg/yemqVMnaNTWqma2QURcNccrOQ4JXJFqPdr4SkdHT3sy3Crrw8MekpNFFi6WH
dCENMxFuLADq9JBUj/Coyb6ikdyt99d6y9VXyLcp/8tG/EPIfO4nNTvB+ac6tlt264YP4spWy/bC
m8PsacIonDtjveCFvkCeI+t12ewf+nrjCImMphTg8ne7bUbeaidgMI/f8RwSUjBW4eoUQi4+MAvE
9d8zLptfD+PuJx++G/QEd2WnVHL1sTwG/BlCWH88ukJlx8iRD9QhPaiWZvWznDzv7IYvZXSJzdOi
2dPE0FfQXDMXlM1jDyQAo40wkM8Q3NMx49d//phXchjbJm7gykHgGIT33uGlCm4BYzVKJ8fgmiPp
lVaTPbEtDBMy8Fw7eqjtBFf7aRAWxonLFxPj210BF+Tly2CZa8Qm00e07PMkb3Qn0wskFkVJhpld
3VDbXXrVmNKcr6/3GzBgc1zPovoCU96WD/sRvAMSsG7M5vuyEDcBoLt2uJ/Ao1M42ft4nAHsgE/z
uyrxL0l7QCE4gq3TWiGi6nrHDV/ZDW5n1/jF+vMXtdpSLbKyHc21p6rJyYfKz9zgbX9O/z1TKw+W
L4JX7/lTr02Xj/U+MQXk9Sq+MpiYG7DKcQ7NOUBx2X1JICJ2QXhOHKDiWqzrnaGHYquyN3oyeyjZ
dojnSiWOG3Y/Uo77Y0jLpxhW3fBfsuncLarVIeZMlmdi2R+ckRrUz8czESWjCZkcbuwRHNlgKqEN
/sB08tlxUZwMvTra7UsJwcMxv0Wj7zmIWWPG4OOtQzbsQOkvyDRke27vggsNirKfXkmmpnsQomLZ
Tti0mDR/xXAPq8UDRXZ21WvltMYoor0CDcoZFkhijhVly2NrTTp6sigmZFHa/TFPJ3v49l2D+lN4
qHe1BoikihLthrwg6hbOydVlBv7CWSqq6rTD3gq/7KEJQk8zfGmi/nzLe8egi+Nv9XFfwK+VCEjF
p1hajzTF/DQBj0B/pAdSDVzM93Wap8t4xy+Y+Mqy3JG2TkxqMXfHZXAvpsX7tmZ7BqkkXXqtE54p
MITUmoX9qzxgFjtbj4a8Dzjnrim0pQqvkXustXsRMSYvqhC7+jsC2q0+Ag1d82JxKlU3xfbe1Wuv
+PWq8jQj0hiuHzDggZm+oSyS6FubD4isPSDD7dL0SJ6G2ZAT+tZCBGVnVNsRjLKVzVk4E/ETTJKp
4Y8lwpXVLMhoThNBiJNsd95sOInx2RmpJMvA7AjM/5kRglSmenO+chCiQ6RpIMZgtHjzvsmCwBRQ
pKHWRoLbbZQ7A6hbOIlX0G+CjVjAJC5Q+02U8SEBXl2JcBoUa10AgAvlN1gu6pH27EhOI+hRhn+s
aHQfYg6sW2d82syB+S/HEp26FVEbMWgbLkyt5WlCruOIp6eIuClawxpefwjXEtKPVYyvSLIcEluN
x2r9NBu2nBjwE6Y86E0Rr+piBoUYehqGPWF9iIT2ZMVQZNP7W7MMRkBCAI08X5tL7Ffvl2VKBAkv
UKiuiUins2XAjQCPzknqv+Zrl0/n425YoqMGREGse0sPz/dsmePYzCQWwHOr5iXPpsbizJmYt2CZ
ZiOkFFdh2lhtC3iKudZmDe822ABYgg4aGet2h/ki6vYwbiKSjKbTilD/CgEMLHbuQEW9MWUNC3uK
ilDpQ8DzsH2HBcTPygi7Fll9rtcNQQVPRXqp+/gHnYefYodcoIY3aMiQ0V6LlDbcCZfRTksNS3sU
GsHZ19X+B2OsbYffpecgDGLxbS5XfOHGSjB8kbFIdTKks/3JXZL3f8MQL4XBgrmohgSezNcDeIIf
vYSRzjvwxqh309Vj/X17XMANCbyI542JXwej/b/gRQbpi8HOG0US8CN4A8fFd4UNcRLtc1/Bspos
BpAF37gUiz3QcmHNZeb9pwPB+1RyQwVUXTKEwo6LOhcYMn0AkyoLnIlXZ4Ito+v5P65mp6Mf4fhy
kvSNsAElUM2H0cQoVjpaHqJy8AAQwfJM0SI45xRaFqjt2U6a3Yte7ke+Gfp5DMrUG/TszvZg/HF7
IjGcqD5iy6JCYlsjngHGpfyEoGCpcJGSeMAG0CMiozeCFoZGBCAFf1BBwWhj6ShnLgHhLinjYyp9
JW/bsfM1wZ2W6x7JR0zTdwF1jGeajU1fzF1aEbCbK2AiVqJIAII3xLKQRYVLURh9NL6rp5aYEAxr
RMk0CBEwfIn9M4a8rQOEBMvIErYpwi7xNj1U9SlRRUA4BtIQVjogDvGO+2jrsZM1rhS9BXbmBmhf
qt5ifIXbUHyGJ8Xmeb2lxu2cYMM3glbwVtQmmwU5nSnfuFEovNCOM60wb5T+yV36OhaTLw5AuRS9
vn2e45g/ktGwjPNSSo3OctVjWgKaTSb4GkYuv2+BnPiAP9b7+z+TAKIU0sbzg1MqHQkW3wqqDfxN
l7hxJiNdOIrKnoaBLzwT6I1dDcA7DGV91wEbjo3zFT08+eqWghPyv21Y5CKak/p7wWI44hzYSixh
bgGOX0PuGUA9edcdV+cw3NtuETRYeNSwLbqASU38s6Eg9M0g/xcQCSEGQ1tXZuOZu159W3xAjOpP
kRURSmwK/DVaGqSA+cb9pE1M5PZfLxHdc+voCMjQ1TBqmOycxuQ+CwfrogHlzLOCp/q9VmKr7CIK
hw5bx53YncZpBaCyJaJqvWvCsFqOoAtPIXmbDoSNVFp6PqY8ylsqwL80OJSHCMnL6z239JlZtAhC
nhT/2ZQyj9JeBo3HYcp9VuSRYTcApW8XMViiJyLLPYsB5ib9bF0wLe425qsToOaKYwOK5PepusvK
M77f3XpTsnIx7w8fwDPYL93Iyzu7DkS6k6uUnomjpZG2V3kodH2ep9ZsSsM9ohwjVjJX52nRLVuX
H7ecZzQb+rpntG7k/whOr6tFY2c8CnDNeW7eQdCAfroQNWxhs3m0+X8xcGScjMkCtc39VdGJ/Pt1
ORzw9Vn/KZH2b7yz60YafI75m0jBEGYfwiy4PXlr3mJlWObMVAd/e5a+VJKIpt8DuZDgTQRzDNeT
+CirVX5O0VYV86wC49s0fn7HVnK/ByB43e/CC0AZfbAuqB+gzrjhtscI2mZ6yAj/F8LjqN2lNa+Y
mjVSLZlQ+sjxBPL5Y5YfhPHB6Ivl6s0CcBj9QxUp89d3IYJ6lcyY3bRwFOpm3DM93foPh+NBj2ok
MlqxpV2Ol5syB0V0eTCYOb3CWNuxPXzFtZxEVKjkTfCdXWrrVKEp2S8//AnMiOvwm8G0MWG3iHW/
y3wxjlEuwhT6NgxYtU+B2MrXc+HDIa571K/YiIAs+qCvAsgtVulVUwuOJaDwPy2SGzyfKilD9hmZ
oBp2Ivd32SPSWSgsjZok1VxK5mSnAaCV5K5TdZoBx/9NQLwbIwmTPJFWqH3PRPiaw2uizRxUU5RR
x7N0Tm2e3eOV4/96WoNhvR5jDSTyGUZB4mi5JNaWD5/c9Bz5cv4AkMubny58N6aoPLHxM5wu4n6h
E6cveBK63QbNyoGvdugc1Vv5bPtFb8pb0KEX7SDmhoN719Fz4DTy3BMBssKP00xgKHWgLad+SfhZ
8FXJulj6ntooUl1iTEhXFuTBDD4Hyea5giZR/tSOydjtvv73WeYLlgJtsO+abidno8RT1/QrvYp3
3LXeKZFa+U9yeqKnqOAprMmehi6JbBiCWIxJ0M3tZRoCzt/5GKkR18UCMCV+RVNXO+s6E5t3l/pl
EKYeebBvw6i0qNuQF4uh5i2xquyfLS9v0x9iSB5LcrE9FeZhraG/GaTLrFd+E3NbU3EYVTr/OKBg
xLVLNtRjohUdndDDuIgTV6yb4u9QzuHt523mPdV8Yq4Iro+RTW0uQcYP67jZ2hX4XBwmYjylLfAx
6owmtMk9kV2rDMUsDbP8i6NH9UdY0ThmhuYTq0HleKTz68IU7qIq5QTpCwVYz1Mt6n7RTrKDNsbw
Zh9Z4BKGeS5z3t1k5yf/kgBeDyTlK4JVJiE+vdN8jyB16vr0vOc0e3OIxyOn+P6H2N8UE3l49noY
WZyGfF3gGeAWVgDtsp1Oe+3HldgEeRfPG0F3vrGvkOLZTsnrgfkdCvzK6pPI4bsWsUXnjjw/wZdQ
tNpijqWKAmeRwdw6IPX0VFH22E/iPtpF+Ojhvmqp8kaf61jo5FHoZbZ3rXI5CVmCNVsQ2sxLDBx+
55MBdQp1Cwacp/b6kt87aP1D0+b8lEl6K49zxWyRAsasyxOB3n8nm+yVJ+NLi1rn+3T/89qGIbsm
GK/ggqLM4yqa1zRu2eb/NYEjdFZrwBWHXkrBJ6hNV7IVoW3MTkhLOVajGG4GknquyaakxvluqMLg
2Ml/GXPX7je/h6lofj9vhv1lFJcT93KgJvBTafGQjCk86a9ek3IdymBblc51Y9KamcNDM+XcLD3A
ifY+XJvtIhnAKLL9x7nzX3MwxJlZnv/rMquoX0uw8TDjjtvgJPLwQE21b9GEtKrBuqMgO1NAlUTJ
g4YaP65safhEIUhwL5MP2hIX32RDx3joVrySiWAEnzZvbZ9vkzf2KbgnpsXET0F2h72NY8QJu6+r
Ys7CDNunE/dCPZMn8RDcDhseybAOw/KXPHJda7MzuozvDPfhrRqlOV2ZJv6QUrkN853vZEt+Kk5E
zmGFZdW96tnrD6yZzFVJcBe237eBsgP0E5t2baPV0YJQMsNlOzn7kjXcwXvH2QSweruWGxwnqUU9
YyETIR9kknuSz0UvM8YeGqhm9MYlCa5Ozo9jH953FACPOx1FRxLFp1qePvMhmJBjSn6B7l8VUXRY
qy84pMao1+Au0jc+gPF9qvxgBXw1d/pwPg92ZEqu67DePeoz8YpE0lByzMxiBiP4RL6V1Cu2fPGb
2F21FBGQpOiD6PXebpYHxlKMFLNHwUmUKEUf1rZ35hOxgYTTGeHzYU/fnVMe8gjknKKij7wXSjQa
usXjtDvc9Mk08ccREGlMVyf6I5dRlrKAujzOVk94oy8YiR0Ad3CpLp6OlQt+eQDOy2Uv2N8OdaI2
rUVSoUNzeu4UBv0sjB4mZmK4seb4K1bqUkchR8MOCjGpuVqDDidz5T1jgeIZ2f8nxI/GzgcbBLmX
ZN5/XnDgiGqczM3v+iMHjp+I8Z4Thu2J5ZlgA3xgt+1qXNojRbOWwJhMCTTFWpc32xoKJGNuaIqc
sfoEDEKgBMemRu2+RjuFX3dtyjN3KUnUaeja3c/h4ZaWSe62mK2jXZwzecAG4VhlSbs7jKUfKZi5
6TBuU3ouCzTkMehMHKtLp+uI6WkG+xLmBeTwu7NM67IRZsKoqttwybvcSDHg1S/VSQrtmmD34Ejl
ltpWCxHZJf7CTGDYj9lToClIGZ3+0+5pwuKty1boV9DhCs4bs2rb2JUXHJIMGTluH8FCuDIJNjRS
Qw/EVSmA8Mg/4ekqneKDNDSdyTwjuEZvBc0KDNY8BcqKRGqIw/PwYEXAsRbjXe1AyizGgCDz1/WU
9O0S/92t/vmp/YIyB+Tch+YKUkANzdTmj4jE7q7l/e4ryj5ehm+lHg43nxzkkqmOxOPyQhdFUlCl
gTOArYNVXFgzEgrerSSdCj7HqqwmvaKBWApDsbQuMaGo+DVl46oFO5GHzQRGNvABAH7TGrnsEqBs
Kc3HR6cudGKAI0QyBN28su3M8QKr3GotqhcCqmrZpPGGdD8ohJsE/9Uc6SITQl1mfzrIHENPQZXx
COUUhTsqq48lY/q9MxSkHAQ/ABfA3xZYALB57BB6eNjKCPNqLoubbVJENh9yYKakt54N2VVTsuYB
2ltwkFFPeISO5ogy6UV2rmrRBXTSEIrN5sl3QAlj/LOtH2z0kyW2rnUTij6Xvtq5rb/i6Reqog6L
IgN/DZ1b2nBtSIpC2XU4TsOahuWwX5Cjph+lACmu4OUDbKRB/lG9BJLIDU2KHp0UhAN3lASMrxAf
CUJIY73hss/skaHqsCLgcJpYkpDVBowuBdFGEJjd3KTlhtYTjKb1axSdNW3olE9oQuoSbodwOf1H
nw4SyvAgEFm7ebWzoUfOhmrJqQOiE1xL5CnBHMc7/1jttif++/XNRHg5GllwkElKDec3vjFtyfB3
6oFwqnYw7/s14hlA0cQDitpDzYvStpPit2h3D+jKY8QHxDauSPP6PrkjE+Gfe5U5L0q1wzJLP/SF
e7IVSfF09A9FdHcdcnbLGt2RfhTMYEry4/Q0kb7Xrb1j305yw7pKrrdV1p7uTB83vH75U7Nk1iF7
LEzpzvGiYKMU8hGY99RH4pc8KBb8Ek5k0dC5pb4o+5cLkRxgtj52HnNA/mlecesQiFBeoyZaoQLl
0T5GM3PxnvBT/O8VeK6sd/zOG2NQwXraxr6q73jjfmP1BdLnCaTNsEJHgqBLk9aMgVhQo3O10pmq
tcyKVP9IhxYMDA+lq8DdU5cAu8BSQ/j8I5iVVPqPdtM9Uwchw5QllnOq754pHAJ5WeKilf7cdixG
jy1UPQUu5u2cN2tGastHVjP20JlHMHuJIqPzqeV2xNgPP5qZS1Ma0J2uaVY2pAaqZaOFhm1ycero
D/LM5t9nq4laGcHid3/rgIfmzAuuEmMsoRitowMdnkrBaQH6tbbn85sdp+s0uBjDfT1b5z7IVO21
9zIBEPi6Ggw9+Ase12xXL4AJnGHI1JZaePYuCxx03jLOYXGJ1gNwR3wJ98+bk06xSYhpXWRnfDhh
x6AtsIOwgoihVHjcBwx5aPWbLAlz76pglBvZelfUDKyqUQV1hDgOHRJkNbrOsJ93YfezccGqgQwG
k6TvOolQRUzR6MzI81uZ4+rdJyR4kxxsx9+yGy0wlarmmAAKNn9UCSOrGtmypyCwKGmphiNecLER
VfJomyJ4x0wjGxhoYwHLy7zTrAfeBPIoID3uPsigw10S3itby0O+YBpuo7+fqFHuaYet1iqEsE6f
1JGkOtbn6nsnxYhp1iQEYLyCRDHiD8MdV89NR1PrPCOYTwVEBscLV2exS5w/45H1893kBddIVkn4
ISgCJ+rEEyAw8cnNqdghFu8r1Dzae+Kuuv+BwKH5GapEKlBqvbljrxqQcO2ZGCLXr/BnbBCaoQqx
8iWxMRolAQl+J92NIJDwDzMrI+f5TxsDeULczv+6Hf4XkX3bf3tzMN8MqYe0Z45UqRldLhhLdn4t
Grxb4wWCakDa9J/fyBj0avzFdNrXI5O82OD7GfoOPmCW6ZRmBQjLtSVw0dyACtgOKKExwmaNEp4X
2RGrhNjKgHV7l3RpIaYIAUyI+zic1F6VAljqIFhRQ8wkYHJsH4EcTloUnS1ukvh8H82F/TVlPzyp
mD88/DzY0qYpbkT1+UfF2ehZgsnXewxcpBpDeU+LDudCveLCQYofGKvoXr+Fz7XiOl7tnPqw3q7k
nDGrfjCLLbSKZizssC/Xb2ztRrmob+h3GGRBGfV1CoTmX6j2pXjA46R414sPoVOT68kr/zI3NPAF
T686ed1PCx7cnyqNWQwGRaxcNoaYQKACQ+rLVULM0vgdZIGXI6Ba9CQLjtJt9Ucpz7/QL6t8j5B+
rHFGTqSLhagzufSpk9CLQkVrnoKW37rcsLqxo3GXWSqRVck8PP7LLfAOhiqrnaQUqZblQ8+x6B7q
urrEkAcLSYH7Nh4fBX/fClp/2KVZYubr+lpagvqSL1msicPE3tSoqfKw58R1exJh6x70QY5ZAGjH
gLrvOpFLJzEWS3zkwN6HEM/MH2KY3gYr1kivAXNZy3AIbNfMCe8sVYyLQCiGhYd3imWaGJl1zYp4
/jk+8whHHexjRKgHJ7Br+EL7QlicxZ0gA5qaxa8wHrA5P4iqDs1MsQdrt+n/BKL/kUd3odpogB1g
TiVHvopzZ/o60xBTD47ifHVACdxUinY/kD6Ls9pS5ANzfK+zLcMyijDJ0tMcMkxa/O0BAPzyzwvU
rIs841pVkGkABUgWnCJvBzsVo0bvwom5FZxCF7ji4466qx3LFLqQ+pv0YHDT9XgAmfd6Apj8WfV2
WeyuuH0I4Kq5vQziH9FyL/4iqaiFJd/3+ZCpb8/YdZjGotA6mmN/E7xbFXvOQmStjN+ajBB3RvX1
JN6z1p1towsR1Jof4Qg2SwhiYCTxNA2hddg5qejbuCsieqSeGXWl71KKKa0l4ipSxJdbkOFQnfIi
T2c9tVhZEWWDhdoCeKVIXnwrkEiZjU/I90lQwaDoNcKgpoW3rmN6kFeO6st7iZrDK3Pqz3epjrqg
e9tg2lUXHjGqoGJfzqHA7+iZwQgjdgXnoSoA6W3Cr5W5ZjYe+jmqaaLoDo6XMpRc8kR0lZIfM3RI
/APnlFtx9AM2JMKkkgR7tApLAcO3OLc5vf3c/VWFe/ILM7IKcI3K9d+V7CtXWKmwFH8OHE58z5gB
SSyeE8wSEEYs0x4f2jAO43tsoWcJHgm60hgr5AV7jOmxOrqAVBAhqOptoyEn+VytG2Bx+wTLgC6J
r7vPtw1CjX64U5DSZEH1fIpgmJZzmuQ6Bb8NIYDNZAOzf8JYFXQeMLKy/UU3DS1HDYIuRaBz1X+2
mH+bWFf8QqSjmnq+rMX9bAY3QxoffSdYk4x7B9qO/M7uExwFvjuRW5Vq5GxlMjfOYEGWL98/jBCi
6BEYguWTTWpKIiDNT1Txpyv9YFKd29SjCbe3897QEV/9S1edPC/ytRk1KWpaGwfbAmJmi4EYji/+
P2vOgR4hHr6p1fnB19WK8wvAwP5OaGGI+eKtNe/LuuebGA8JWAeJmeif5lvMvypUdOc5yNVocdxz
B8JFYFJaLT+YLvFFk+HKOxXKYPYYDpLI+ZrXt+Kn3OQCZdIzA3N9yM/f+/nJ44S5CJYKbRrbJNsl
sV9eWr3tZ3rnp5uBHRRXTQUo4oztiY7Q6dRvMOKu8H0TBKpGgidq1HkmMRgpp/Fcf2lpjDY8Gzn3
Pu1l4tvq85GSqJaTX6CDDZxctW5LCRH+QvAZb8J0/+NVahZGbSIy1JizhG4yjRI2vpvGrGLHtaky
Q5hwLvhgGu4gIXPYPBppfTMtxG0k0FF0wKuLA7ZSubIbPNrwRSC7WCrUGSHv2p/gYk11T2nf3/X7
lYa4PvyeT6gnF76MEHGRg1BabYlRCFexhetIAL35Kw3xNYXYsR1sTj6bn1is3ZpurzLNFNR/o8LV
h5NB/IQ1Xrlo9akShs59MJiCbdvksIFcHrjeWtV8Bw5BJ1VliDB2ajufJjJSf0g7GfybP3pOK1iv
aOl5tgucaBydAfUGjU5hpvGK4ZdSq3CMjgjsKaxd8psNUny6o1ZinK6zZNKoTnSevlO3btAcJIcm
wBmdKt4YjzMFEArx3tXazFtW4Hstwgyf6OIxO1NmVvZffVGKdEIxhFD5hnk22sKqS3z5VzGtoMqM
c91xiFAdCPtmaZjUEG0G5gv0trKY5k8bXW6pzLNpv4Vkk1ttrg15w+KSIwjLDIGMPVm/Y97LxYLL
GSFJtKBD6ce70yZzu0vkVAIHDZQuqf7yVNJIuoQeqf+SMnJvhyhn99ylmsnfbldZ1xDjsyA4aWls
Z33NfERCHPUQ9upPVWfsi7JSf9QFuGJnn8taBuqP0qC9ayQYorsAunIQD5Toc5HBDZIwAesyw7i6
LzCFgZ9u7fbtQw8RdsChqRJSC9DAPHcvJDQRuh50ESR8S8lN66lICnABnAVfbKK48tiPOv8Wg0Zt
yNIYprOtKQ4KyQpPBH7LClOFlerOII0o+xfwSrQJVtlEUtqij3pusjQXPblZB94Rz3jWOYmIKVM0
MjJ+c3rRO502CfZ+UF1NpFCd1D/iNNgNMZzaSnPlmFht4F1zWoUfgvcXWaqNCI6F/W0CCW+NEs8p
gCHYizF3TJkr5kWuhkhVvAsY8oHLwxmMcNcHbEQ2D+jPblV31ttgDZ+BEHwaDQgqWuGCPvA1gjbR
1Eq7UqvR8Kee7mi3l9K8NRdS5ZkP9+Zf2joFO8Sv+rpQ9uslvy6bldDBr24hbncWODRIjtlIvPVv
+BB8tqLv8Jb/zT58y+g+wlEJIpBkD/Xrb6MMJKxRcFBzsDLG6tvn8JrBdcmUvjBaAJtIGjn7zsca
nA0VvVTp0za2m0QChi5VelbySl2sCOqezOP551EfaTMza4hs0fisIg3bp+RtQC1s3Pw4J4BoxbJO
Q6SHD4LGmu189v1Y7AOtHC0QEujkkq79vubS98N2z9FwZfVZJ2jtxewD5eWMYaS/Zl0l9lOjOzih
Y7188BeA8tZ+vQCuPEkNgkvCnsDkJpduWF6B/6fOaS52d9VfneuAkyJMsFY/cFXQzdqg4mbMj1md
ccv/US3QiUrB4TLspnAUrruEOBJStz1yF2NzMK1zNYYECbKa41ljrq5zlEHAv2wdId2KhaaSRdRC
BfBhrmzHXVj9JbBwuUBeWFQj1r1ffu3G1mdOo5M6uc6Z6HeWMMVacQjdmc2WclfmRxY8IeKrBw9K
s334m18/rrbjtxrXSbm4u1zbI2NAhBz+68M0kdEMOuOd1nqgiV2A87kxhbMGEJ0WIUvpKldIgNkg
MrDrMKDc9J9SKodiUcnwdFuW8MystVhn3IFwBB+OPcqYnChDBkLj+wLiHWlNOdQjZmkWN5bZJddu
O2mLZHvd7TbMYFhmvsB5vfDBuhV4b31kae3QJKZKkD4pMy7SMxH7zUUoiAhzBy5+MVEG63JrfpHw
l4tJIJZAvjlNdczvM3cFiuFNU3TDctWpwzJBI5lMUdD6Zap/p05RwFUNoMkQeu5mpzkumQ3Ro/m4
mu3a+RuWKp3J9wFwiHPPsSIvBrFnNcHbP2kKP5145+IMnqn1MXl3e1GE4Jvfpk5GtVVn7HSTva4T
qe3ZkwY9QNF/h5FY1N8c8NHmaQKf1CXwZ3IAIMBApaEO4G6EDftdEwLq53ZuA0lVsteGOtkWUNdT
o7cQCFDCQtfPaspnQJUPtUnzdkBsFP74l2NCJbK7tgsO1/MaJ+1p6V3vK3HNLAOQIrjE32K3YIFb
0g7RRVoW4OTAh/zSkEdUM/rDjHqpd1vCYu7TClBLEjcFIYUUyEwDNsHPsy/5yD0GaBI3u+nT7zRO
K51ootJsoSe9aV7ChmJBtRNmcX9opftqV7dl7Skvyzp9AwSCFyWuWZ1kyaI1hYv2Dr99AmFF5v7z
/MiC54eDTeMf+Jk6JWGdcKpZlzQyn8dWNHzaoqeni5TKj2gb2bw0wKYnUIKuadFBOn2zR8sFjGlf
TrqnLq9iK/vKOC22LtdirAio+auSuv+lLArPyG4WyedIqgahty+kKuWXoPy63GD9/rWOLNOch9m9
TzdlA8barONNuXsHiX2O0KdPe9NfgEXkmLjEKSpLHWAODSa4iVDlc7jEvs6x65riV7O4JT7PuLsf
t9G7VbGGm13CJ0HWM/C63n73NALNGiVnEdqg6wdyqZGVIGmtXBS8ZFdXuP3AfnwqrJwx8ZnOG0JR
8RC5KGi8eh8ahh8XUEFKr+EjTGDKyQ/w4MjZdLPwPlcmHMbHXOFyaLlglH8ntFLrDjn8WJi4PxdG
8RKjg1FBHZj6Z8J/uufgYPPWJHty8MdXJ20Wi43C6J6G+MID9O3+38lMeLCMCNq8Jm+WMe2LDQpC
s3Yv7XsOCf8GoDgnfTGE1pkzx5HUwqkLoGkNpX9Zo+e2HvuVPCqljOGoShEK7olo7zTN8Gn4LDwJ
VtWXqb7a3vwCLsKD342kxU9Z6euI76xPv5gRz+QTCq8IQ6o0IfiDrB+NearhRC0Ly6533IGw7pV2
38Pw/53hRtbLfdpYbh9wxE4Ls5VbIZmjLCqNS43SwhplkBCE5neUoWApJ7+PZCzAJr2tn7ElJtxt
Fgaqs8cwX7ea+cOfM9frS6oDrQh4zBb90VU7wdbhkH0zFBjAoP9CmCxVBAreehywFxFWRyRE47iB
uVrP7rit4Ncb9QSM7n03a6PU2NlVc+++RimiplkduJyxu7YR1zip+SZGZan2CICLjci/YBKpju03
EHx+lUYghEVYW1xS2sIZKy+ZmP9Cya96TvQw9nscJbpo5lHTKDlT4Ew12Ee0gcVPJ3gz+GnutvRW
z44hC551oS31JryZZOWIYh46ACRZHaHpj80ot8cHfFISUjTIPcP1haJrEDnEnWsBqyrILEE84Dnh
CLKllPNctm86yfw059dKFI76QP0KoIKXB7AW6VXQRzg3EVz3TnscG8MiYM8fUX8i39XqA+Cpt9qK
nCNNBMyPzTTUclx0x8olVkvhmdp6Df5iATawzvGEqIX2/Km8sqaaGkPfaI9omB3PM1O6eJAVA21j
ZOpdtbhKR0PUgBpCo2oC9+4gW2VRuOQg+ptgyfoFKZ9poWQuSff7Dagg4OubyTBcmTXqpbCaJzAk
XmzcEboe25/VrYboToXsp/T2dnWqT5EhCz4E2ANuRmz8btW9QyAvI1/xzy1DiZ78SV2vYv3JdGpn
Ir+pbwNlM8W+LZllGOegKrrLICKm95m798fBOSGh27bs/UB6QjN1DygndwFJLN4kEtmZhW8Ncb+A
Dx6ngBbmt0gUALDnpH3xB8xoZJpM/XcU7Ukl0m5LITR5Oy1ayaPhs/A0ErKKR9jHYS6xJ423dWuk
7mB197Mx/4zne8IPm8MebWAkRjAYzDj5oYgrHHI76lj5UxaAvdi9GMfhBFkvtqhqx1Gx4H+a94We
aXH7mGRehPGQyAi/3iUiMXSIIEpxOp7kAm2zjVZqTATrni0ieIu6HRxDc3za8guRvMUeyrw4zRYK
p4sHHu74uW8y5Vx148Ois2BXPZDrCJUSQ/I16WfEDo+tdW/aS7VpRRBOO4n6OvwpZqKBMRY8sMXx
H8T+9n7zmaXbbt0cb9iv0kcYi79uetnm0tpuTUntVNstKgoAu64AkyDdHeU6/GecNc/D2Q4Snmi8
iSfw2UcQ2M5aJbtizT6qPrmdesCtBIdCHLk4D23110wHDYbir+KtkkKX+8PDTYL52uUUgtz3Umvb
XuUbaDnkI1XQAFJAz2Sf2BzXk4wBsfX/kFxOtck3x+WqAzqCGgGqh5hqluIokOCa6KOyBbRestFr
KM5S7xchOylQfVJnxFnfW3THnmNFOuhMbLeliq2MlYb2UHP3qHsKtMAGsbGctgGynLQ0rroxd6/z
CuRvjOSTAgjOieSFrNOL8BBeEzHiaU52ml6RGKQ1NiZ++bZO7/dxh469nO+iTJWfCBq3SCwXbdAp
ltq6eQu6fm0qjm8+6UT+46XW+8qJzsBQ0rmYTvAbOlItMIWWRm8gkKy0lMrZavkGMvVaEugWCOwD
nxubAAFZalbtvUw4dcmw4QcNFie1GZsCL7pGU+CLPFzLnbushHgx+Td+a4ZqxAAVMK+wPTed5mhY
xVogE5t4cOjIZXy1rzwqqjzWcWdUoCb9z0HdBvWoNNcFJ3HIHAbR9TiVHRNTKKHLx5KbS+c/3Zl/
dJIcG5LwcSvGYT9nub/R/OohYpvKrixHkFx7tvZIN+Lb4/rvxGwDydJqdqqbQ/nmGTeULA1RoW08
m4Mihy2+Dwmu1VtRq1PxBJ/o8IiZSB1o9PhkaMjfGFX+jybRKJS14ebwB7LTmv0WPkxWWVMlM5ET
3kxZxpj5mAoLMI0eg4B2jsch0Vqv4BKeOWz9EaHpKVD5u9y/0h7P5zxylApJpv75oEeygvr25Mb+
28xKZoEIZcw8RmPz/bhXmmij/UvMy0mrsYkhfGGznDqbHmPKB3L6IJ68B1WTMD6imEYw/t4U1joa
Rch8IDV43cNv8Gxd++roSknwF+jGS1DjU6MCx7udVLfDgXXaSxUMQtxQKpoq1RIAeeKMi6+QRYF+
RD3umhSnMHja8IvnUtil/oNqMjvYqRE+l71pdwcypl/O1fxwwJiqKsimNXUvC8NyfkwwkEfIbnmB
0StM5rVwh+45OpffMf/gFugOFdIVxPyOMlttb3oesE1ht+mvRA9HS9VDqhKdW5dKL/Wcnbn4FTko
minI16mdUPDtCBXRIfwltdWSjXTLAVpT0CTug+tRjy1GkIFNlVlrMyo6R0Hl1V6lFE/fv41WqZeR
/Fi822CjpRKz8c1tnSOvH/mcUAN5dzcwqDaTB3Oix3/4I7ftFJcqdLNK8rwckpacUt2809CFhsEw
GQzGU9y1h48kBosJPzTivDdt7AA6pYD0ImaFF3FRYZESO7Z7uQTQKrfb9nng1F5PrTc8+NafKYCa
VziRdNEvw8y93BSxvNm7UK/gkXiwAZQi2oLKnnoYK1AqfeCY99+Ltyljyf4VdxeDchA8jr46zu5f
evm/ZfzEqCCRFQEuAEvKr7lBfON1JYlZpx50kGyTzH+f2xwFBscYasdERba6lhf7D/evN/wUm+hs
gv6uF7cx/eDd3YM5UNAAQIssHG9YqSt2bh3nc2J90PgtrCpE3h7XjQJDx9+Xa9hd3rEBwjy77LNW
UAfWTIjJm5tUssKvi+aDZDFVZJuM0hzKPtzyMXGjo6qEbcEqrr2iDVCNypUVT8JlAlWBVbWKXa0c
GTcallnuYyH+/a12AycrsL4B7NfwNOL+q+Ui/XpU1EEN5u43QyzQogTir556iogJdMDqsRHPsAc2
3UCecA40PFKTTb42jPBZ6Bw7CjqlYsWyNizjsZrR3ckboYFZkhXqWUjuSv/GVE1tQu6FeQg/cpwz
YDPbpKy8LmLp5wW585DiRSpTRN4DxvciW4MUg7pMbBAQ79ldSbWWsyEKW9bA+WtgJ7xU2TJbVxoa
5DhEzZUkKL98ZbqNaagQff4PIopaBL1UtG4cygOs26h6B3s9qJtp7sqA3QcwdCHLGiVpPSfYdane
GCXCkuVoLrArqmbUkvKTYoENfowp5WJBzwAvFQS5wP8KGExe9GF+tN/CZ3FvlxI9BVYTc42K75bL
3T7SVSIAEqYpaQ0ENGTI+BhQZmgqqM9nXsbHnbJGvSAVikSh2W3ajw03ux8SNf2zB9dP/yP2+HlJ
VCocOOX64/dULpyeqwZkMHWOO01SuT+GBBnTUAwFTMymyE05S+XJz11ApV6Hg1xIzsNkXyQqouyr
KFKX17yEA75szlLuBKdnbLj97SeN6X+BuzAOurqFB3nRN8jyWBPzrdvhEsPqpBTZcfyyLWqdQAIc
Uf+kowmXPZHUhvoDr9IJLLtywRfOlcECRAbHLFprNB+ZZIxtX+3oB2yDbU3J2suKmcJlRC5ffNm/
oR4VGyv6ZtBBuGV6QqTZjvS6kzyr5j3xj6zq1m1+6Fk6GczDheIIj+vqJ2HimlbYJlQGIlNQaTWG
Nq26PFNbLqAFVVlktwEz41r+oKuT65C3jDK+wGX7z3HGzsI5aBwc7FmP151qryrdBJjr5j7Mq2xM
3XLUe01XAPQ/hO7CIwH7D/+Pbp4cI8iRLCOAJP47vxzgQRx+P9eivhhrtIH1hY91x+LJi8uWIaaU
VGrygQPediLJBDIcMb6Rw6qSnWydx+EcNEdGqJ49lNrm7JKMA4SGt9RceB9ix/7KPlnHvyU+OLLi
WiWzhdewyt9PH4TwA3hm81pvZmC8pSxBhRwY7C3ey3qjf5mV1Y9+phPpuXi8gCpRZDDuv24YnkaJ
DkUpgpnZtrK79oMKE6CduVD4nRl6JcZCd/C2r8ZmxfpvUInyF4xMiWSiHpkPTD7GMnCJ2i2b8LEw
EAioY4DfsvwZEZvXPD8FUoYt16djxw7RBMIRaRLqLQxoCfBvUysPhv4X2/kcnAdle5nIExqOvsNq
7Rx0bRygZlSIMaJiSyvqfd79pX30pfpzPGyNHKdUDrR/Kv6aVjD/vParLDtYLfDZVI1/8Z5tNKcO
sWZeXEx5M0O+IPAjn7TapTATODmH0CEFhBWhR5EQZH7LHOAg5OcgK7OGpIBmwPVR8I0vARKi/q5w
lZgLsgXgjiCwgt4/TwAY9ruTMW2fOB6ImKl5seikh/5P3DWr/h+h+NhkcbOY+LAuzbdP41RkB5ab
Z+AEUDOBAC5goIzRyNIh3diXp4A3ozrZEkI8rRxkehZHOeOpJurnOJCGJUxri5czM8aZ1IqxSHJg
Zy3+rrUXholQ5QTWMpEn2lNt34ACvp3rXJ4dSaHBriy7WEhojAuxDLshyUSqcpkOYaz+aMlH10rc
0ojxIIt4MzQ+6NTrKCYgigIDvtCgzNiffG3n7Ef4AmosW9BFguJCQMMnRjrZzwHxB0i943lAboct
sOF0uZ8BAD9soS5WMEllGVFmHJqWx+seYJlbkUXeYZjB2MpHUz8ssmSHXHQvbDSoDNZ3K4IGfglv
l4IwEz6e2UxjUzpRCAQaqcJOJFYV8KL0itJGvnfHB0pLIrkEGSFu13hbmu14e9TRIktWe0tAB/v4
ig+JDiXCHCGu3QbK08Cz/3G9Ppv+6XTbBOVf5QYN+fbqM/IVRycr5rJhDXLcx8bbdgv/+mPGbeVT
Kl6EEBeW6gURWA+M49f1YFWNHUilpOf43ghYUS3rV2LQtlpIeTWikOnhFZMSrjC7ziv3iW+aqKDq
KmVGQvciLrM6swHcmuV57eITLsFKaWtf6AaBmSHyUNewfQyqyuNgnsAuh2Tw5ZBXaAZEVfFoDNHj
SNAA0MQ3YA1nxY0HUNjkz+B2FxbVp418iiSWpgp3wZGB5KGcxIpquc5zrvudrJUtlRLJXcc4Jk9c
rvA+G/qDWygGtQDympDLxA+x5HTuAbR0NjMY18eMwPy8fF7hbsgFT8WcAZwN00YeXOsNjTWDj8FT
Ua3SfvOiaJwZKIaBhyxzGM5ykVTlpb1oTdRlZzvZgReK30FleFxLXeyMOyqRzYIrb/eQ4l02HCJz
yTdjoA0RXbsFkqgodWfcU4zd655LVI+wyQYXdLOhx8H3vdfP1aJJhu8XtmxkmWR1j6JpBOe/hTMf
wplQyNNEgx14lIdvvLGHzTY7obi9g/tl+Fa9Oy14yqXdRcRtcvXKXHUeqxg/a+K32aqQML4dYrJr
yftFeKoDTDarirtWQ3G8kH5lQtYksUxTgcnqdZqzJI4CX0sbDA+LMDt6DZmIKIE5HaSCU3X2fIDH
P1ibqcLtGgkBTKEEneRT7ci2gTgMB+WTsBJe3j/K/pYDZUhWajzbgUzXQ1G4r5VsuwGT7VxGJ+Mi
54mTg/WmASeWSJp3ICNMO6k80QDLssOUvv6f1R0d3XYidKPqpg0+aDZizaP2QfHYzMPmIUFMVzLA
yI9kknwpjdYnb/1GowjoA70pgFvUs9fwVkz35ZpWuVhYk/cTghUwTIoMdLKa1teuObE8uTsiuny5
noFDFG9+DWWiFsY5w3BPIToRFF9rOnAlqjGCRn9w6OKeRJKXjIOyCGv7RufIgpXPUD0LHjUsWS4G
xqwf9EA72QUiF0WSSPgEpn6M+lvTODsR2WMOYe/DR3FawFSAZHbIlE9nYQPTw231gwcmyH024mwg
Kn3lBXoCAUqq53Kyjfz4R7M0OOkiKXKTlJloOFbYHuycD6woZ6EWbD9d3+NHgzsGAXfPxooz6TRD
HsqJzMi+I2jvxcYi8v8GTWaQPrW15/thFg3s/jWbrHe7/Cp0u20znn+B5RCO4V8eh9eP3kfvqb3X
ICmHDceYuEnQOpHI552MGJo8FxTTU3P01OFfkaJjogmUM2ZwvHV2R0+QAj7FrXPLWCIIjHzPYRMi
PDKvrW2knFeqGWt6JBbx9aVKeEgF6HLQoXzQH26V5d/bckW8wnUmqTVoJ8PDrAwDtQeJk131uc64
9yWY9YqA4L79/b413nUj2JupT74ceKaQufZ40Lbp999LSllWSrN2qykSsiADo/slhM31ZuhSB7Wr
ao99aavrY6tXNb3t0aPSBQLORvn3QZOANtp3aiADCtkRuJrJSHPZxIRuXUOm8hTRraXA9W9RiGAx
wnmWa935c4GzuVZfvNAZj0GD5xRul/4gF/m7m9bBsG1ZlscY6garmXWHd4xnkf+AYKtWgFzga3yK
HZ4PI77esjDzC4W3dZehqSaLYbX511sQLneZSmO5nllNUwlKpsPwHa/kOeFUkePT67oOSHWiEJha
oZ1QT3R6aVoYhgXZW5NyTxTvGdja5v4DFm/LkRaGM205R8AZm2sR0Ns1Gp1RcNCs2rcNMehdKfrO
/EyQcsxz7C2dwHpMg1uCZzByEFp0fvUC7HyLSKLOwtSgT3exzIgOKApNnoNDvZpvwCLvsieehV8v
H4soFmKKd9lXYkbG2JVQYT3/3OF68POU3C/IbZx1+DVpf10pM21z8lSp5RYfZmV7Iq3RltHiuQB9
3hH0Tyigh6eHudDOXRQZeQus+E4p/gIeqV1APrMAWHK5Bp6eDMemMujDEu7sR5Qe1U0Qs9bEz6YK
5hJKzCdE5rX5uwShdBovrJHgUu3P8J6tFw0qKKCtMz7K++I8pOB/eGUcuY4mGlnqVh6m0yA4SzUZ
HPXGdlv8puSnTS81kb/kTyAAun69MyE0t2BuHBObgyswZobDy2a3t+PbP3LPmcFy3zIkM6eepp9Q
vHu7MqMZO7LFO5TD9wbVso5gdao7BlB7v7AKDcSvSEwroWLb2kB/ebpS3spucQs7p6qbHyLdfBu0
52RxCLYY5vt7kANAg/KYTofSaDMNQpaWb82sxTVTQy7sWw5xCGjJxIsO1DeE1AF+lWe0WLQ8PbpK
Qx34N+td/RwGGvHqt0Q8bTMhm5JMFY4oyyfdxMrmY5lOB5q+nRGOTgLapLOwDwF86z6mnRylRJGp
ShFtTIEKUlKHuWvey7JNLJybHdsp2sM1Gui+2z0xZhx6vL2mUmc3f/HOIpj/nnWBmxyQOzYc9Q5U
zjqL2JeV+cUoUjpYxuOzRE9kfO4DQHFAw8lS/uLJ7gjyAZLNK3Uvi+fkXVlQNCYbTZa3UilN+ISi
Jz7BKGWXIERuOpjyW/4VHOq59LsFQcSQpvfeg3k8lSBGlAX4VeMCorwJJS+mvLBunAPjzR7CMjF8
KQLM7xJfanFY41RZWXaHLp7x7mjoKHJyJOrzw3FO1QMG0vnQzQMPXtV3wjJLg9EO2VmxaNEQ0s/p
mjjX5prjXw3lE5QuZThHdYPuo3LHpofBVdFBzpQKGPiGE3mNfXpvsQ6JA0ZOeyh2w957Umq5ugns
52VGSJ9PjfMRGHkej/AqbuWA2VY7qGv1D3J9sEhiZlh4wamcQV0sz0W0sUZ2acJCiamtQuJB1llf
Q+fF4K6OG71RNCmnY7mzvmypmpWsaQDWsud2auRUDquuzaGI0xhm6AmHPncs+mcyQlil0h6H5lSp
EGxuH5Ssoot4mB5TmMCgh1k9TwmYRXU2H1TeAzjmNjAG9vyvVc2pMSkJI+msEkMclFSv8yvODKm/
4K83f/IYd/aJ4n1YE1X544WC54KCIchj/H+HYsEmCRoQ43u7AfttnubrtlElLdtWrFTnE7ixeq14
1JgjIBo7r7wlmdfPFpW9G5Wj2XH2hsrAA3u2L2fdJY75oA5mnEZbzzmiUM45jTDCmSJHEP/XdER9
66KqfXsMAyMP56LwZ+Kv9Rb/hDtcgTX76h0txAvswSw56Tc/guvBP2wDVPr/RPCV8+QhfTmeATY9
Hd7kgAgQqAQ+5XXBTFXcaA6HgkKEvTgaJiOyTjuGEogyjPVhhIKrp1cuahew8l2pKaNILacRvjdU
r8nqeoJM0o5yHlGyygG9GU7pG7qUuOLijrSo4Ck86BdUuEv6DmKykSQQy8QNiqEl21A1eLDVkNkW
iDWwvnPaSq/SS0JuFndiAcCxVMYiRMRE09vJusg8MesI+cW46knKZvw7g9F/BAEm4gbJ7BCNgB4c
BhIezMl+VoPK9y+s8nKblVIYFMK7rqs3Gfyrtlpu0cm5vBTcaGTtdicsYmnd55xYrQKaTJNIi+0h
t1fNvJdLEsQmNKYGcA2oGpmL2s1dP0q/NQDwdvPHF195wMsoN9xjnPj/OwT1Mb+Aa1sWpAphzexA
8hDZNAWUI3RIVDPsY4tXPKWtVZnOit9crhNPkF10NvtBPJqkYKm9wKEI/iR5SJBSztU0DF0PRgii
q2oS98PJo+SzHOMKI/6/4t0S/dtFwFVnxd/pa0dPf4/GoQCNIWCiQxtbDSxZ2c9mwakKcGERoXEU
jktv449x/t4CDIBFzEYTvHlY0e3Kp/3NWlq65xaeOkLqJaS+SqIQqJI/HcSjGVwijCWwbuiYcKFk
b9INs1UNdps6tKTn2gkVIHdPybaRZz4T5GHB2PAR9qd0WTyNy08DB2kttjkBIXTy8gBEW43w6Az7
4tSImoD/CqFStPkryBSC9aH4F7dS1uXatM4F3xINCqx+Y4cl29KD4NkazmxG0M4DXOYDi4mlrMxI
Gy4ZLALWCmoCmAh9BogerLSqkbWPDsj//+pxnVG1nBXTAcGFZKTbvB0CgNkeyYFg1dnWT0wRkGj0
cEuxv1oEr+3NZoV4yP5Bawfo+fXfeokKl2nYLhYvrKe0vmkeSP4CF0Y3BcQ6ojUGkOUyYT2H4Zg+
QMQgmuiytFv8KRN26x6Fk4/s0AJyfdfPWpP0qNLjcVYVn0m54tBZ5J6aB7F732LaI6EjT8QdAI3z
pvJxEjQlhu2R7ZFCfDEVMBAsPMdQx3XGWRDMm+eDIQnJ52aiiydG4TXKKG6nG+CYAIvbTwra6LAp
kEa8t6B3zMCw/ATBBOK7XuE5AFxQb77CbxRVUgPh3hHeo7B+h+oUivWpp6aTRl8JURFFk7b/II+Z
8z0mX4WFiUKYGbfhVQ5eGS8UivdKIEb9q0eJkAw346H5mh1ekviKyBm8lUDZg71ymRCqeasMdd1u
hyDLW2vlbZHg5P4uXQaVm3bz+wSOEZf+83EOPLSAGUbNBSMhT0v0xLMbkLFtOuxsLTHIZHCs71zW
MCN+zu8x25YhbeB3Nr3uYvpZxN3rQqnHlXpSOh5QmEVkTD11Jz36z0QeDKkM8bTlk38sj6n3CeqO
hytqNnHS4RK6y4RkL55Uo8B57oyisKcXceLSQoKbgctq2QxljPGaP0USIqt2JGpDdAP+xsIJbPoS
c3iNTNnHbCDSYqZfJV/12QCfvep/TqUZloA10o/hfK5+bTt3uaobOTFjrTlRwqXDG+J17iT/fzzv
ItAdyrvbIiHeP2igcAbMwLByohLtD48xPO1pVIu+/IB8hpcOvDBrG1lKm23lc6cPjser2oonnq5a
xcyxp7m1OOIwVe03i+RNS2kLUyccLv9bJoLvhzRzV/bY43H82Di0uOZkKAp8mxp+IbohEmFCRDcr
wA4Aa3rmGovP3jl9XTy3ZPeQ3pKMfFbxDpfblJhm6TxunN5T7BxvLDgvaIwKNpl8c69ehEya6Ypg
QzqkgKiFKeQnDbOGX6Bn/ePlnL1slBVWnEaGVLq2RH+N4WB8Kboy0ExMXYbmUlIUu/g4fjxz/rCB
TNkRDSQLbNSU/F63JELbieRYYhDU5iqdPEhN4+H0G+S44uO96Tv+lOjp1e90VGtQ9cid37D+QfWT
iQrfB9+cGn74QQP6oOoJA6MWR7H0lsUTX2E4S3Kfddr4Ln4W+/NE7HHpYkBHojlZQmg/Qrf8fI+c
gnf/IqBYwXh22btGQWoAqnUFD6q+R78VA6CPL1y1mJVDyxx11jbPnxgsf4RGBTtZF//4/Tg1JeRJ
o5uCrGzl2WhP/RFpmZmLDxxHBeqtN+IhHpqlr6z1cxQhWzmTVyoow/gnPkiCk5yoev3eI78Mtyhc
NxoTYu7h7rF4naPzHmmTg0m+xib4gSdnyRSCCfiErid5vSKA6fJsNs+EaW4VkVEO7AR+0SRdYwtQ
JdsBMntKyNJFqvtnx3+ThSBQbdNx8GXu1/Wja9Y1VFWMMAoIGx0eSiK6WAXkn2h8UnlHIwOKnZPt
Gem4deDfjg6QHUXBoT8A+/tUgqYGukvyFGSiygtPaPU6FhYmb3phh4NqZA+TyAdQoW4cOtlkQzzo
BoHqy/H8coKLhD/UKOlYSb1dt6lNzqRhbaOfFLrOobNL+fxp0dNcFtgvXArOA0FWny+rk658ycjX
JVMv6Qq8+qVNT5ekVF16KyE2Wcu4FLTNMYVqTWDq8EwAyUMVWTmFoQxQC5xmHk0i6Z0j4lmnDYdy
VX8S6bUNLaqOHZBcKn0BidOIAKSXDXFm0w2I6BfdJEJRmd48yN8Uc8o5RAiNPHnSwUbqS9nPxQQL
UTbHeTCTgySfNyMPcWG5RgbmDKExsZvtkhLDv4hW1LlaeBEKjdYrhrIpIzCy4k5nYfBcQ7s0d62f
3l+Ub1e4Y0vOY+W8XUxef7Mg79sxVUYLi+7KHRnSpEsKliUIQCvoNqY44pkuvjC1e73jeEsWj8ty
n0bFCxNdxUbFZ1P+wzw60oXtdFtFPJ59HJzPVTui1zn3THkzTk50b7qnQlzF45T/J6Lv8qhugGOh
ehX0hsqmFNYSFVel501oHGMBIwzvAbFzRW6IN2XgUQDErWWsRLAMEDoEa95ERN/921ln/19xZKD9
LrCkJhHEw2m+Uztrv6lxZScG5IEPYGQ+bFbmLUWZj8iosXYRmY2EPhjzYlOCOJeVgegeNNf25T/c
x4YczOKOC951PovIA4IcVN1XMhsH5lHrhfFptXNHRDc3OiXsKA3lg6ClaDrcqDvz4GoF7N1dtT3V
GIVFvTMx3yllMQOOqVdbnRrP4uzHoOYwB1U8L2CrwzPGBvwevQq5+xpJsNvJlle04qFQppNSxx6J
fi6ouGjkjVeYbkenZuaTBadc/gSSqUI9jr2Z/UwHqYKFW4wuRIeE87UwyRPl380+Kai53Vq4NYKO
D/6pDR2RXDctCHxpOPQ0joFQeh3aR7E+R0Kt0d847ft3uoS8UXraQBtEtEAR+HAVNYUjzmD2GbZW
Z3YqcfiQG6uRswllAEpvSRZXWR46PhEP/r5L+ue7e977freC403TzPcjj/HkntQCH40MKXvOZvl2
oVqspxyku5YNL0lCQzrIT/+CimvGPyUMqXyO4nHdRYJ85FC1+BqswgKP56kUwZmYPSLS/uAT02aD
bHRJoIr3XQLJQGWAQylUdpqYtsqCm/CJVn1Us4ptJbrNF+UDsMCKDZF+nM6GtgmFACkG8JphC4+t
t8yQufTjh+t6GNWDtHz1aVsMGXbajCpxszMyl/84iSDt8LvsK9nEX86L7eo3YFWdPsz6qXvwBB/c
4sYz+DwLKI7o1n43f7kmFR5D2N5op3g5Q1hHlIlpZNqfqKNUwehK/nBtny5y5HZcCU29Rie430sL
0lljUd+kE3ksgjNVFwXbY4J2SxfzJ+oG6oIHespBJWzF8JwNiVRY/a1T3U7f+VY6Zpu4rWsKRrzd
0dmYp6SgCqDbzfZF3ZqNChPwJK2wxJK/vwK+AIxIhvwrIAwoFWiYiBjMsNFlIBaxwN40YJeSuaMR
saaMuDZo4lLXExoZ5fZAYqwltledd2BDlpZ8/T7VkVvt8Nuisqj4CX6PcCUPT6CETHL0pACy5BP7
yL+tRXQeOZMb8jPTeCj8jow+ysgbZAmdT/CXufEYWd64Ir9AgE5BzmEh/qM880qm4dY0cBAkHc/I
s1rFWW2GhUmS4vlmSmH7As+5sF9HQPAZnI8QIY2gWTIezaFas+h582wjSF3FFKrnd3luIdZaQcMU
H3l2McmFCt/yUapbxk2vg6mD9iSzzRSrHfjGhp8/qsYx6sUECh0zu0OC2ov7u90hwoH60Yjak6Rr
N7eWfFF80OZDEcYTQ5o75/Mi2xBN3ZQ/iKCCwzkye9y5l/2C+x6WIcvANaYDkSPnfxPGcQrtXoOz
0XH+ZoL0YWexlu26rWxw7R2LW3pVtSBpgt1x8hr7E5IDEBw6UZIF9bT2YtkrHABYU1wJJbOblL1Q
bdaP8TUwudVmSE8UgUHXPF8diAiI9VNhpfoUDBgTBQt2ybH/CPVBYmW5MPuMSYaS2iBHDiCH5v1b
UHTv171cx6FiF7eThQGCz21SouB0d0bJuihvlpkSngfmTLVAkBkLvm0Ki6L2sg7LL16GgGCZRs1t
a1kYBa58wsIsazgr+P9vbblzuCJX5CB97B++DsHTkNOVP4l8NXFCZVm5GKeQ35bV6j2UJ01Ca7O2
C9Fq9VYMACcmVen8H5642g3qvlUodmNAhuy25LNO+sjDdu0/yFlrR3AEhoS7a3P+dVHc8QNlQeLT
2ViGYEdZO7+2bNYRm0g8zlvmfo3yXF9ZxvkmflT6AQ2LnH5dlcv5NfzOwKMvwoy0e3yuEqSWZ97y
8Uuzbq+0zyIwuhFx/60JSNKkYHL747v/iJT0V1YtROUwYrk237lE3FweWpNEyZ8Od6ieV/eG7lwe
7VDM0ajXG9mp+Ec5m+37mDkNVIV4kHuvCYK4YIYtpEj+AN8tEwk+zxIlVnmwIYE9cXTo+m6iMxoR
ifzV6DqUPhesNX6Yn2BD3zKz7MuAhSzAowlC3Tvb3T/SnsAjUhWFp9JRSozBTJsmVfHfUYiXPdF0
QBowTE0Zkp6W0r95aENKK9P6VD0tafaRXYmrRt6bWUCNBlutCzma4N0q6o/UhglcHw17hX+qW76e
2sLKKeJl7z2rWOL6J9Caw5MUl8+RFD5li9gGVag3sblH3RCXQjDu2gg5EYGt3SQPKub+6hMzWH5v
D+xbHgsCYO0ThA6XxRJR/rL+XiqY1dn6R5WOXfymd9b3gc4CyRd54WUtU8GWdixn4nZgVcHkkwS6
4nieZ06mR0TTM3K5hR72NHF0FNFp8SQqE8VmTFn1SZVeoQeIWFEdvaMz1QzCkUjolBTfVzRNcGAc
ZIH1MJRHfTEsVigEyr95F2TuY8cZ0QGjBoRABuHoCP5nW9VRvl5ORPlBLDSTyygkrgaZ3EjGIpZs
Yv9waGtNrCy+LyTMSN4Z/AsAb70SF6fmmyQtGwU4E4nE0YXo8dT9X4tGLsUSJ8ngB0Ah7MUCZ66a
ccAX3bV74JVWHBlnhHf6n+rt4wPdOauDLA3uzW62lWc5Gt1QuUS5tmnrsvmwtKGsbgE3aeRTGb2X
tN7yLK340qB1bQDPhl3gGw9RCEVUM/7Dr+6to6Nz4CBTpi/+MMhOUfNePljaWJ+P703xKGlxvnvs
COK457W9JqlaqUJpbK+82hyhBap++pisZZvo52u5hyCta0UzHjQZAg2Co9wS9xol8pjWJSWxVjKd
BIPa+CExqrgMuBF6RkdWRw1pJaLB0s0AftEENNOvHOaXFz0qyunZ6LuDqAYcTiiX9iP9KwFBNT3a
gWMXpC9Fj4p1AUHqBhE4PqelHav7FpOFKrbNN7pk44I56eE50BL2AWGATre1UQHczSaDAta80jvd
Ljyk/TJtoYuez5FkJbZvEfJtH3KYQECboCAUHir9RphH1x1oTHn1rC6tVetjr/uVzL+jU2qD/ZyN
9ccQLN0NpUycYxL4bmDDLJm1n6T8u+kVQYbCTR8W9oDXXdurTu2fC6dwzUlV1x4K8DcxAKFoFidA
R5t2D+lnqiZmGfWSxMyrlgbz8GVaJ5wXfIESckEIYbcOdQPIbCKhKIXDa3kfpMFMVSjuSFHBFOMa
YqEPB9L/So1OH3ADt27AJqPLT3TH52kj7KB+UKJpwyTfL4pyBPv9squCait3yohFQ3wmhOL4xC+f
Kd6cA3RQjlUVHhT/SwrA5MWQBvcF/BNCKrjaG/maBCBjzH9626ZxtSji6xOX7/GzFmMyc2/AMeTt
5u4LCuIWIJBAM6k6nYWLpMnH8Gq2f+kd0ooOt/nVKq0e5vn/ng2qNhZCWy4Sy2rGTY0WkeuBo34o
x+0/0Q0C8VD74849KBtr54kaPmNa80p7dzd+1bm206gjlkggrtjkQhtNr7VmCRUDhLe+mWh6+qs0
bFrM7YWiiNujzoyGtwja146RZ/uLXKWj9kqsr3kKK0Ila+mxOtbyVSNX4W7+2P7vtE4gVhPuW0mo
AApwGJdWy/AmRf7DNpHIEmvwcg6c2slkMmc1k/UYRTrpIz5R7f38w35wvGks+j9VnpqU3Gh6zOvF
ort4EM5Ey1ssZLabbxlMcTiUJWZIJoygxSEFBeY3gc7dLZqeN62a0jrwdHZGHkPGP7goutsR1QV4
VBtmnEc3n8f2Ufzms52n41nrCEAU9bZJmSNlnRtjaR1QOJ5cRkf+Z6m55J+SWmBWNgBkatSzYlc9
GVa2N6iZkyhH7AFoe9205TnRMBRkR+hLs9StLJWm8mVwhLFJhYMk5n1GeTfPmpoJxP1AgEqhQzKy
8IT/pm0A+pFHxUU3AclDfLqT17AN11VOY2hDH7bfWdAdUkj/iW4AQYX3Ssq0hy8/Wot/+5CQfxBt
TkBUM9zNl1b9Cbm7S2AIDSxXI+R+g9W4TGd+bP4D1/g/kMkEcqEFnZ7Gve/GnsxpPOnNfCOzkTgk
KNBUK+FiwE+rYJEXIKgXRfHc0RtNVjvVC8EU0k38Rsk1eDPOff8fujDgjEGsQTOIWW43yTFBcFC/
FIBfQevru1u2KkSHQMM7L9+wCqbg83OUPKLULvi2cTc/1R8CYPpvsq7kaj5N/1JIoF/XANQ2FnxR
c/T5WiJSWQFY0pPO4fc198LhiGGTGtwdTn899LQt6CiprCmXCNxot+bpNCFxoKOKfcBkecyWYX9P
ypTbkbuzyqJO3WFTd+Mv/yrNfMBHn2RGgTQPghkaoj8hi74ZDV3ZfGXeWC0WeQInhB6rfWd5U29/
FINiQJo06wvw2Lu/72ly/Df+zHUERauO973rNOoAJ3kHa50HddoKeXrW+fIu8DhnvtccaMDfcVYN
fD/JKrznvSNgF0OrRVHrs5J2dBhQC1aTd2Juwh1PRgiA/qIYrmXx1ynUS6CI+76PCkExydvgswSQ
awNLipjPY6FjPbX74bjIP9u63E/8kAaJhDWhsip0DKNJG2JHyxywbyJv1e+lEH79ESSBorxj4VhE
MmAYS6Jl5Ezc7xuWr6+8RyPpoFzTVtp66ckaUoG6YW2y1Eg/VscEJIOBug9XHN28/140omjPWyJ2
jelSgcsc2wMvKblihbSNMVsu/AHiDHIfuXTSUAeYmhEiSO7k5fRAk5h09dZwIkFqNf61N6JO84mp
nyRIApxmaTVWlwjqVYo4pcRrykXVJ2K6bYkmHf6DHPNJv1IAfogB4HjCqY9HOlcDqSS7W3Ca/JsK
+Hm7CbRrJ37VnMc8tBQ20FM+8gg+qRyPutC+SvmrdJGPcMFasK3sageY/QCnuyUk4LurtfIUte2f
UZGj0f1UDpMFLFb1ryVpqTM5Cg57aORoW2BpqPNRUKilxdFVGc+r+3Kj/GjuQabWZgaTIwLIWO+K
YPiigQ4gqCm9gIjz54P+KxzmYRn1ahg/UnNC7Rby80y2FvccXQj6o+g2JKP4emicyZij4AAnhslZ
QpbS6dmyGpZNTogEY5DSR1HZNtIxomJTFvEVSFfHNk2laRQsmMhUSkDoN2zAOwSjBJWhIJo9qI6i
eM5VQIL2HSOPoUXbb5gibXN7ytFNIBZQBYtIuaobF1TW1aCvSCOgs84Bt66DK4KEsUy4Y3+BoGta
0ptAop+dPMlwldGGrohH/hYfbzAZTB0a2Mv+IqJ/REwD5ttCkYBVSB+E+rMRemHtCXrKK4M4rj2M
EhepW91RtPmsSMKHyk5oqBo+NA7M01VhJpECAQsv3Ixwa5nAFZyy8quRRz9VGyO6GohvuwG+i8kV
xy4Ms+kMpTvLKq55cWPKRai6PcSSisIzJu8Zuv09KMWmr96EgG43tbFJwkL8wO1kumDayAQ84XsU
/1cQ0zOHGN+Au0l09XPeLei+1vx19AhgOdx9L/x0NHpPLJXE82fQSs35wb5ZyhP0/2yGMoYBIClf
LfXxjwbfp77gH566VzyEre1qzsnV9j9dia0Dou7gZxsFeBCDiyVAw9eJHp2E1qCu+5YWDN4nw/dy
nTwmel1LPUKgqvozdQ8EGJhKa2CEA3QAZ9NG6k4tvUfLkIZ6M3qOab1Qw2osUq+2egndSiSp3aah
cMVEJsrlIUnlqustpBT2XNx72I/gm6HXALU8vNQRmtYz9WM+OQ/eEmJfjn1T82LZ75NchTHT7PMI
JZroQZjCkohNtvSSWCH4FsSMivXgMiLGjJp8byygZjfAMSFpshqIIJp+rWyPXj98CSyVF4wo1JYT
zKFr8Mye65PNNa9yjG3eLa26IRipirImb84XFjN5vVgtTyenWDyJZC7yH6u/nYMuwPY/nLeC3Py6
g2LUq84icMeBDi9eHe0UoOo7TZi+QpiJ2NzsGUeQ9Sgf1jBsC3PsAuuF8rU0nkcBouENYvRM4HLZ
5CLTw2oQ3dkdG4srZrqx9Nj13D2yOwjfbbUdxLksfB1SEofGGgShJi5LUVpeFjFcRqe3XGtFLeGF
xQ28aUNCF2el80DK4wWpslY58CegcxMmgiOhDASUTpviAJcS/7VLJc7r28zl754G0DhvtWAUgypH
q7cXE91ubOwEdrm3GbZvKtzE4ivwtEJneL45flV4fyr0ENa1xh2lSzcFGN87nLaroHX4gAdjydM5
aLVVcQRuPzRaskzflq94CHDvcm2HoR4wPKs5jirkLi/TCbIQJ6sG62qBLHhgpL8dpKVdEC7uPI3O
Gm1DE98Aoebh07mVaRVa5x418UB+ZtsJTdKUFvJQyHMdHMa2N75fL805AE0Ltjw9sg1gXKg3FRSX
2FbfCM/XCbelLfW/IUfbl/wd0h4nMQMP/ccpxCJ7x3/kVQfMxYRdbzU0qf2VidQQ5TwL3DMPaJK2
aUvUOvnF05fOvZRPaXL1uw+AS6AeXtptgkaAzl4knIKeUrOrYWd9P1mJ3zdC53cXZERvSIFaBzU8
kfXY5r+3/Q7DlciUqZsUnrP0d1nqkUeyKh/VblmSjKjSh0/WhWsm0+3O43ko+H35wIkjzbDGTVp/
kVjM3wRKTm4mwpOW1m+a20qfCVsVnusGDsOutjP3p5hLcol9ZjA1Hw8uk6+TIlSUW0A1JbyI6EGA
blB7KcQWOYq1NjZV/KI3LF99AZu6GxwKCgieX6xXtm/crIU4UKPpuj8m01IpiibiNdaXa2SInb0B
/K/GKMEzJFCgSQS6TcFU1r9PvapPXx/z2/AZoeFVqQbKTyr2eGt/3fYh5kIUcEG85oH5NytVoDKM
mOWWveuByQZO3gf6TdwXYUk6K1pAYvR1Kn2AX1P7uCsTnoJJ9T2hFaLkGfKNMoTGJOTKI6A9b8Du
97iBh6/vk2jwcMsQ3vC2eGAqMMNceo1cjawo0d1slNOJRQrJ6N5f5J8fOLrAFYtYw6cqLsm5t/xH
++p1JM8ggprHxYBBaqPAFmQJg/Jqj9bJsPxpY3L/96UgAV2uZh0nz+oCFKt2xnKD1K9TYlamDO80
HqsQtbcxW3jlpC4Zfj/+fEhXhHn1lzwGhH5eoMHK7JCT5PdUHAOMSLuLUoQpXQjMIsUg5xCC/46P
5K10S821usUQIqOK9b4f5CVsH61SrUENAqWhrwdW4FWuDFYL0VzaxhBLpb58oO65ZAMMxsRDf7F+
Pv3qtECC02QSHMMHAs88uRcpUvVUk1EL5J+zM9mh9JGoSjq2GkH4FWUbG3H5tR0Is/zb8fgdLT6P
LIcMtE35qz0BIGRrOhzOjHzEpPTWZuzwgSjOiZhOlUBOBtMUHCLVVzh5yQpd0+Qmi4h4+Gg/WAR6
0bm6J4Gvs+ViYWSnN+tpjOfFDN2DmQZ+Ml53qdxHEQFrjA2r9JApUIvy7hRhToTwJqc009zO35Vc
RDDCd6IVs8Sw1sincFF1NTlzyteYhWN1RIaux7/2Xc/K+6X3Mn3ocEfg290mrNffR00Ucu5aOAmD
SZ/PxuiV0QENeSQc3KSKbrEzm/RfhWCK66y+4nKCQRNID3yDNOg+FnFHHGSMbpDbc8ula1XdAG6B
lBpJxnzrSA1rDOHD7Nd01QDtsyLHnEv56uiLtLr12X5drrx+BGlU6bbnmQy5BJqsRlF9pZdkhdcL
Pr/qP+4g30/k9aZgmXitF+e23cIKVrL7mEpQjmEh5m1rP2tRg2M98YWk1zAbfb96hMepOM/Z4EGM
gFDYHqPyQhG+ZHyK23RZM3iK6VUZ1DJS/rbY/1Qo578PBYVdmK7M3irkfyUcgDMDVev7uMpQkXDW
kfu2cZ9TBnUVDrKlTlzfN9BggcydQmcQJ5OvJ7xW7cKwOJDF33J4H+sFgrqL4zHzub6fre4AL3ud
Olz4AvN5zQ6HDi4mLTrJrNnuRbe4maA/buqacxSqCIleBNOeb97Y8krgiQf4cZu4mpwc/tNfn3rY
P6GYIbTzU86iETjwBrMKnGJ+4UgAmByY7kVa67Z2IuVC2tlEUY8IKoxChmeZJTdia8fjs1Sbavr3
DxnTR7yzteBlESrFIy2NUnFktQAZXbRmHRJSARzclH6sTHREidjhtF/eKYwm4R2XQaNL6KlL8URs
oKcwboN5pJ7BbmnHTSlnNtHjkS0zEkza/lzWOXmiPQeWDCwBcQTuxt/CRACFEo2CYs95Bh4Xcs9t
Kis9feiboArO9TmZFP+IQ0HgDDlfqKRPmA5WWvl70KUsqV2cJVza0fLlt4vZbDtZzsHzdP/Lh30x
VWtDaMcVosHDjr1KFZdRdBN317jCv2x0b06moBmshGVvrHTZq72vJCG5x9iRahH9MWIySEnNrHAs
FDkqSpmLFkyo5Q0TOQFjaEARcSyFysaQ23jUTnkUyegav528NEy1kTZYf7qwiOCfhwESjwvf3lzT
I0gMr403Kvx184tgEAE6d3TDFTQzvEewAD/YhjezeyqHJH1kH+hxXYG6DorkxUnrqt1He9UZXF/c
JiwK83/F00r81CNE+3apqAuD/XgXcbfttYflHOtsyS/e5jkWySgs+c3gUlwXjsZI8jBrQdFd/EIj
B1nYLwn8KoISd6J0mRmi3VUkN+PSJ9VDrsYOSbPCTCuJH2gxsXUpOeHQwpf7bdVRAOqBP+Vhde4h
yAuhsZaezr8U3M/ITN2wVYjokqYMBLSP9rOu1SMVVr0gbnWkoWkLzOSFi4jOARsFrgFHbfKCpuI8
95Piis4CsiG+rUECO5iBM0APcxZzysSJrLtZbqGfvRqR9Fm5YfzvUqFG78YbuZMC98rIvWLrD09o
mfqgxHltyQ8KNOgYR98b/kVmyHPLvfmyvWCWPxJ9/k6xNKGN8q0XIKam4heqUljszg1bA4ftYEyz
J6kqHZBbmWI0NRlABtHKNbCWznK3/IYAUnH83qmF7DGrAPx1XwAGbXw0G+coBXR5UAZdo055G5L7
6CjUn7zqMhT3Ow7Gwhq985Dhg1IE5Fn3uAEyTScjKyLF7RFzexvHHKH5SJjQoijqILPcfknJFIUr
KVdIkpJhNyjVOWMIPegCL2d3vxjRnXsP59esWZxl8KNroUi0pWq/bkJwvVwr7iu15TRYnar7x1HR
IPPWBdJUjh3pIqRrigFfqMhFezIdzIX+Tqn2Cry2nYGsfSx2cgr/XU3NdgqXdctHS5h0aVWYL9FM
imzd2z7R7NSYc3H3neq6nxC7qo5hBZOwx92BR/ETU2ecCqPu5q9gfrJFrjUT46w+rXJZAJ8sPWNs
gUjwikg4sZBcvlsAsHsQagGQcHQKJ2DJoUL6HivBUkUjtEbl5pW8EkFumqtSH9UL9nj0LTmOIDjb
X+53bDVeoOV/venKqZDuilbywlt9Wq+EC6upM4yNK8mLJ9C3UyD/sy2yKp7pdKchsesOGxTYuCx8
rYc2RbKOhg2XoI+DZdho4IPOVPqzE4MOCHNeDM6GglrgTEaiP6mxYeLjLq91mW/5sDG/4N8TyovW
q54j3S1QGP2a7mPZroqLqgGs+xwwi89tnI8AovNMaeGm9bJRY56283hebMzWIll/SVyZjdMqd/y3
T2zeaJpmFlfvzOy6Vc4K6oHQIZ5VcOzSTQZrzNNUjxTyDcGQ1kTUh8HZ45IWTuUDPSz98CuRuN56
j31BQAOFitRIdDzS17wcidYwxPEj4F6D4HWsu7iVPC4PVRUgFWM7HQwTrELZlC9hiGfP+fvvDr+j
UGUg6iVja0MmpC8f7Eu+R62qGw5v02ULWIYZB7BwXhrnGFjYSbGRPZ6TaxuZI0GxeROAvs6oDFr5
gXbrvApP+mzoIoXWC3diq6TVuE09FSCkapMb+4mIqy2hWcB+b1pJPWXC9F1bYeo9y7i4M4UfKDYk
Gs7ADFHUqUJ2CLBeHWxf3EylHsCb956Dw0AuWRnIzQzq4THfM1m6WCjIcjuX8gwQRU7XHN5vEuC5
6S0VbH7n4CNG0R+6wuxJfZdZS57w1T76+xFBlZz9MR3TY7l2HmK4BMQq1AbXzNPSe3u52/EF1/YW
oGvhdglkDohMxPnWtGVZymVwed5IU2S8aUNqc2dHRd+gASi0B5e1In+F5EjMi6ORp0c2s+6lxX3j
N+06H9adGid2qLZxR6t8iPKndsDjsma9IGrXE3sbMaMyGswIjSuid8YDuUvSfG9wBxFQVcIKso66
/iYLkk1Lvj1hg9nEqDEuV7GBGkeYcupmCshpOpwrevdiB4/crtkncq+JfMzeXGuUteLpIOloMH/o
A4siC2FqbUGmoIAakF3T3wSGDzturNsXFTvdHWb7SW7bwWHBIigtRCYMTqrHrAnxuekSr54eGZqA
ATuRQkQ57z/QUkkbI8df7mPxxMtasdBQ8nz8/oZ83uYjeLupI267thBvDfgWlbn8lDK42hhAJliU
3kfhVAf+WD8u4NE/Jiywn16rPv8wxdgyraU+zJXDORkrGTjhVWYdjt/MtGwnHNJGFhtkBihWXEGX
MjkEL5rz7DkXfmTcloAF39uD0qQHmb4ED9qXO7okKHomRn6HWpirGGZjgiMlw73PX1PcKvqgjeYT
gVKWuQGeGXJg296HMfpaRAsVWJgM01UX7GPxtx+emqIBfEtiSwRXMHyR329XpT04UOtkpg/U8n4f
JqOwm/YDuE0i4sfmrvDVKnGroZrL2ZBlqya0Titx+7cuqElYvQnIfkqxnpM9hOmBYjpdGI2aP40r
e5feBYckORd1snFWQTapZfqcdZg5Z/Kkex5f+6d93dEDIiX1oZffdnrLlZng4Oj99LZcDphG4wf5
0ehURzlTOUPQnOqu7jRoawlZ1DhZi2Z2Ye2Yw+puXmYzR2solWTGQHE3Nghp0fNw9E+GTWocUXHz
QXe67BkEHNUZ2z1soqe07f2G1xmr/dnU20liYraT/jGLbFMUEN6sTFHC4qmaG8W0UOVEWqi10146
E/Mx+Nr2krwBSV0+Mk93nrllQDRd2DC2bXxbMTszFOzZb3+OywSBWI8QI6yBhzclv3+xfRIgdKg9
i4N2tzdOq8/6l7Q3/j15nK2FH6q6t27OLnoheUCfTGKjpLlHCCe4rG9eujh/dKt0Mr4QwFsnwQsi
e8cEK/LGiz0t9IOC7OQX30Mlyu1mtDYTtP5dzr1v2TysIjzYkAfQxkktHl1F/R/A80baeFiNvXmp
jfsMbjaejMSbdpzF32L8gw/wEv2qmlS8bO6aBhL1f4FigdS1O9Ar8NjK0ATOmWnZ86xIeY2yPIEa
I0SoeNNUNmQl+ZG5it88cOkvVeOvLllSt04JxmVj6i/ecInBb/wJoe+4yoRFL/6QQx2ggyI4fbkU
+K4M1fV+oMj3IVYAvEUAmSVfV7oM3bfn94R4Crd/Hh2lhgM2t/Vy+pqcvgixaoA733IIopSELjOK
BT7QEyjRAGCJHYusM/rY+jTA0NkWMVBUnTTWpVu3E5kCV7Oxhh+yJknV7gUXakGOQgWKQ9rys244
Q7hjpqv+FndK7FOsI5fWGdgl/X2LeO9b2R/b6nWS02n7K2pllaeAloKEog6uoS/ctFvMjzMXGwRR
rTdYI5q9z5/BZIXXksfl8LgQEUB/UxYQzbx6lX5+MYTs+BXpSSbO8cfAqZDVQf5Yole/gxpJiF4s
5aEj8AZBgmxMDER/X/+xOus+6zQE8lCIJcQcy1ITxq5reBc9SkG+sxbAWD91q44zWItS+XyVMQhT
AHsCnEjTC1iu8thOsT01SM4HR2H6UqOGz5QtErAObnNj646wdvgk0lKFQtSF2CPSubx/iz7dvwWL
1ZxbOMSFxJjQ0mVf4l8OFUDBi5x0A+wcHP5qy60oYXtdEHO0HDS/lWxs7Ffgfb8sTzy4XNQAep/X
L11VBY6uukkypW1bDGjGQR2JAF8r2dnJeMELVA0HOh98NUPq5Jflv9yf7HnmkVJ7zAbSJnx+U4+o
gm3SGuRax9VdfF1uOJH3TAI3FYDLfAj1pHkANTOk+KUszBXJu889kYAs+W0BRYp47GXORLXJu1XW
bxLbUqgSl2qLVXGDemKDFWFncu5Fjec3X3PmMHt7e+rFlVpOOCXeWRA5lAi6A5yRJo1VzuiQgoby
Up8qr9H+FVDfkYTlfOaFIg9XAHAXXp8elKxs4TO+1k9vPsrhlYMRrNnKDSsGf3iF2RHZsaTKbVVx
W0mcJ0BVKx4Xh9Adoc4rI6aNyJwRK+9wuSie4Vsw0iJyebMQArU8pg6EhCgYKRTgDJ5+6m/Ky0za
fkFs8nZ/x8tOZxJLt30pQUoSfaqbgZfA2Rub5YO2hmJwq4YCPZ0L6ox4xtnIF1k97kEAQL5CZ8Fd
hADlldgKEyvpaKTmOGBLWYwAND1l52RU2+TS2/qC6nwK8bFbn8cMu3faz9ybB65M44M5Gis289At
CEqoIaex/KieLh00SMjAMurUzc7BuVzOCifRYUDg4I7kRB/KNGd7O4zCG0aEdJStzWMLz5Da2o0m
PLH50zrBh/cMC6SmObPK3unqUoDU6os3X6rdSVTy8b08HekEz+AfqNDc35IHkkQqJx6LjQbOY7LM
D6WajBZaTSIDM2SYgZS/LWxJUBrMJxgBc9sTfSH70LsZ/6wWA+YjMFOeF1lKxmo1MzDpxAqcjPqJ
0PfSUT3VRzRmKEaohiOowKLBqAbM50e1P8STJqs3hNqTId4DItkPRWn3N1zmwxQs2hXpSkePJL3r
jiWCoxdiL6abZ0SK1ECpYAfmaWVlfIkA3uW8XfVFL6sI//ftVBpI0JMFt4ToaXWnNqb4FGoQ3TXB
Hjo02DeSkazo+UDXNkBzySZ0IHWQWUWMIIjDk5o831Zq7vYwmmADfjmSFWzMrp2foEA+Hg3SZJj7
V8ttSItpDBxJZkvG3E9tDi2tf2PnJvXp0OS0ETzxh6lAfZTekaMrn4DSEXMhfPA+nJkz9txkz1Xz
rehxwcMMhb2sf6CSXECN/syWxWK4BczqQlpUraow9Cp8SJwCjOCi+uNti8CFr5/oTeE/Hy23SWp0
RIGN7O4SgtiBm4xkzplum2WVH0wFhs17mKDvC05iZfC6TlrXsTF6Ph/WYxBKnHClNnFx9dxYriKl
jtyLJoyUI7cyrEgC58C2ZnT2G9eNANRx6g/Dn46AiQ+9C1rB7DzErMW+0Ah+aj+W1/sJWUaZ0nbh
ya5ada7F5Fbugn6QptLe53vki3K1I/BfTl3xtzqr+lb7zLxJfotQIQYfG7T6/Vx3HULFDd/6fAe5
Hu1F/eqm3vBzd0FTfBaUaELl20hLYY1aEc5ggM1AwuFUrqriGNkn9GFEdGQKw4SMZwcrpmtUF43d
8vlsNtoiFL6tAL7agpU1qU6sTT/fMjdhdxv9q7HHKo6cqvsCNaOxvEz+duwlGG0yo6KELoowJKQm
5bbo4P9nUmfuIGdsCnFo0A8tnAbIx/5xZJF4bBY7bHd/OihEUjvZwBbovFM6tT1j0iyYRqvAlL11
IM8NBiMDGN2DmM+qCL0J2vMNb2q0b9HK+kgW4oLD+QFCi/Hl0uDlpWaifpYYkXbQ9y5X6KjmfuL9
UA5F/fhyDGsk99iuwUeSjVVnoz6MD10x7bmYO63uabmPOp+z0HgBfAIPbftQOO8JEpN5vC5yYxNP
wAcG6DR/ciiVp+RolPzsOwq7bX4WnZAuesNWXDAhVT7AHcmYzQIXK2D66l8KVMlBxHDUJ2fevxQ6
ZgpryukFyTR4i85m0fju4KunRyYLuGMfGG8b/EsnyhClZLx7E/eIx9cYhqXw3PxrBZlkO3wnPqy4
xKIZroASoe/Hk/mpDkwNhb0YH8zXB7MH21UIkqs+ADLBlPmhVGt4jogUU8FTGkzjZH5eqniOzXZT
MJPdzCvgOd6yqPmRRgj4DG5iph7JNvz8AXpNQPZdpXKJNidNUWd8pCCUiV73NU97/PnPRjd3C6e8
WmdCbAGC3mzA7edaaWJ/s+aJpV0NYguXz68StZp/DqUf9F9PM3W0XX/f9U5j6f/6HZeCOchYl0bl
GbJEqDE0XSivxGcGTvS78ekNaEHqTM0mb43jAA0s/LSUASE80NEuLxKxQONJJzQ1seZK3yFuQcKZ
T9cV1XdxPahSn4knq5PZqpdblTMy9zPuphZNTmBgxpgHFhcnrB6aX9nDDl/nsUQXYWaTlXTXuU+J
N5lpxnzi+tagWK5erY297lD93RGG81CYSiiNBQ9m/6cEgiMWc4AqEKLrDooJ5fMbIMKA8cmZrTNX
o5JcaaPkqfAkMV1nj52iOxYk+D+GRiNFhZss3UjWDghY9jW+53PA0K1bYhnnOUbSon+0bw+xcssJ
/Q8EKsNsQATAONs3ZRyP5UGtG/3CnXZfOchdv/j8X3MhZph7A3kJBminYGhar6CA8SRE6OZWc4o/
3aL472GXi+jI1hjb+T0qBGrdTLHKbVfbZqW/yhaj/TXTUKe5DF2D6iCLelbhBxHeIW7Z5Vqz3q+R
/I/9HpiPLtr92F6xoX5rZmB0vvAVivCB20IuQsvkxVj9vpbovD34LRl5gckvbkF2eI2jE4Vq/rnS
+0kY5LmJiwnjia2Kwx6JnPcCsMkWtHpHgYmravdjC+m0i9Zd72ZWC4/EsRIt5XWocGgr5RhVfDaF
cB4Jus03SvsHugSMqD8J5nI939mkij+t4esGYaAxuMFKBJMM2+jKT1MZEeaslYetjPxZcksIiqdy
EqhX8kTdqgKOjnVfVH/D9uRNKpsuUOmwjYTEe/V1D4q+CG884yT6kxLOOSczOzZTRcZPirvweRDl
u39+frK91f5H69VGydpkk3z+5imQfdq1IcM9/ecBim3XXK/VEmJWuAH+TzZsVhoqMeRQVt4i8eQg
aMh9L47ybZ42wWCxIlJYmreiTK2c0SGbwALmwtJWIe81D2lXxAF873fKq9J4j+Nlwx1ZgYBE3MVU
pABOP1/l6ZNE7PM+JAlSIq3R+eVTZq6xF9w9a4A0u503QjL349zQLicmyZH79UToeyRAcD3dN88y
aJFLkO6G0FreyJLucqZI4SoX6m22G1qwn0BJfODfGMXTr0mMyCZiUNWZnTzn+kjc57EqHHXPsKD7
ZzmhBdXfPSZ1Uy2WIvHz/pOEi4VIl/NnbnjgHR/bK/TxzkCOb9ImOdNs4fSIXf9od0SMtgd6X+7b
QXG4pQ2ayauqCbmWmT0nZGDY4UgFPr28jm4oxseGEhlzFad1wcsds4DvOgxTxtoYVhSf3yUJvZio
0XSktZdtWWr3MZLOGpSumStFKX0rYiiAZxcsshdeOb55/7rjMJ+9bYr2gZ6mW7rxg2hdb6AIfvZw
5T79erPU5unFYrJlkF5E+Bx9RTAaHv1FPx/c3TabDQcm8Dnk+Yv5kMrekQxjF/PojEZa2WBsbY48
fdEHGrHBsfl2KM4r1gxmZYREG/OyJL8xEZj+AAFaWjCPLtmGzd4OAkIaUaUy6XrKWQbER0/EM4au
DJdQ9Z5XEdd2WAhepcKgQzxv1fuvw38A75zHGOpkbGllzAj8eVSd047eGQObW2Fr4IaPLALECfu1
4nkWMdhG1DGMji/+ODZICNe3ytqA+BlJUeWzyJ2ecr3nI/H43zo35erJKCohJf4I52UUEV37VFrl
xVjdqvLNh8FLS6O0iOZ2QQmcjHYKGBx04ZCyFbgz1PFyYy6h2ov7cQjZoRToZWNSafi3UBcPTVFP
8WiMs7dnOCFumb1/od6FFYZZrkl0ejrpniSIsrlon41gyFkpCHMvi23Aix/3VxvLusEkdWBcT2w5
4qojVZI4kAcg5gRNuSHoFS6nBf2/7F3qh4a1aMpEg9f6RGj9PP83E+PLeWlGlN/DtKQrKZH2/bg9
Q6Vzg8QhHh16fbanr5d0YNyv4YDoMUDfUM96ndePs/L/j4t6q0Bd0Vre90nY+D7m4oyX8l46xEDV
QqeeGPsZBpZs1eVAsT5PjzBo+hrQIb8+6AbgPpAuveAnQ1d5/iHUXxQG6RNtlSTX8g3LX4LMiOL3
JCcz7KIE6SISDS8qr84m5HMr0ea/BPZ1/Goo2BkrIWepICvoWUv1zUe+q+idM2wfmcnBZnolcKla
f5ez2uhYu/HgzX+t+gXUnKjALiYLOZHCu923uOPaJUCCQMpZVbBaXNWQM0A+hSV4zhq0daOP6rJs
u7Vq78lA6G+VqGPMKjjFgMHGpKy90h96G6lgLKd12/qzqEKdGm4oqhjl0oFhLGTDGOWBVLe8xuXU
bI2Q/y2r5Qjk0wCyYhTV6LdQN0PJSdqq2qkxXqc/FlGXi9FJzbqHO3gZ3+7/z5hXIbp+FhDb5Zpz
i1drKbguF5f6v49scJ9yjYKpRCP3erKtjoPPA3IF4gIpTjua60Nzhxr+rTlzYYr9DlEgvciHIJHO
Ex7WpIexaRBuWb+nwFDrhs6FGPxEzqfLltgzy+fednVzlB2Pi9eqK1hGglpoAmyX0F1QzF5Q+oSH
59CFvD1bk3FNhdaDqkjkgsJ3HeRQsXtsEgG0winUcqJlsuElszEYrbMmXUq2NsQEAiOg5DTrd8+s
yO/YwitcLBMhGe7nbnae25T/GSkiRCURBnnXuWQuPgIiA6r1qs5lwK7B/vnZR950UgRybDmob+bQ
KmU1bB8NwUKHmBNx6I7qTT4xzyxa850GLVfhSgjZteGwJQaHj37dvJzXBcYaB8yEUJaT2zv/LPj9
rbQEl6qlRwcdmcn5yRwP/BU8oWlMON2WtVIJp0T5zk4TCkVNREKm+TODTo1yafv5VifMVROm5xxZ
I6roXq3xPbPxbTX87rw/79mNQpxRc9W9YexZgiEKrM0J2/v0POwKdg1an2JJwxCSW7Gp+h+77mFn
LCS+6Us+TUIdJvy8ubqJHntpadEAL4vVLF77ZryYGWEJsD90jqP8kjLgRUqykoLqfpTPwBGTQo1r
f7JNDqtJvUfHRANeHMrvEJbqQLRnuhE2ezyVtWpyGGsVW4uXmTf8zT37RU+ctHFOFoGNI6bTEvaU
6Fo0NTkFHG9+6WYlzXwFRO1B+rEtk8tgs21uUYfunTZCeoU8VVS5EDdluqyhts8DSJkAZS7VuDHd
GxPEO8BlzArDZfKUIu+IGh+gM4ym9T5PNGXF3rvtd1dJsvwdtfXEl9zw9ftb3hiIwfOaGPtyyXby
BNR2tVcCDeGHXiQ2CddAOmbxXhgBO3rrxs+J3lwNOipxZf7chv4m7IpoIrCtNkVTkOBe5CB2PkvT
ijTxDryRtKUvhKNtfy/a1sCUcDvQPS+QHmlRC8mRbY3NDOnHqPotOaFXJ96GwyM2EOdUuv87LX6d
lnc6+IFY0ypggJ0JCUNS/6NAyquUUYStXVESOHjq1ECTmpxouaB+cSRSrGLNA4LCVZnP9/ac0LeX
N2x3N3kogOZ0wrTvzh7y8kirvXBXDBrm7o9u7uhQfSOfW/1nYGqpKRM5d3mF72rINjtzy2oNwgcI
O8DaS5EKCor1aqWkz+dLXUKHKGKd1FXAZtGDhciBlUK2ZBS/EwRFQujcDFJemr+x2xGqgSLmaHgu
/eDh96R0SZwdguTX8IBPJthTrxYeBSgLdBVHGYN7KaitG8UFA9h62HQPjU5EhX2wQX0GTe1hS+Ml
vXoE4ptLPHfbC7gr2BjF4B7XWW4s1kC+WiL2T4tiAUE2S0lhn3Ou5PDo6Mmyh6iXy7oNw3hCHdBz
+UZNuXNspSQp57lNgVFDHFSDO1yrtzULYo6iBtX/mN8IWdIywe8z/BX7FG9WLrNP+BaQWuMFQXtz
YN9ccnH8teQwi4SXi3DO+DBQMVLpE4et8T51YKwv/JlIkL2jkIKeZOwcfAHCsbp/kwAAyU+ajwX0
PkrPxNJh6gRtqWqRvGxoksc2YWu54kl9NnUhp/ktdetHIflSRpJR/7sof5UgHEeRMh4cQD01tpCp
+yyeXa0Mn+gN4wOqLhuxNMWj4lviCqule4V9KDrEBGTFoyaqBRP57g/KP2iCrmCLw23A6X7ctIs+
cuBe3n6QYed3lpAbpvpyeQdg4taYxLD3QVMARU1NlBCVtDyhcJNPCaWBjfyd1VSqWAa89XxUYMyI
2laO009APnB+HXkO6Y04M6/PSfq0n5djhPQecCaDXlvN1N1YlU8fOhm4ptubHwjsx56LDDXwX4vQ
aNcYMpTKk03gkizZ8avbdyTrEk05vyQYSgEVuWxcouzS6vzgW8J0S6OZHCbZYzClcT4QKh+JOQga
l6BhQycKpQr0olATGcI+Akp169OKuNwqcZN5DA13iX0zaxtyQE/u/Tx1n3KW0J/U+F7VVl0/qtiX
UDcq5bhQTkygJ0zwAtBSfHbVvE4OmC2SEaxZhmK7M/zlGczFwuKP8QZ/rJ/VdkpxBC3C34mUxWUj
ylT8ZuNzRHmZ5VKMmAXjX3gfeWX6GQmnmD3+Sa96MivS0FSdo/rpVwjVJQZ/MH6uQhTcBAQaFU1V
sBdp1ap0dDOXzPCO87J8s9IXDBqEA7fWXR/MCP0d8Ax9HkRAkpJSH3i0pHLzVLjhLFtroTF54N/J
qzWLVgt8Od0pbOWU60HCUGH09Drej83uMH7iSH+u5LlA4T8exgp/nSYoRpUn3XS90po+ph+ra4s4
v9ZT1umv36S2ycV7CrW07Hb1LXHpbIU2LlmY1j/M3fPT0cZnS9stUVJ8QSXWFVrZ/xvOjR+STVXy
FSJcU/I24BJFi60Sii/whgx5XhwWq0scOf/VE24gwhQIr27o7UJlwsJ6QbUxke/b6NzTMMfPZUIr
IYa+GjLykbuWpMiDrLtuUlFuuENPqpleMHxZSxhCgN1GbfATuMqMvAUOAGkypjtT8A2F6sD3No/a
M6X+yn5xug6A/tR32OBd69evm0bx50ubbbh+/Jb4fLqJtPvGMfc2SrHfoijO3/J6+tZy79g7kHCz
kndb7cXXfo39tagTAn4Ns8shAtC0bGPzq2CIA+r7D0Mk1kZkD7QT19zw5OcnziRIhYPl5xqMyAkQ
Sb0nQ43xytexCu+HjpCO9kvhwMjKLaCQycKFtRnjg5Oe3vofJHsSVr5M70ttoU5TnSWgL0wQXRPo
TlW9tqiRbCkXbzg0JqV3F0mpJr/P3LHeNgdVgrmFfS4u8AAw/z6rLonJMTS2dTxkw0rBjrwHG7y4
nh3stSWlceiu0O4cNYSEpfVpUHsdJQPY4MJwIgBEQJ5KFJeCvmjMGf7il5yW/0jRijFZxUFJwOkk
tKX9EEmQaNTy61XpDcbl/AztMMCewYS0W3L6A2tsGdXegjaqm6Biai3vb5HKNwioLHqr4pVnkYpx
n94Q2MsKnAtsKEgXUriD++7tPHpgUwHs8gHH3f+jAdDgpG8oXfvyH7NoT51d1aiAllTPWx5t9Z37
86Zhgy8COK6wsTZhHQWhE+5CQ4WFzNQYkZXUOvY7YG4QJ4282gf95FrLe6F4q4WSzRGvb5Mo+BC/
uMOKRv4Sx2vInocnS60B/LlgS3vnp+GM6lMnRjDpKoRtqBPDUR3azkstL/7I5/g9mr+kersc6wXp
JgHQgYd0hq3BX7ntOZlCvJu5GcYzJX1QZZKPd0PLlWHTp64AegExu4TTlQvKZcW97mDciPrMJePE
mRXrDUNjOtfJLkly6fJ7AhJBlQy/vq4krIh3+ZSnvNxZahXz9115kyuIJeoQRjyLpVEkTH8qNZJj
HELuJ3N+/+LtJatCUARlHaNZI6Sgj1Blyq7hiSIdTU04LtClowUg9YE46bsPQF4NuIDYQoNFSrX0
Py/6G0gRBu3QchlAKz6iGZtOJS8NiGk2WjBTMhyiYlgQcQpGgxeSmvrI1oTtsw7H7JI0IQ9JFvH5
mTCk5by3+yqdRiAGItOwarvIcTEOtyOJ98yBXOjc6zS3CaJ2VWSGk8SZNqjtO9OLq1eJpSSmDhrH
HPa3w5OibPbimfp5LWKBydthC2oRMRuBTwIT7ZDIyamPxwjitfa4oYq1u7o+bvXzs1/5sk9PWuzb
v/i27CCCkD5SnRhINEdBmxV6lFvnVTSCqB6SpzWJ9vTjDbjmR1br9VJUA9uJILw/iV4nSWmut/DJ
LOQ87c0EB1xJa7hW2wX7HCyxH10xAg7De12MBwdwnNCV/UnwOgb6KEoow3O4I4iAQixGZ1T1nbdF
eIS6B85WwD4w+zPxN1tKDs5KsF4CyngS4wLdEEiCRyhWRe+jRjYcNEVzagnj/jvRQ8qeshj9gAc+
RjbQRHQNa8b+LgjForoJEp4uOYHmzb1547qBxgqJjq/SXS20v8rKtJqtvRgqy72HfHIwGxCHt6fc
59aJ0RKOH1pdnnYrMm/PX0xgwzDvv3XYKNcu1z09SN+eTBXFFu9hFGsEAqIQvNEGlbNZmLzG9Har
uUIIAyivWWpvtMxvyZKA+ecbmTGZVJ4Lg3mtkIn0+SeEDbjs6J5lKqPL2y4kJ5betpDorDQ4+8P4
GUs31/sYMYMJTfpUhY512zxGrLdgkvLln9AnPq+KpMacNnEgNfZScWt41mu+GqDAaveD0hwJSgOO
IlmIWG043Lh5uWKkpF938IHaL3KyeIi+N5aHWNhakZVmH3NGQix1mAIX/LD7w90YuW8Qd+0xl/tI
CJP6fWBKM42Hhg59I0cSaQ186dGVcXMz5/lZSaD3gOF+UZxK8kaCG2SLeGO/ArTTyQ5QIGXWlWFJ
AV8WL5ruu6iAQEpUN/vzWAdJ2/x/F9eCMrlLulRk2+yRHHLnZd8WY5pWy3cbUHr7ODewEZUwCJ9f
GKtOhsaJMsl7yVdhyKIhqStYQkaxs3Iz9BitoR3r+4Y0yjXITPPbfocCptIF2OlYUdsyAJW0+XpN
MQXSapVjVXPHual4eLZjbjZJOJlEntzJouxpVt4+tZX8AtAZKYYQh02oCqZq/m/nYZaYsTbivyas
KM7tmH0PsuK4xDEWlZX5SCrDoNk5hLe+CtDEpIHx4KWO93KQVejNpKNZ6v1aYVhSHxYL0BJQ/FNP
JfkBdkr0lmnLUvLq7MELHEHPymRFdwWAfznF78R0F7L5aG6G10GH94bbKRNY/UBR1/qt/ZyM+auH
Xf2h+5GY0P4C+hzzflFr0vIXEFmWWIza90umeZwyflZmeSECSFK0lYDXmfXffMNdJRQDHpn6BPSi
rM/cSzNcG9BH4qTtfE748Y6dDDUVeVzvF2H3qQ2UFHjF/XO+1QRtieG/pA24ZVH3T0Mf82fX93Sl
KRFcKODjeuoh/K7MtGdbcy7YumC3VHsVRVmd5TpAnw/DJF9QZeH6EUQuiHKaLU6hlgyP85MfCXD3
zgjMLCJP8tf7Q7gjZAcUZlPfjq3Qp7YBBMeukf34IfebWe74jls8wta1bbjd2VSg2HyDeRx/OIWc
cxgz4tYPuqgxpfJu3sJothTdlkc1CkAaepWTgEfNXTR7QZn8etw7qRTo8iP2Gp9284p25eV7xbs4
5/slgSFK0jeTdKziE83f7cQ4tK8+crY/m87+Xpt2RkH1++VMqFKKQZOdtN00S/oVASjU2nv01e0o
hl1N9VI0/uzkzBrO5EImbH2LQkOeHrBkhT4vGNZdFMImIGYb50oNuaU7mb+qBnZhFv38CdI+V94V
BztvAl1tVxa01Jn4p1y6p+Mohsvh7cmavBPxAw8M4A5GWMgo4e11k3T/PpLky/AvY1/J7mno69NL
++OfowwpJlOP7xaMaVUN6juqzw1H3eeAkvemWoDCal+9g3zyz/hvTYiQSc0GtJ/47F0o3YiRSvrR
rw4uNU5tiWLgTWEYYRqPKkV4lsSoOOZOQTluNKXzce9LKCkwHunAuwJ7fZZZ/XaaSuFoZXmf+LO7
WJk4JMmiDaY2fyr4l8E7cDgu/by0ngNCytN/V8zOwZ48FumPHtKlYhTpIgto1ej/Keqd59j0Vyj0
jeT5TxQab/7gLDaSWPnD2Mos7PQ80CbACw6nl4jBZhidc+2bIdCxoqjMvODH0ledXkS2JG0ht6sb
Sn4CvK+CdsIZ0FlzEyG4WqubGE0As2jaVjbPe1uxRZO1B1DXvvhKJLVbeDsq4cjK6EkmmXjTjN97
H17BMgD+Q8uw8Dx8UOnZeTYR5gUnKJibg6SeE0RgrdEPPQrJ8CFXE7oP3CKgWxS82TVisQrSmDb1
EYQ9Qx79sLi9Yheuh6CJ7pid2kGepozOIf8RUvX17R168rJU018G9ZoLAMofb/6nvixlrVdKVNDG
K2E80YUtdO9EQydr/z3xTt2sxE3pUre9iQlJlsShFnlauJM8g634gT3BYgI1iM8JwSmlChJpl63/
EWM1x9S+UeCP4tH17+IbC6xTfvhOncLTFCrHNZwGJJJmoXbz1obMtI8rEuaLI0l5Da2rpmvI7js0
cEWR/YlLsksDr4Qpbr7Mf9PMqdg6dodP6vJQ4fAlDXx0e5EYcQCTedzbfrce7TQyV487eGYR1Q2D
/9Q67GwJt7aiRi8sKIb1QYj2hSXBW28W4BJbNO2Mg7N8rD8ibmJta+ZogiqDiQQjIK1tqe5XQ7ZV
wDGdXbX4bwWAJewzL5mXsm9ijoQySvMTRuThttEZBngemjCVSXcxLzM5G8zvKWcmb33eVa0KVSFy
pxXqOyK+qWnlgBFBRyL8SMOm3+iGjEDC6icdVpwN4AhE7Hj95tFQEj8H5/0PHEVmyReHsTvuKCvY
Mz/8UlRjWzL2CcKfGd2Vw/0fneF8Sdisd8JXj72WlNG7SNSp27ktS7hq/PNFyu5kOZge5k9+jExy
aOgVPB6JgVUWb4FhTM4gK35LOdrCHIc92TRPKT2SJ7E9A3ubKNeXksJSDVApl+4BnB+K0rFH3xKK
5s/f/wtoJzb25PTPVJdf85R28o0DGhIf4BE9C3nKgN5Hr9crcEFmaai6jVIdEhaDkNGfeZ0R6e41
eNLMCqg0YF7D85jAdutnGQ57wg0mxR85i2zwO5CoQsTJygdS/YPrP8EJ1cng65akLYaxRFv4iq0Z
zSLU3hmBWd+gPKLoRn8RDmupZEqepOb2y80d13r0cFXqYiJXk3W/CkkeNhGYxWm1rXrZtr52Zj9J
gaK8yryS9haEto+pXg+JMCsKVQO0jb4SrA+CyVjLqkcC2bC7X7bvB6Xr0Nvens1h9EACXPdxIIw5
ieVItDJEbTFnhl0mvDLjQejELtd7i+5dGsMSy3249V/CIylxLp72DXA60r/aZa6zNqnADkVI9MIK
SAfjhf5hCrPzbc1YI/RUYfZR+fDbC2GXL9glJLiu860f5pjsVLXj/8IflHIynZcStpsZZYDphT+M
Mb+ESkgN0kxKtNOqy7RaqKEBHiGBniZgTlawTPCdvp0iZCuAeeTpej7u0fR1tp4az/G2L8+L49X8
KkM+tnWRh69a0KNCHjkKUP3fcvFFbNcRbfdU3WcQurRJkycsouQ4gCR44hLaLAuahKNtETqB+MFW
/BVv41KN2TL+BTPak5jRPLL6ID3dMQLKBKl14LsSjLVJv79SCPdrwMuS6JToqMfUCuHs8Q/rkpsV
czQLThF2/64H0q9Bgbk2scMA1sZqEVgLrQWZ+Qx3wePHg52hO43oC2QNr4Q41fLfxQUc9zkOWBmz
GJQSFQvzd7YpFTuTE3CMqdnl2zLq7VUO4/JxnyKhL3ZNnE7J2mAV6FBEpDR7vOEpF/HehUq137Gq
hsX3XClfhzHE7bsUezI/Ka3w+t3Txkusr4AwHUKXYSewHThqHHJ8Sk4xWznmAfW5CbstBFTTpZkI
qQ357JbMfDUoUYw8AA6omL49d8SvLZAjmrklREG+fdqpsc2vv5YRPVn+48NQjkmccJ2dJHY/mzbf
TxxEl5D+UL89MayB3mksn4N2IGXJO8aZYFbVn17z41Dl6RZFXt0boMHyw/e0M1mq0c6524qhupiu
i+WrBcVyHRe9sDKEY36k7s14656ZwcSs1t7Koh/A1HECKGyJe/2AN51gWwUGZuWlCI++pzQg7J53
F8+ReSIrJm7CvCc96LXjFmjJY6FeO7RFlJfLMlmOlm2gzBJu65eZ8LZkj8E+FO/J4p558RyaSMA/
qt4ME3FpNena7IaGnJGtb3+jKOYjfeBpwpnuL1+mRRP9ENlPCflJrwdq/OqMDlXNXchyBdwa758p
TNCPPc+3oTJ4vhJt7Hu20AhK+d83BLm3mb01tgbQUeiS00b3l2TlAXchWt3SFVMwOT4RndY4iP0B
p6JfzKjoOJG+GBmk2WMrtes/ZXxrHcun5UDGrkU2Txnp4iGYQ3A3FoqbBsREOTfbaQ4sjOTj+j/H
7SRrjEo12eynU7qaXEkm1gxyYY8QyB4JKhzA0KVpZCTi+jpcKgRDreabbJIb5qhIyj1AgcV5RD9J
5nGkkGbkiErhBhA7G71QVv4C3MrdgmKCE9l85LSIlLxdGPRa7hvvcaHDdGzqT5GrxRrOiOch5IGn
xgZlYRzBoipncW6WfInvY+nG5T5rjaZmdUZDZz2seNCb+/N6EJfu/1Dt1SvnfLg7LgTH7hLVZWBV
Pwe0ImAy9apXPZ6eJx4iJ08ozCEW8qmIF34w/IgDHaqk+VYseARH2BBGbiPuq2fM9laI6U5Kzy2f
59Wh0huWpyjJC9T0MlzhOb/OB0mOtbAd36jqYxt8EpmrnGQ5ZNlShssRg7K9ElP5oumY1MAdoLIT
s+zRFC+hK2PaUrtJtSryoRb3+2TvyAO4tLRY8SJsjlpz/1n0Vlg7Rb4i+oxnB4ZoKe06MIio78Cg
5afZUAHA9BxH3RAbWSQJZ8GDpwFvf16djsPZ9pc2KawTWj/msIE7gKWUHxFWWdyR3aSFtTmBvoWL
/j/sthZxh/U41jW8NdchoMLbc/x6Gr8xxwNH3Zch+z6tujHIqrEsP7Eg00Eom2EDpvB/ww9gU7Cr
5LF66KJfrwr2fjVOu7ZVwCZpyT4yJ2p04ItGsHSO1TohzdYcHIiHv3Ceb+0pUZwhWwlOF3x46Xir
11t57CllZdI6C+OmnSCPsHCYhVqbivpJHwUxI0xBJejm/goGZHrR6sxf+KnRLKKeXj2az1vhvAIy
AcX2NrDRoXLI02bDbrCAqy2Nb0kOiUNLJE9qezmsgb8fWipERqVZkb+Jbqn+fDLvdd2SIh6K3+80
4oZHn1C9JGI8fWJAm9YsfmNdsRkjwnRHKohmI+oAsCEOpIadLFd9c/s7neJKIGkDRsJZLb5cWhd9
u85SRIVt968hYGCh47SOJsIg62VkObyNA2C7MUgVQp0hcVvea2QwCOnPEl2v1hcSeVYuwvh/zAXT
GNB6chD0Fsk4hsSRChReKZkPrt9G9gTXN6tjL4kCZoMHd0DNo+ApDwa37X1KM2NXVxfF7vXW2iJh
g7ToqpUvZ0nrqqaPg+VAzimdx24JuF+wv7ESUFRZyuFejjgiTqevmQZMcdBjxlv64Dw+QK+huFKR
KWNymxJr06kgB+XRVrh5x07bQha/s8dOvyoguIk+BGS2v/dbqxDw5nYX/PaGieOBkIOkBwgNWbWl
DpO0OuGw5sOoxrp6Os6T4DoojReagXVf9v7ndyOGJE44CYUsInR6p0lg7QTNx+XX0hSUdA4dbZC+
cZavHYIGAciX4tZxyogo4rimR6ZXQB70dGd3+zDnEVuRYkZ4WtFHFqU6JFB+DsUjZ2vHDLJEp7B1
bNn0qp2vOz1e7k9L8R30bHnbwd+wfkFnECP2gV1ljfAV9fLGgTf5ntUW3gTXkz8VgF6+GqqZGz8N
aXWqnd8JzwPAxq06npandWJLtgaBpL82qfTO1+huXMos102zntoLv5uQxh6L3u0w9m86RrSAIGOP
C3tlxts0pxUKABXNaQQ6JLnWQ5dh+8iCF7GR94tCSqJcHHKBkhrDHLlcL3u9lI8jWk2oGLBRAaG5
SQttMLhMulTTHboN6DjNxxDo6Q1z85nbo+eDCdB12BIDSVlkT+C27XT/P3bReR4hii4YT7T4cxZP
ziixwac7otggv2tRis10fg6H2r/K8NUsUUgO3EGVPdPu8W7saBb8T+V48e95aEO8a2yNXiJo5gQ3
M0gNPOHvN7VNx8rwt2m2RYz9hIiSb0VVI1GSwNyW2Qfl5i8pidDz9PgEnyF0gwvMXgedeQr257BF
7cxl6O0GGqSEPDNQbwU9rsP8WzVPc03x16TlTlLXGiEnGcvvgDl76dpekATW9yAi68RVRNxPCVpj
89RdipI4WYAACkDRvXgdWqQphR0WkkbsmZ+YxXxuXKsE6cnCC+YYHhE2TG+nDCCZTAKli3AuPdn+
QLHyJvKAdC/QTUqbS19Kx2UIbfDj2q0liz3Olcw/lboybAEXzhURh02PVrZAzKy4qc5oACJHZV7x
6tpMETmV8EwUkPo38TkV12MDKsC56bOCVSoDepJ8FDh+HjsTYJdNdOvM8VOdFh61ZH1AxL/ZOKN7
EWsKgBTNSr2teYyLTcRKDv4zzwOB1sP7JV7cMgE6E1jBz/gAc4aDuO5IlFfu0CYwNTL9j8BOMPCE
BlFA4trBNoMe1LGZC2IvS81T4kUnKQpT8fPho7lVS0gPGw5X1kezEPDsnpmXThubEM8RyaX0OmOy
htZoEPhaPwQ80RicKUfh+ZqYZU7o4vQ7GuLbgtmej6UL1/OyS7lS/6x6o2Eb921GYgvZzxZ3b2oT
IiJgp7V7An4+yoUA/iHqsoCAmwYHKYMuml2LAcsCXsdVdychdCrTSw36zB9ykD1cho32GQwMygY/
rJLIuybUd37LLc0BZZ2nsGg7tI5QC+TRVNWpvdo08rO5YbPSXF/8+8SUBDHGuv/0raqTQwRB9Z7u
clQ1mGLCxIGtl+/jKeX8kA0HLj/2GPESbspiVhCzzB4wr6zixbG770c3ui64viqFNS9yYPGq5o/O
1jO+eua8U/eBr+0LcwsKaaHbvNXJ3opJfXVOMyL/0Fq1JxydMGl/8X8ltPgG9gLkwW1/lsF4Gt4D
pT6jBLc6idHVmfiJDPUAA9+NHrCINMpLJ3RFBVHs8OEHw27GEqIb6zd5KZo/7i1uGvgZJIFWdFe3
glVovbIcyhFGyqq22SwRMK8mR8STdFafEXU1uE940tHBHPp9aIZUIlC2pVjKo7SyTlwJe88WaLqx
R4XwG6ld5MXTydGnRh9PIrvDxK7s7Y+aDNUraQPWgCx8VEKN03Lyo7FBbbw2fdOUiHPGKGR/c5FD
9FjrmnD6nZ5UgJXgKSzrCNk6YT57i0lr4vPbul8/xeeTArlFlTS8Y22G11XmI3LXRMEc6FQjRYXv
QVIFsJlY0UWtmt+uo4yP0qgBhm9nJUvcmBnhDfuMIh6dMargtN+jLWsONtmb/YFJiSBmHKc3c0pJ
V7HdzXYN1lsIYTqWV3NN2HP7QLaKBw7x3TmA7lHYdHtj5BgEhbsOt2jyaBeHqEjdPuaeMey8zuWs
+VfPkewcV+rprJVUClNM9BpkHgy5e3jdb2IOX1Xtbzujvc1I/UwcZA08YEEoF9S0maW8MDvxo/Xd
pmfauNmAa73k6OT7/tpgXTb9wM5FAZE5f6PuXcdgtIEFr9lHtZ7drB+Qbw7mFwmW76sth6wInKs7
vpWY6FpDfl2iXV8KyKPHJfMhr+0ZiS5E79xspVKK4SqHYjoLyyzOhoo0nJhVb5Gue+2AiW2hpytX
1BESWmmTT9HMuqev+iiFjUPYG6MDsLMppLwdqC5Lu5CJMw0SnLKaR0MdHUC64puStqX5MiOcphoL
O2F0acEbXLdzyL9o9eP1rhWK9V9I968JVvfRc3jjjWECKBgy13Vq8hNUAw4PT22ideqp1stAHawV
BPhbPh9IjUtOo2dqaHr7bESpsG6BGX7W8UfuVrTwyeixQzWA2INfnpBPNcK0GlUzwmMtpRfkO6oK
2dh9GNVRRL9LIsx1c2w0xOrjYZiwV3xp7oQbVblywZsYKk8oXAbv3eXPFHfmMyo4sRC5wIDX/alV
Fr67Hg1XPl7cnXD7ReLl/xhOcqzhvQvnYKek4qY1z62Zn6lGEe/okWZUgY9+GFt03aRr6HRe9ZTc
Z9x2RQUrZgjxSviOsG/8hfw9QD5c9BrvG1dxeZ7m8i5Istv3vGlG4fkr7uM5T06wAuC+KbB2lTh9
wYINxOmUDX5S7hrLya6Dky3GuALRncAyGtkX/Wo5cVbdG9x78vXAMMwtnbK8/xt4cK5v6D6/2F/X
dedRmmdWeJR8iY2WA2PPzWEqunyMhdsaEsupRcCKNbKMFSism81btbxS7rfNpqOo+tcqaoUp6JAy
Y6yC5pDr/c7Ck7j4KyQdJdrdOf1eSYbGv4VOwb8MqRz01zAK5TBlF1cK9eH3Kbiy+fjOTmEU3M2n
VUrclTvKcXTgxPGV7mO9/G1KDKKdpVGyaELv053QRVlDMeWYL7bncNV+ceAjWFrPoI+FlVe+XoUg
2J4r4CIm8ncptayOJwXmS2aO59GfJMm64ep4hhbDOFrCoXIMjzxSoEnU/tTX532OsXR+sgrL4rKB
X0yiqO1X1zNaHrUX26uS+lKEtwjENHU+zfiSnvv4iSBzG9edpJtyv1xRYzjY5dTEvaGKq1mGSKou
e2aFV7aDf613cEsyGaV73upAva/w5CERsyLP8TuFku5LbSzdpaVuSuN9L9RIlFv9ExOPgJgR0jC5
b3Y6is0Renocbh8bsU12XX8gGnJH6UtVb8POBmjZlmuh5fNbyclLNKwD6E4vWuQldCVfNs/DOvOj
+clKMXhRL+b7zHWiOX24ZeK/qJMBkTD6VRzLIacvao3JXFdS792Qiipt3SKcn6wo1692kRRVJhkq
gWNdMi0uEoBxHxwikuVRfEwhbpwQizp44IYJT3x2an+nehDVnnl0hArugKUhQX82+eURrxnbkSjS
NPQMgcjjSREN3cDhypKuaV8KjI4JeuYy9K5NV8L7qwyQDmHUA2FNVPx1XuM8YiShHscARXTtyHVT
kJ+EOxBr/mgGnuP3pOo/ZeLR8g6UH+1Vt3h80F1sW/kEX2dENk2UQ0ZEZsvqdv7kw/35QxlgX/9R
mvTPHYQyzSDGpJgBbun/0bVaLYdXlz6zTE8R5Y0d18p+w0kF4O+Sl1YOh1yTLknofZCi4F6sHzoZ
JuQNBl2lFjnn2CIFiFlmCcPmpS4lC5k75z3Q9xnrohEPIPdWEXhe09jyfLgjsMLigpNnRlB7f1Ub
2PHopWU3hl0yEoAqy2w5seqcfFrfCL19IgSyn9svtEHlFDfrVv+PRqBz+WsJHShNpq3XWODdYUhu
riJmuivD2ypMVg/39gPedolBYSdyy4dx38n/xer9oEJbSkiSG8MvZvhpuOUGpGnDfEfbluD31UxN
0XCHmZcyWHHKc/Ejy97ZQofsouAhtrAyl+LifEe1qlHPdUNsoCshuWVvSMN5gSyeo+WQZD63Rukz
iJOp0fcmGGjSxAZQAf9aw0Qm4I2aYUTXmhZJhAvfrjZYuHJJOTO1sKyQZ5PbNsY7EC6bYDq75C07
il3uDTqtH7ZwEG35xHikey6h62dHiFJ3A7ckXiQqhsZ0CMDUlph5l6lgnlo2LodJmL/0WlfVJi1x
N6dj5a3qdHD4Jxz5zSOMCL7kO8595bpFgHcRzqThPDwiHp78YdADvL0FfqNCCH6L74iJ1McJVqF0
sHWAAz5Vep4LG62vr1XU71g2vTbfZlCSWQYyUpd6yeD4BFxFrWTr/draUltopkNTLxZyy12mcCV3
lQGvpI5R/eX/ww0ZktWD+KugrEx/0wbKkENWs2/TThRtNpTN9M7cD85arMdLGO5njkwT2kYbGFY0
6hm4rIVPWsMo6WmlweVR8OFjvHmFWREtor9dsta9SpTxeH/KFbpGmXug3Df1YmEQ7vXDLZ1ZlXqp
Iy9jhZXMJ++pSVrTgz+ho7oymLiuvcU1jF1eJ6Gsqeloz4bTuwYCK2GXwTy0Aya3M3onXlH3sFO6
yNkPgamfEkDKYa/tL7aqhTq23GMb58sy0BfdV47Ni3rmsHApLyeqrmm7tbeaoD1JxwDQh/9HLluB
TFshug6Wn6F7lWzNKa1mQ2ysrNyV5A+SUpjxyRdob/rZYMO1eCgHY5OaxhjjaWuu6ZLsUXdYsh0J
pMIwmX1n0MoIzgEM4l61yTXNglFVTGuJzXkftmSsOGoXWoIpiBLaB3f7GlCV33/Yt3HTMeddr3mL
UPh+Vfd2lOS75wr21u+2Y4m6y7p/LrfDYbFP7/x3nccv9nXb8e+cgJFElct28GnsF63AMrsXIC3Y
fRg2P/aT9D9/gsHq7JQ2bvC6oiPtA/74nPclOrJCOpcjcqnvcrPKJ/0t1bJch1sVTJHdarRiq/A4
bDZXthBvf0wIusyioGJGu6RsTDenN0FI69mW9wB2AJGLwukZME0RY5zUZlVbjkmxxMoRwfdWkqkZ
YIKV/3SqXi5r80j9A6+6iGJ3/ZQb1PPbVOGR64tUOmekHU9CsC1peRKsSK2A2Q0vydq+LFbXXWPC
gZLL6CXo/UkyinzBx1YHFYTQxm8pkMA268xM3x8huCVdknBhWYAcEPuL/1dQA4czt9ioJ7Vp7NCr
EMkE3iDm7T41dEJTy1vFGXR8Sxv2mUZmJr8kepO7hx+Vsd4pDFI85+VPl+/tJVPWcvZOsMz73lyU
1+FWo/zad3jLBUNECqe13xACxiigEqrJabAizZAWylfq+jQvAk38roEu5DCReKuX/2CKcPkRRQns
nvik/uxp1bQjJe5LZLe5zhwHCK1HDbL4CJiwRG1C7N0lPNiaAVreJ8jNo9fnjDKqr1qvPfz49QKS
ImIx2aP6whKsLQn9aXyYiVjr6pgn7UdhcjJDpcICXj4O6xvMoKCVjMAkMESTiSoUBQl4u5rBFjEw
zYs8resQjs71zcfglfPUwMqV13hWjx/WMkHcnTy7ByCi9mtgAX9gVmui8rOSe0p4pmAYyzHikOyf
xWXDMw3i0SeFIw8EvmanDHRE6OZAv+RK8RRP6pw/9mWaL5BG0kDUU3NEolimqCETVr4RPCpMFzE5
JW8Zp1hoICGEvOpVXNfVR9hTaGNDZ7IoNQV1sTfQCCNL49dJRUKwQnT7kpV9ADR5CrkaKqIlpstb
JnxH8IdxoWvcF52qyj3SvZc5Z/0uaAqXpKBue0ku9hV4XSV0c31c7V3N1rgZmQdTtizy8p+Xn2vu
srseQ2MUAwWfa8laFH084ZFpR7gQXW13x6LO+YfH9pN1+NyJyOgzOKcKZlXM+owfI/P+Z9zHrnV8
E61ffYZdCL+DzKbv1R2r1LafjXClF7f1pjC0N1cAuJe6eHjAbCG8KignJa3zbjo70zVhI7HkYChq
X+t/d/zCvXZ7ggeE0sHK2RP0oV7lzzKBx9O9m0imY3KoEbRKovonjGmZQAtA2q7fmA+rVdsShWnk
GVcsSkOqVv43YMCUv7ViWrMKgVfhzdyl+Gi9rh8oWVGzcNoLGvfNQd/nqAoxKmlxkHYKCTmT5d5S
vtyILgroS2yoEyVYdbFra9Vd5QPNr9ZPkefMTdKZKGDxclbks+aBAyCpw3kbYxOGqYA3n84XFA0s
Pz/YYrEO92CkY+wwDY4mqdS6PrEjblasswiBQstnWW1aCpodEmUWWYFGMZpNwMeKsPbOOfS8cF7H
VKyJnNa9khCnuYn7s9HLneEnXaHRBtArGuYjwHPlsCmdOUQYPvAmojW4kgBCthwFnmVkjCyIK2pk
dKNLx/mh6W8jnBGUJLFmIacD/5aJPHvDXsSrfiQ5AiJvc5Of+3dbmwv3V8qxY/AWfHgnKlsShTC0
XDlM00r/bWoIyh6PAxOWNPl4lWyHY0baQMximH9b+M6oOEVOp4yDlyiFoZEtPfYcSQt5oH57iSp0
BvChKINc6/I0mr2zfq7rsPe0Dx/OcHgWhGzbL1KKS6WFcoUhInhRXf2wG9t9xH6yG3vvG4SgHwku
6d1L1iWf3hnXKRmkUEIzpj1rZfUnV4FDOGgajxTnIyFb6jIU/gxYmeQqMbP/IVj2ssSFVIqSs49q
X+xPqUuyggbUtBvv8+0xMuHVd2EW3hUSAmlz8Dtha0M2aN/WHyIjBfqgU24H1xQesh3LKA9BuCSt
Gb7pYaZUknX35+6Yx7h4cMjgHyETIbjw+qFXy3s/T4CdBu4kXBhh8Ssik2mqVtWV2TSOhttCMbDF
E30vqQA79dnzBVQ8cjWtcLleuiv40QthCfbdVwZAFDxY7SNYoAP8stHBnA70WpYes9LhmAQN25X2
j9hmgpt5YfDXJiLkK+pllYbB6IVjyQQ/Cb2XIK2N9C3M50Z5quok+uIYK+VtSlnBr2or+ASMMj+6
EFv7Zb/1zq/HWz1ZbXNZkbcUDR8ag0uX55opEru4r/uiu73Yb7RgOpZkmg0g2AKubGesKoYvabfY
q1DN8PLN2Uq0ZnixsWd27dT0Z+XEvcNcRRCPt5OZK7RyMgwaNhhZBVtxfO3qEQJP8nzHFshlsS/Q
/O4dLNF4ddGduYu0CyWH2UGReN/mqhY/+D8dIxUFNWdm1p94R4222/fNYGVWI22Qhkh6aYaA2NxU
F2Krvkg8FvxRrrbZbZ3HKyrszd1YmcM9AVS4JGXc+r2arm4fCub95T31ckYX+3tOHgSDxQpAdJle
rBCHJ1sBSWQZgh2oGav+0jm/bpXVCeAohx5K7wArkycy+QoXKCyirCKerRRe+KupRLyXSKPKBTzc
zeE6C6DvQdezs0UoTRrEqyUjGb4DJ3op8RqpABZNWkCofYDnLsvyywby1qd3IgrhnoHKw8oriyiF
Y9ksqOGrIelKwc/iEIcHwD0g/4s1IRn2yob8OvQKLioRM9vf/UZGojXNSGow0tBSFU9aO1dz0v64
EKMU6LPtZMpXmFpkrJRBuEg2t6onXMecDJ41ReKrFJsgZI7/62M83QpUIwwwr7wJbo9UO1zbdnmn
I98PSeYb01owCeM46t1visAs7Vr/AjdJD+M4f7dXttVYhfKEKlqyqNcbVVVhzJWnp518b5l7iQl5
pnrEO1zCfr2COGc4r07TgNaPkW1JGc07uDs+ENhEkQ/pQP4OUxWFReFSYn299WyHJBtx4KxgGF2Z
VIlojSxDTm26MqaRFXyVsvfYUXIrpqooe2vAXAc666NfaGURZSyYBlO5dBE+HLSrQDGodvTVgvTn
GS6LCaS1QKl/QcmbyX1vNQ2aTLlGpNqdJcMHGZ2ZcrVZjhvy3vAP12gICMZ7wA51bq6XOsn9S2RX
XfsR640a0D9bOiFfYYDrfDYjZG+nlGuS5K6YbUXFyp57kxQUwN02lsAb4TAOwM5XILHPJcLkQ0Vt
iSFHqe6AQ3XwE0FU9IQEVIk6PV3eYoC+i1e4OZA5UqF76JasHXIUYwYWBnOc7RLIEcwEq4QyEfcF
ll6iXEp9tVqrN+0Pooybpe4yktQuZn1vWvnOh41p6goKCx+9F+kabeM0NQZNTvYrxet2HEG7CnvR
cm5n7CGBx5Ts9p1h//K5bYDDzH1guOZF1VIH3vZMcSWX0r1n2fslozDtrqVIA4qrX82Bae8ycqi3
VxBmVoy6IbQUR+PoxsIg/t/wbGYarr17rLsEXfRmWWyNqitI72EeqboSUqNupX22boFygvvNsXjV
Rdew9wp3p1eMgrYEwkXCuzL8WtNvTyFzh36YJ9EI7RXWIK9ZTGM8/HzTddfcZhTcFcfz9jbtfD9Z
r0HwdNbpFeP0acUePFEVzuuGyN5mXLzlaHe0Agy2DJmTko55gdfgcYqC8MIsaAykvETgqUagei0y
L0z3mjDdl2Pd+bdKbYUTlSy4I3S0ujCxgCXjqRQK0dbPexg6ztsqUfOntgg2EzIBEbByLyXJA9Ky
rE+tkY87xJXoAhdaNxjdmnZa4TSwusKqMNFdQ+MZd7wjmEMyu56hgKsdUVAWn8dg8lBTRRl4/edt
aTYY7dzBc5g1Klb6MwEiizUVK2WQ7ujhmG4ty9RKA8RaXr6tKrT60nopGLwWD3VEmFCip0f4Gtz1
PZLbGWmNWMcw9+p5yAbXHc2oUKbUEgK2izybh4Ulu1Xtno32IbQ//qa3xQNxo5uUoSryRRKi2iby
ibTghAeQt73rAxdbqwrpVTeCx4ve/Bx7pHcbqKHSaNVIoN/YNp3FXS9XkdpuZ3iNo5n2i90SY4Ar
F3DtZTmacBmOgXmHMw5B+LooMr9rXPjzq600Fc8l04Q1zfD5g4lP03cTBSRkaQtagD49w/fINJSu
nMTZI3AXoOQv22FsSnxBRc9CIYiVl1e0nMCoi6ydleGjWJnJ/vmcN9VIYWp2t87n2jTjQMoV15OM
RnnnA+KT8Q+B4RdN0xZkDaRDEeDeg9MwcWz75qEDwq/VM596F/SSNFTdiQUei7/3Of2n3JpYR2yI
Arhx9l3S9T1x2gaWXrXOmDCUMX8UrtmHyP4bmnKlkLgP6Jac7lI3B5byrew4beu3Iy362g7Ne6PE
5CrpyH/ZHR6Bgcdhpxs0TrRwiWdVG1jQJiQBFEnvP8u3g1rZqnvXUngDBOeS4ay8xjpIHsfH6T9N
ZaXEKzs/b94Vg+h3AMGNWBkRERxDR2etm6Ot86iN9chxwh4lsFVD3oLA2CTGqjVYP7GuxMNws3Fe
VNUKoNaJ1BpGVv1v/wFgjG5KgH8zI62LcHF8mIshTQoSEGf61AvlyrdhAoIOaysH0r/V5JjB2L69
+m9Ycc7/LlOr0Hp6lcdD0DZwdysODk0YD7v/MK3TjAMPzE/SeB84i9x14xVilZ5vwcopNlpx/4yb
8JmExTDk8yBJ6FYjCUpUcT11PaipL8RzhJkVp+NtMTWzPSv5MS/alxfM3E8awlE1srDPqH9rgeJj
pgTR3a2BQh8WudSxwCMOD9+T7dIu0LNwvePFbTFoASx1GQd3rR/X7nA21peXCF1fohRS6bz1UfCU
qgKdDPykpI4ypAJDriuOXzggNSTSz1/YHX4YXljPzBYi5QNcbsPr2AIIIWMP4i4JEE3L2O8twUjc
RHMNbTA3VpV6zDtPwb3b3i7nYP2ROkPKzeJrq5uwGjZBv/Ca/ORjP5znkVjV/FzihFPCfmVwPHgJ
Wc4e1m1HDFF9rZK+N8VCRa2q4/rP+m4lOdNK3/CcaCxU2f5Gl2McR5iuZHYMFvNQUSKpWjwUwjVl
zZr/cHIkOc9Py+9fL5kFOONAs/qLn+d1NS0faezvbE8F3rv5umIunaOACweoK8hwLkQYSiW9F5Ub
NSdksnZJKn5EvSS8GyGI9N+p+TkxkQAlkdYtHv827SfhbGzHe4cshytP50GlliEIUsseIbntZZBL
2Od7AfeGAjOSwjAyHqhpzcDyN6kwWxkz4IKLZq8dAK1SR40JqSMqJwreJKJzJf3Ykw820mZ0e70+
DVIDXIpum6kyTWrwwvF+IsXBDAoOcfLlFUX80R/tDS9xigvC6t0/bFeuZNF2LtZKqLFWrNVeR1eq
txDvTApnAA0uVujxU1O3WjshNSlz20FmiJWjHuwIRJ/cvrlHZwldNxMcZODTbNozPLmgDb8BKNo/
aFJFrpuL3VGoK42X8/bWtWpbnScb7u4kcNnQzjHwN4Tqi9mdlUn1vUliTDTrjcjkl9wvVDiyIW1F
vHWmXVjw3SEJyuUfFHE2Zgb2AC3RCKz9mE5Cc4HqmW4z0wEOA019tznWVXhmwUbvGEW5tuWbNZs5
7q4iXqUJ7siBgKDVJr6kIQSLSTueroIKXYkL5SuLaW9g8k8rUPRZ4/Igdfdh0FbayMQHEOb+ad8N
LKdEvAdpaag/TCL8y7fTdPO5YJiplL6iEAIO0C5W892+XMYCvCvDeuLj3EBKxl/prpT+J23OKgp3
dPRE9qAWBfVuQJa3p/gD9M3Bo8PLA6u4AtmwW/kPYNvAHc+BSoGyeNo3B6tHFGFoh+4iilZTmfQR
ACmGNtzLQMFg0FRsFoohgtskTCP2x4wNwm+ygIxs8K8S6mcLAJr05RFk/CkAJnmKeNR+5fsZZSfn
ZxKUGXgLOQzqf5OIeAYkOxb4Y1zohD5E6iMIgpqeXY2OW/3JAyJWLRD6hPuerPsADv3jIphddXVz
xyH2k1OUPFgsCsawqfcWhHEg+6YXk22n4NP08soqwsXRcyPLGLyVTicm1C+rqjIcTkWQaBMzQExk
i9wzcEG9oLC5B68Ch73tNwDxROXBGe6hQB0r7CdwXuXLNP/qg5zfZEURPG4tFix6aDABac/cagqu
DVEJ6ltZYHGPw8m6Mk52r572Jkn8PyS3U2dvp7KZ/ZwsS6YS0dSu1PFpbh7N3H/wRWPwFls9KZ1y
ja7Xick7GagJ2rPuQr7whpkmxnPNRzB24Ql9vaAvJgVh+uvPRjl4C4oWt5oyecedhXHGnu0tE6li
SjA6tYezoy/TCoZjLJ2kuxuSvlFn2sk+WEUqagoZovprrljqyJUQD/Bc+2iYHJs0DIJiVgW5ecVJ
xoCqzrYOW83Z5vdUpTopsQeo4fKlDyw6E1UpUydsodyGm9O7+TyvsKXjKLEHNNyyxxrUBmNMMS29
ab34OXGmYs6fE2hZE9sa/eknyu6CI0nBc0XZaK3yng1paqMReFLsiAk/uAWzzrAr2DBp7RooqXWU
Rgpmcde8+XYaqQUmiwTDSzuvjMO2PYNb6tiZRE6A6NCXs5g2Re5Ayd10QiDNoqZ8D4pGTVslelfz
r0N/rTkoL4VCh4bzGUluvPtBlCnUfdKmbk85RXCtNFejmgqvG9Vm1Qse1bl6S9VVCLSRilZig9Z8
p2OTDlZUVBIiGDBQHJXdT0NBKfUiMDfD49Sn/2lK2OPzoCaxG8TxT47B4kSPThw8o2FDZZ/AhHt9
xtbm9nwBrwZsQvzFEzZgTsu2FtVLuLcJJ+XAHmjpSKyiGumdpC5u3a9ka8ViulkP/YbHOlSyQnUW
TC46qPof4OLlQSbLYy9mUA5LrSZqpmL8rXBnmVRUKQOa3xY/lZK+ZjuFhh3D8XlHZltcUFfPxRkq
qWWJGQ2Lyr2KXzIZrMbi0TmRVOK3EZrhXmeKBlMIP9Ljf6LK/uV42x/vDnrsJmSHUN7qOsWYgtxv
rZY/EVnwBsBa50hDPcTtQ72P8LF/8SMti1I58Su32s5O7zQUCRF5IDPoTtPOmtY1O3SURN9EGcLs
G+o/IKymZptiDRO/m8B/Xt8dkxNdcgyqyFOXU4GuFM6+rYPlLaFKlxL7EysMATPtb3Pu/qFh7LOi
ov3cHmDGhYC91GWnv9c+g75vPuVt0l6m0Ea/cSreerLazg7tCXRj+GQusLUMGrKVzYdRp0ZGKe7w
jwsBT+Ms3SgB9j9cl15ZgoufjOtKbvW6YGQb6q0PluBQrD4MkFPVoHHz2BANKmEiWXFFEN+09u8E
Y4jPwttOo/YnOI65MqgINvLGZhAFaGzFtMxIPe6GUzyqWEXbJhWnoP2ZGyH5G07Phcg9811tB3g0
fk0phOniBgOGWACl6mUekk3/1At2rdqJHXDmO/PP+t+euQJfAf/A3Xd5woKXJrk7FBWYFXRDVlPk
O4PiF7RirTSfH45saHi3L2wxBG1splpUF/iUhnQ/9wBIMd2lGJB81rbXvD808NnlIHBbS3cjNgO7
zurpLkUyc2thvfckeSuu+BeKCOdXPHmtj3Xwez8u+Ta/bZXqTCNHnLdKh1VU0Gvpex3LTBiTX+wY
6nS9tHl+VKQxY8Ls0OlFBN3Pbs7nDwDI7xlUqmaFjdthNGSJu6mCyLWsPqmlSlCd0Eg+EYhG4Cc6
7wymAn4L29AwPmHQwmO7A7erI9AJFApVOuEfFQNvOQ1zY348hDiR1e3ly/OUN8o9wdCHFDtC/DdR
KOY+PKmLfkBzjEuCn9lMExRzcHRv8Rx8vbGoWJS3V4lj2D2T8af18Wo8VS0N3tTzUKCKie3T5107
qY1YmxNcz4KeX4ft3e/fdZeRCzVVbBfVfsmd1FFgVzRLrc34CFSGkETky7ihmWcPLQHTHQ+TlyjI
AKI8+0b7t4yqShGrRlJDkh2TnXJpgKHm6YQU1ZeVpdEh8Jux7F2iOKj+GboU3d761x5gt9iJwFVQ
fhtfPo/vgx3/WcnyNNQ+rvBgtqkmNBDtXE+DvZNPl66FtLwnMQXE8FdNc0h59i2EKQFm8Bqw6WKH
Q7wgPsztnCGj3tDOd6mpzsZNo0Cvm+gghOzl6Km03sRVmcKaXp4zIIHwDTB95TIHPY4BuEq8C+yv
mTtNh/JiHFYZd8Ld3oXc/hmBupVNzUOdkXCEb07hbc2qo5vLGp98n/0PYBtb2n3QV0kum8+YQ98v
UiZitgjKexvnsjRL/qyn1kbCFbHPKATt1fFxe7bZR7y0k2OpxIPZtbjy2Q2XQNMk2kJdU1/9iDHz
uwV9DxXJXfhshlM6euNE3pplKqGnawy7MjaVNkDCIp0BlgmLzB6GCxGhW8BteC95CzMqlakOw3m/
fz7RuzcPluvW8eUQIRvArUJoDdxcXYS47MRNLjmXDb0HcSr+9t8vkAiDGJxuDstKrFquj/8kVe34
QaS1svfEqN0NmjgccvNEIETHJA6kmv9/6dm4NgD9yBwZZvRXp3NlleaT5MwjaDNMUzIyozv7pKUJ
n89GoDou27o6nujWL8entClEgk7kt/Aw0gD+64FW93MXzBqvbTSbzmHWiRssOXz0RiU2/j891dxf
dnRYQKKXUZsd0OF0PJZRfR9u/CFNMvhksiCVcOeIeolpcz8RVpkRTbb4M3sw71fhnoJJzHZr/m6d
5/kwjAYnVGRoa/wvYjjmBEE1G1dy8bIKdVQeKVPAOAsTa+vODB1FlEZqFEfwz76ggJbMzhs0hD20
9TGA5iC6PGmxVa/FAivd1OLarlaKpX93Hf6kFuapF6jw/7LYJYZmtBlOZtYA+BYqjNq1a8g/J/8j
I/e9WG3r8JmbcYYLZOg/KNCxCrAdBSqNUHioWKXdKpCs/OLXz+u8Ohzj5jjdst8cx92RqMofZOKQ
7GPkv7ywmYLXD2sfmJmCnMqOknxqYxAYeed40owgTgEUP4Ulg3VdsIePZlNcajIzLy7u20Bgk109
MVp4ysQMBW+vY6BefFk3L8D1tdnnVHQws2iqUWS0J/8yHTKGDMdTOULU1mOr38kTMBjOVdXh5hyD
Cfq/gGrvhGIZWh6axzWCMX1MfWxs+jhZi1yFmJkG1WSiZ/s77ApGovU65xXF2ta31653z67Ginop
kmNjYnvDtpMEOwW2d5RSGP6HnZrRegi+nGfEGShf0KXR2VIHXrMzA7y7ncFXoMjMmCwkWYLMZPxH
DBYAyaSmEPcPlhhDDNbu+2P/XgW+KiOQRYzayFd7q9wvd6XvO6xqJg9a1oJPw+cAks239COgT6k9
4Rr+CAhcSN0YWi5bBDAvDITjX0B64SFeCqtt8gFdnu9C8tt3ix00C88iLFLLsUZcVHZJNbWg7xEB
OUV+J4+l/1Wxe8TuVqKcgIGCIWaZF+q5C2nS5BzecaUDSksG3i+14qDgu+HOF6DV/HJIDumdKe+h
dVvOTuWvir8o8Nz1PmQjDV79u0d6iIyQDhKyI8TWOBum8Vmvjjo1qNKihL/41G+rQpdtcHWW+TEe
kEWEhCq5oI2cKM7CNOXH0DnteQcRQ/0k3/862aX/+xPBPnyYEZEehYfLfpo6UpAyniG2H1FFmB6s
HuxxUwAu7gKOkAq5XHurYvCJqI8TTEJBOXQJYPVOBc2b7vHFu9YwQPfyMkZSlP5b8PGdA5YhnK5p
IuTtcOrgvg6bWikhF5BK3qRKpVKfgAzwIicO+UfUQeglfIcOIMM03vPPLBlwjdfyzACHT49MQsGk
g+GTII5/fcrEfhNq+bOEewALoTiH0hO8i6goGSCcEYwIVD+rVpHRJvOQj9i5OmaCZDHdYzZwNpse
LTsFyp3MS4v/d+RnGTYBITTGuQSrjprZ0Ly5whPRYChDZSSgXtpBxDkDYjr6EcON/JIThCF/848m
4+CtPKHGdMXN9s07jMBnbZXRocA/mZNBdilpEc6KAHXOkZWs8N+H4hHzY2KAXIXQ9G1kyNKNQQaq
LEZr+d0gaqSBhwr2CSryjU8q2IGtE0tdRkg6hmPxAHaob6MbyuRSKJv2gO/D6B2JLSjXDm2RDSum
ZLxXjrZQHV3U+Dn61sfd6fcyp6nn4cFZ/RtpWPskkRkhW2bMK2wrKjujuIOHDRGR8H3o4MICNkSb
pXuCKO0dt4hzNE7WGuRqjh+SsCTecDDPEe6ifqofApenrtoyuby/3do2J9UGgU9YpQOTyne0Wbj0
aeq+5olURtpH4qOEpZJs/mVCeumnpVMbngJsAZ6+DIId3HHPiZm36qL6mRuYOplxfQnUCIldHR8H
ZfizlYBCs2to3c3SFhl5440jVUZUywvdirxbk7jl9PskS4h77vOGS3oV5g3UkW2qePcC/8Mzvi35
qSEFegCWaIqtFOJIa0cK+ZKYMqMvicDzCb+saqmlyL0bX2M9NNkJkNhRndVkPoQ+6gqxGUBITiw1
e1nNOy3yuIOA3di8SHkn5mrY9Q1ppevVRm8Vrf+mtJNH5MA2dFNdIRtkiot/hwFvs8C5btqlvvuT
pe7gdLMxtp3Zixk7EeYFQFlx++gRCavxNjldHXCIFVqIFavCKvXyah+AAvyGTTj5n03Tkl4z2xsq
gfMcSdvfXfydltf5yRR3pfdQY25V80COJF8O+fAFw5hMzqFVrkvlFk9px5OH1nGllbebbetRz1ov
UDI9LBmZ0OiaK0YZu5+kjBeKPQ0vhx09QmCdvzoCgQtS6ryfnR49glf0Zhp9SxDKWDQrncj1RHUz
+fm5xJ4xkF1b3MzOMIgwUptOUWa32q4kIQMxmbScgu07idTE7jRy489EvY1VbMRc7GR3HRbZs5bR
dJECWAi1ZZy8kw3/zCHgN7RSqfByi16ES6ZsyIBNVbscJ5PUi3rrNt3s5mGbVInRJlo8cSs8vuVO
hkJPjD/6hMvIrYr7j5TDGeNG4PiBo1HxC6PzbIuWzOvKHuIvvippFbLjSStWQErCWMkrpV2EN/qA
WAKEq4r7JHF5hJCsB/g0dP6EAwWA5QIBuYO1f3IvH2XT0EiIbm6AhDunP2cEz8W1rmRYAe+F58JK
o0gfzDKjPrI1QU0OrWu92nBOYykYYVZaNZ+WsmgtEu0GJp9dkXrn9mf1XmvrPXQmNRL+vYVpDLt/
4QRXrW17dMLSNGpgpMQg6h4GHPjWDS6kWYxd/7prSBR+pGF+v7fd89syTaq234+v3O+cGuTaT00S
zfYgi86lZw+FP7NEcAgNpTCV+ygsog37jfH0XYEIN3WkVhDkuekbXXDko9I4VQX2KsGEZC4cg7A5
+hTISZacFKVxUbrFAOThhasZ4d1dwpiMOWH+p5Amw/yyySIx/ROZ9fFtM+wmpE34p2lYzvbBynMc
2vu2yOKaAqPR89B7WtmpMgbpfSxufNDHam6DAW6p3MEt1hw9YLB1Cas+PdRitpJhhgpGjhnrQJEX
6Gq53diZeFdA9mTiQ5qwnSZLPWpeZf6GE4UPwxlG4pwCxRhGxfmTUtsMaUaZQNmOe/RObilBvRxQ
RFR9royFou18XdYDALHxgMcC0cmCmk/PdnXgIYSCCT7u+nMrkNMd3t029MeNw7oAei5gkMg0ORQp
95CLPjiVNPiCAUa+7bJ0rcoxXrhv9fubd3hnhB+9IgYkEpuG8OunNzTK3e2GtZEteJQC/pgwRv7R
jd7yQoIbDH0Fwr0M9nPUETAQGr6aKfiS8bYlObr71X8sULNpf1kPEvbkLl4kKKr5glm1bAAgIho8
8TLEYB+T3gXrt0zRdmGyCk5mCY9sok6LygNXDZ7nluWnxhfE8SB0Gm156AuivXuxBy9FbW3Aum1Z
18ZBdcIJ6Nox/nF7oeUBOkNdw4x02omdQImyPVmlhLd3sl39j2Uv6UljnCQUVaZGb4EISwXw9h5c
Bwwv2WlyZ6yICzc7f5n8586dEIg/4xI3Pn5HhBhBh0bpyDRnNzJ9s5TGc+7OWIK2OwjDITXyTkPk
mAhuZ+GECNidJTortNAAsJMX4ShAcl9FuNEaVmn5YLZWy5wg/wFFYBFi1bAH8a4JSIyaQT4J8gJB
U4ECUGDohwDaqqTY3NDnS3PKTmQXmvOJcSvafCoEYgzLy7zydT6jjaMZnaM1ZhkGrrhSLVGacAPk
+f6wax2t436ABQRbInDtj7dV5FU/iHRLbxN2d9elklbvfNFoC73Ch2AkN/a21s+U0P+SVQRlaiX8
KtUqpiPF9HaiqsTrJU0dyx3A0hSvewdJIPu4oFPqRK2FAXR7zQfXbG+zW2jXgFsJX0jB6pCWLboZ
HUX5l3SDGer6no3/g83Ngph6IV1ORGpleAqZJszjd9i3AoYcpwtGV6Y34Wdfp5l5jUDqNwMJxAD/
CIhxygHFis0CjYYgQ8DXelFvmiM4I5okyeVbmYhjnwOQGpnCi7lC7DGKz2OmFOpeYvBqGFKgNUHw
3LI8q7BqMVCP2PePaLY+uxYjmC7/l4VDmAnKQIEooSe7bU4gnbNNkkDGYAiEsOMr9qoubD6G/V9R
P1avakE/JYtG5Ni/+8xObUWizhj7oWvrxn1ge514wi1llMtaC7m4Zs788FuLx1KKdKE7Jm2Mpc47
syIQ51gj2NT2qrFcYdGel5BLISCDPdSYSQhpYaPjaQp9TLHyuov/aV6r1GcG8DHvND/jKvC6xTV2
nu6voi0kuNBwEhHHddYWkNoWnADHef2cnfb4SyAE9Jyc6a9xqEIf7g9QsC3NG5hNWROlu0xg3LYM
HtMPWanhYkwZxVmLlk5qIxfukk+xjeHQeEixXVrVizNrjU9dVeRzYA4YFTl2Zf+x0yzUrWeooO4d
D92Q7s2GQsNY3geK/aurFoatm3/F3Ql1jGwi13lPumzayy68sF/ylJQ6p+XPpxVk5QDw8yIDmQZk
NMqHGDVpSuedcK/Fss+lSekaNI65IrPlzp9kkRKmI54pook5tuLMaZpLfVFNjno8fMwcsrBfGoNS
E6DYDE7feP0qQTVe64WVq/GtGOHopwjxq1Cc1A5VCYu2hdlMsN2zM+QgoxvOIy1C+uPyI2GMrjI0
gWYrBIAedj6FuhDJs/w7LiVJQL4ayc12BH6FbhVfA2MXaGg0uOIA2YU1eA6t6DKxpNvvyHZNAa3M
ozaOmbpDPjxG4mKKszbozr4vJrBN2vpvWfAUHaXVRdLk581Ju5RGx2KUszj5GyoLbWPgVSlAs1Yd
GvITa2AkcTsruYKTHDwZ3hOyZr9gbH3Jkgj/GnnssZvwB8hbT+0Y/83iWIBJJ5S9KdJeL00dmXqQ
fC6FwHOUkZy3Gwkh3ZlZMl2UWughM91C3ApugoIQ4usLeFt4IZKD5GcBl1DLWmXo1bBhFMfjqSaN
rqpbJUj0RuslOw0T6hgnJwhMDY7CGy9lR0ghrfjxW+YbsY2DkuLFRhKprNLSTjHOIRlH8h7eYjdr
Tx2hLZION83rR+eYGhAlYQX3jqEJ+mM3aePs2f3Q6sWKBwG4sfhdtvIQyuSiCAgoN8QIQLJYed1+
NraBbk2AEhXS5Has9lZMsPENmQewpxVnFNGMSJ/vkhs0hIg0oV6QeheATZd8Koqn8P35ZwPzZFYH
pVY20hjs1wADJuiYbfZIpbvX9DCYYtQ+1yt9X4QWwyEgvjLb7kX4ToiH8oIkc8vlHqC1G/LOiirM
nR4NizRlfrp+DQ2K30rWXxd1anV7y1gEEvNTNwmDIBf68yn4dvVmmBWWkAbAgnoa0UFM8arg1512
7uwq9PiX/Vn2XaXW6HA91MSF3T1eFXFRFNPoFMbyJ44YA7VCsQGuqWHYG1qpWa3L/TJ1heFWF+en
M3TL/8EpdY/ZeQs5ZLYcqqgYT4ssOVhGoRCBRVjhCls0m59qdlGY8aWTDq5ZzOWz7wSU+a2CYG3y
bpWXMEg0DO8rZmLVeH94Z+MU68ob+Ba1Gnga/oGgOIXu5OG9gqp7dClwgHu5CvUzItAbtzudaRXh
SRNegyT58mxALpgz1qsSXW9gKXK12f73WiwrgjMNfpwvHHSEKJDwMqbeomVJlTowEsil+/7LI9ua
XzhR0qlmVP4dahPD2hJ7FbF8F8cHm3qPhau2snpcM33NdDljzxrMhSFvkcsJrXN+eiGQSmNtguaY
rCKSAaYpFyNpiw9/N3d7HiY72AYq9ZLwpN5azcNNYTh+I1ukyHr0dRS0VSGG82iOu2mlsMKd2hSL
JxmucGmAQAu2Aow8WgKBoYmBQQQfvoOVyRqoLdjBan6vvXTBTUL34EYCneAsFvdEnij2wxx8CIh2
xqxLt107ZYLYUJyM+9T3R74fOW03+PALRny5bWOMZ/gDui3ZUbt+7i3YT8nW4+zu5BnsgN/o2gIR
IMaqjyiu1uhA6ngz3MToxaE7hoQXec2oN7/NsH1arc2GzRMYegEzzJnVSu5XiYtWmglCwnXX7pr1
6YPO6JqvmRx0+2OfcxrnbBg3jicJypLkdHTligkexmY1v00dqyhKgZIJaU82r4C52m34fZhKUIOF
gQXuvm8uTXHucRkvTxvE2JAySnd/9QR5HipP56PEWRiwa3YG2LqeY+OJEGgnABvHDQfRaJLKY4/e
IVgJMR8zVUGnwfethbexdJgKfJmYm1gcotLmNT/17M5agED58V7OQqI5ohQZxSIhxnOSHdg5RZ/7
KUa0X+DW9UdhESO0GXG5DOF/3yfvbzPdcQH7nzMKt9ARh8FBkJY9RanUyKS3/XTfqmDQJ4b8C+Ty
PVIia4siMgXV2LWBmmbn7mNgeA5FaGL1YfZAy7axF6QtVy3rl0Lcklqj39HNRFBT53ot0vdu5iz2
GE6qmvd7QbjZD9UgQtfSFgs/BP20MrU8EtIFdekzrXJ7rvJmiWBuvm9m6mtNlvum1ovl8MWDZG0Z
cRkr5Le98MvD0d/mMR28MkQIlqjKTPJZCUg3xaBC8efHrL3dIkyG25phrNxihziW2c8SW+p7Xut7
YH+uK7aPpZZpEcKS+Z32I993XyeZ64rgPKcYEEhHlpeRDTM8XoosLo09eHKF5UKpoVMpSxtSRBVR
pgiG7SP+99VnCnP8t3Jk3/CcMPNGjOP51ZvMcO2ykIcx2Af5/nIZMgVd34vrm9BeQGmNDeBYcIm3
ZD+Y2lJ/s/6JpNkRItLv6xVjKQx4ZScU0kJeNyi6/h0SIXiOaLLwjXtRmP8xQiOvgEgZnamU/xvM
suKem7Vfd7PuZBdgAJNNbfxhMrmBU4D2rMJ9BZoRWOFmeo7TB9TO7TVzK/xfgI1Lry//FmrgsAwF
xiIltzmSgiUzVYtid7EDxM+ed/y6P8AV6aCsdKaXa3HCD6lp3OtNfGdE+LRR2rkXqdqG10sDug+u
M0sn3j2XTehrT7rWjc3+vuFBDbgWfZz/paXaVbuq9li0ZKyS8UxMNtYANt/4OnbvOCPETtu1Ly9I
2mcB8718Jdi9j49HxdCfbKDD6OfFksugX5S3c54GsySS5oYD8S3TozcTheIdlaos6IUlRAj3MWy8
q5h6LtC3nIXUAGUQfHg8/s6pmfNCTGaC5CRTPq4U0baraq8CfjcNX+0t5SKR8DDEGoO7UktPbdli
zk+D2ZnfbSQVa0AJFg6CQnkBiYz6ZM8tQvsqdyck9CwHrAF4JVVysQIXNhdGtzlHwU/QgLd6evsn
SbId7WDq90Hy88rlEIv8G+xl+wx/PwvJHjGQyKL0PmyT6ERegsB5rFOl4JomZsk9K/X8aIdtxvHv
VuLGF9YXhMixcpqat1TYR3zGyQXIWd9OjXxClNMqJogOgCKf8UwSPTLw8d4IZ85rpwVzWeqg3x+J
lp1G0tAj+kDw5V7cvZj7awqr1GXAJ5v+kgNGgdrXof5auxkRxORWr9esoSUb6gaWYv4TRjmOBZ3f
W+CBiBtk4EOKHwEhleCWevkgJ3RFhTb080Z7B7OC/Wb5hnVrUesGx+CGjKHcMYnpjFKll1jwjfkc
rAFCeDhvoW04orR+cjNnU7R7IuF3WL/N/6BVT0wIuaG50Lc9glHgVEkgP2npdEXZjqFnjJo2QKfm
EBMVx32LZs+WFTgD5x/0LzMiu1ll4NxzNGnEBOZzgfujUvtCGNKpCtuNkex42GuU0TkLUxRvkiFL
QAo3pEh/PD1CM7lzlUIiGrCaB+vC/tbPn2w/EA3+w7OGNiWzOLcV7Wn5IFQuCUR67UWQSe+ZzUlQ
k4tw5dlywNMs9YqtbS4xWLZta25//urYy0V99iCAnnKWBekrPY9f5KjcBv1/u63ilFH60oHXeHY+
4I0DLz/hDGXn2Vci8KvEtBRVcReAjEQeMBH3l7XirNBb/65a3zjaUU63kqZ+Bd65JmnZbh5tahyt
/tKZQ82rqCBOxup1rGRWHL+XVsbMLDNL0JZvej36/WNbbxj8L/99eZTwmGCEDqFZWlZJnEWiCEct
9wag5UtniTdXx/2XGXXlV7vbZNt+/6ud2bJd9DoLT6j6GLL4mw3+gjTgdWopxu9d24GPVL9zhvaR
4J6A4Zjvgn5sPOlFWz/Eib2ePhGvE1AWHsX6eNCpaFCNG9/rGQwYU8g0V9S2MVF0I/JlTlXGkaEq
RMcu86P+qfQYRjvWCA8xkK7vQA/UKwmfSsvt9g4c9orXiQjadVMXGfe0YKRDQSG+sxCOtyDXfBy4
AOIQsMVM/qHY1WlAbRMiy9rIZJQ+MVL0sCz1tteR8X21kZoFyqQBqc3NG3Rz5HqgGC8zAzepgtZF
rvqZH0RlEl/ko9oMYkLzBcftCfp2KWVJdXVKzGu6jJburTdhEywqrKdg0rpvdYIf/WK24BX5/bim
UkH/5Ki5THydY0WDdhTjNryAOYvvgVJM7iwIAwmD/UmLBZd60fQUAPemQgY0qEDn14udkfJhnmOL
7q+Ik2cR5RbdGJ07Zr7GJpfpYPQMvWzVLVbNcgQcud0QxQIlpk9xIGURapV+Uq7Eu4Xj9vlJSSL6
x9vjZ7aHeiNbzp70/pbJjGZv7tdL5ipsSfUE16rqA4OvkEF9RZs/cEv8k3EQXVzEjqF37CGgHbx4
+n7YtpFTtD5fJJCzIknofk2+A8HcsqK8YJ1Ph4EqdgKGVqUcfU1kFCS4jd2bf0bW/0ZELDAz9/Ck
4FJQd72OZAT1+1lQCs6+9OT8CrsqrcV9LKjfmbNeWDULCPFOCGpHWQ8I3DMEDKO8SNNiGGkU2y2I
9G7bXYeigwNucOPDN6mgJYdNwZYW32kdOWipnaia8qR7kgFwIdIt1h3reWVgW3/zN7ck8std1mY5
P81GGDan9RY6Aq4CrRpmvboM8rbGa/Z80LOuRqxGk9ppM7kEMgdtDZ3VscnCgqTd4oqD4syiY7sF
1Z1Q2UnLofmCbXQ5y8CsUk7Ad4n6RZ1Xx2U14RLj2kVAQIys2cL1ZO4UfXxv4ibUNKrImL0++Lsk
eypwsC2df2lQHuOqPxtI3tKUdOOkDRYgKNpDk1ILL+I1Yyv8JqsydpRk+LsStelP2DOZ8l0+TDqm
qVVexC23UY/qN/yhg1aAUKT8gaZhmNgII04T3MzkgFIpru5JePYygaEwhV1ewHd37hsoFugjTKeJ
AuiAOxUcR3PWMz3sCSoeWYBMBwuYQKGb14oC4WedhLb964EjRCZVZ8qfqNIFkztSqI6V0wATWNNj
+JfbTIfUkfBj2Jv+uA8cmcJ2cOHNW3IoVjqZsh2XbLzA2g0/mLTQeJc1wO+qWpeqjipliHnTqYij
Fm+DfkaDJgoTUg3r0o4tUTozRPhmzehDw/HrZBAsH8p1Kr1jg7DGJYtNGmaTJFQsdGzG6D4kSxX9
Cfg2ofBMIQ4T9RrtEao9+Tcp8slG3O5fRtomrW1T7ZR5tO9LRZDjZedhJJ+DP1Q942+IGt/suN5S
7vWnTZ8smXtKtYvet0dNhYlaHqa2RH3DvBY2lQS6e7kclxX4qzrxna9/xuKJX8pTCph9Cf4Y3dUQ
yJe35+2ZCclRU3BZI0B1nTqSPGVyvgVKyHsTXu4gqm/h1Ss5cGE9F+SXncp6EDCdeIq9IFaxrllF
IUygtRz5KZj3+GzMbX/EYve6Ieyb9vjWw1FMtuqGlRu6tevp/LKQ0klDxSsCMxXkMOgKpKEFgMp2
wXQhKG3vuUCbesLfSsYTFiOvSmZw49Bn6dAC3q0hpQS0px8nzrLBqOZfyfXqSHpx0K0FAOUhPNg9
idH5Vf/Eb0qU5EuhkYm0JHcopb+Yy24TqVcIt/6qrOSaiGI3laVcIryClRTrRJ1T2O8iYKHOereR
g0uKG+dLUE+yxdvK4QcSfuMx2qJSLjLbKtOxQuCzWNe8vyTP7o0gVvZ0a2r4CBzEsSjGRTdM8j0H
5ZuDgssh7ff6tmnozJFZ8ikHZjQ3aXyuRN678EiRavc+uRCv2H+ED7OaTBYlznftDBgKPoziaa69
1/i/W0kzsLtsPnhW9Vo2p+3GNCbAbbEtppVhx+b7bn0NpTsTylbr+ChZr65j+ClNj7OUyxOYpCso
Dyb6aFhfcxog3nluWgUuC5JE53f/NIAdIgbmL6TNfCDXkdjxpDGkfP+Qy929/HykJ73D+J1YUSNl
6yTvaT5/P8HIwgSsxkXthk1qsTu7qj4/5k7kJs3MUpDyr9iZ14H7mTOB5sToEkVhQI8MOtTct8Wb
PodXwyGyg5qnxCF8rRHMc9bkHbmY1O525JDh9gERrCcMkb5EYC6eUH7xBm9+MHpgYPKEl8iPomAF
3azO25dUFAhci8+5NS7vMuJqUXvfIz+LLAZgfugPERA1riewMy+gxLb9Yz2RPN7CfwTnUldU0SR+
2UWCQVJBEfCXkAp1PQycMo2VB+//zEORVG2wJHEGgr+7Y4UJAwVAPn1XcPNKkq/vMngYyYq+ep5x
QfuFc3VwiQ539wD0qDIoLH0Ca+bA1Wf5S2HQysVpzAU1VORRT4t8r72Wgi652pb/kPMLVvoE0P4p
dsuWiVkKRSJWdtOVPMTrk3bTYfigFxWN2GU40pvfBEQTZXEltf9JhcksmguYcJw+FFDSlVhqrFqC
3/oz1uEyku67QdQMCgAYrSFRm1H930TAOGNoV2r6k52q/VSXUOgiQT2sDVDUbRJqCWWw7xjXM6wN
pxpL0wjdEejN7iGAU+7xYS/BxIs7449mW11pYhPkDYcUszcj1QeMbFyZqUthjoxiY3aSvcc6xXG1
s/qVTYpzrzGDx+QsY8+RcAnZcCycFffbFrKdCIwjwgqm6+Wbwypvl5NxuaP8xqjYdY+YwQe+8684
7iuNNUZvhrslNnEwrZkIKRjduVmPtPE/D2y2xUbl2NefecI+/jqAzMtuN6+VVYNdXlkZ/ahF+TDp
TOXLDH+msjSqWLwrZIv6yF4QgU70MZktSOi1C4iwG+NZiYXYIqZIu3SZ3Njnn/85ULmuc9+vusG3
hcbgsX7tBsioH2tGPneaFLsa3LCDGU4U1EJjPZ3SDnrsLS4KZ7mFOl8dNxFqE95NNxzFBm0Ij83z
o+fcMeVw7qdNbxhfMhOB3VMeRdQhE+6JXiKpSvejlqGavcGXBmdxdgs/mZaEFh/YEyvUyrJ6FSpQ
VjRuKFewfu87pPnXHc7T53OdEPdfTmokMzLrsOARpAlZ2LxIGS5sFA1pDmjii2flOkwtQPuXny8r
1uyY/vdWy26Y0TeJGRgm2jdwHzDcpbj/j0NgJbmUCc0IwG1FHuTXIfX52Io8ogj+41Mqjh4yr44z
5wQQ64fawlnnCcWmYVPzOxgdsX/7ueE0FfxJKzJF+LBaCZlaOuaOFpNTLrJicBrvlzMHfOKHMil3
4oqkcdpDIg5rFb3zt/Yqkjki/1zjkX750XrXufLWsblqAw+lexAxJVoQKTlMMUAW0OLJPuPxe4kv
PgHLWCltUGqquUirQ9wfbjFzwgUiRHT3IMiNZPW6HWeUuDtp4z9KckiSpqIWAawQRWP9i7qz89KO
BeT/I4R4SOFRUZHVoj8FLFPj58hqLm8dpbjYcp4qbMUA2tiIaVs/iBdxLfeukWglrhCbGSUmffgW
JvQFnOgM06RwPpqNFSSDlvRZ69snbdRJAMxtw4FrroMpRJHlFL1ls6Mp6GOa49hRPQJnoiiReZK2
rB03cc2Wufxbqoj1KsglSpi2Ee/E7dHiRTf5m7/1grpskk5XbduS1eXznJc4g3yRxHpCbsGhY8I4
1nWb2dZNbV26mKrmL/OyJn1Bj2ZLfgkZOM81Xgz8bn1Tr/jKmoLMQiEb6G/5PeKTvFaA/zEy9fjb
V0/EwL0Duea5UB+6oEQuswhUPY59y0pv31/c0wuRWpde2Vc1TTGoSbf6cMK6KIAt8EmrNgKRcFZ8
7ofJ1IRw7y3b4K9dxnYIlYsJJJu7MIgKEeYNfWfjY+tbvsp6c80EAR5SzxZZKxq8rMyyZK/ZrkRw
aPydcYd+Jd5eede86uXRmctik+dqOYdyyR9x+HTbBy7wgEOeq8gZxWmZr9vH22hG3UPUAcJFBPAL
C+in5EKHz8sj1Bzjdi9g0auPXLfIORfwoEo1JnMUeALqvpSZGwRMe4vr32C5sa8nkGj12cc2Xm5y
3TiDXLC57bf5ebx3/lBEIdreEbax5ojpc54kJGRFV4+8uDYJsQnpZo9MFaPsBBr+4T8ac+Hv1jVX
phoWzlz/qY2UruEPcPQE9WJFtOwWM4OudyH2YW9SgJE1g6q7w3zT85O2GryMmRudy6vQ7ayuSbcs
adUn5CNkCXcDoRFCihyHI8uTFcxoICavAifrNVuEjAFlGfHkZxsO6gdk7O4pT0kPV0w72axK0rn4
wiYR2T8xVctiTDrrueJnZJULqyeoIwTGRzCG6+M6PC+voCGl7OUCT++5NMy65F4E12XA1gOICLPq
wmvUilNbPjGpe2CHTd/4+B8tN1jU0OKsqQqQL6pMkt8fW3kXDsU5/dGQwMbTdonDzbvacmQIJpRL
1vWhGX/MC8nPWPMr1uatD3DT7BtpU2V5S+RSIDtocBVBakCW/edXPuN6LPqMlsUtmwcAuK92+SWC
x3Y4LmeDU50GEbwYtSuyxOuQwlG8qRQCgWlWbQFLN2l0WfRkxSlh78BhAhCMotNeDZ+JSM7IALRU
r9YBXseO3VLjg2ZtEGSRs0HkjXb1rWIxUpHtnjLwCWNpkMpNqiVQHy4635+N3YJNg4wVsnQ06bPi
iul80RhceH5CAGryk8VC73yaYctOM+Fj/6KxTbE3jznb4VCea2cUgQ7UaI69Tlf64yp+3kXjxWFa
BMSn4Us4xDSf7rnoORRK+DWuMeJHuiFa9chF25IDwMGg2HkpeTv/bg3Vh9JNaFUUecjTKRULBxmW
SoSch5KC+JSbnrOsV6kLgOiC0cNOH5pNO5dahcmqwru9fUKX0GeNdPh6nDF8E689v/4wVyoxypl1
3rODvOcU45tWZ464gJEFBJt2QnZ2D0qR1h63g5/3e86eUqZ+PXmnzkIdzAKz8FnBnpst7IHYqSVl
BMLKsk6vCNeZoC2CzgSwbJaU7XjH1Ffvx1qb0Q5B75gZaVQK8aN2D/H2q6g2I5PKdtkz+8EDDhai
5wuzzwGi/OR6l48fQZLqcIC7um2PUlFRoGkTUkZUfT3osog6BfPXvTeQZmwcI6JXrMKFqEHSRN3R
+k65vPq7zEyKvdOPT2N5OluiBB+yj7TMfZQX+GgwUVc92Q3/SpslKtkSzQDexsbiCA4CsAPAz8FE
GzgKpvKbZJ5JePNZJ4pEdcn/2okJbY/O/i9EfxTASgpqU3OQliydlCifC6alfYFvchSxacFF12/s
pWebSJmdp9jhiR6oZTrDX5b+dmmQSMQ2UViH04aLbseMOzCnYlXf5yFhKS4ulOvWTcLtRwt1+iz+
d/WsFWE92Z4T9PqrcaMOaCrbKpxa64K8jt+QfyiRVQIFAnPHp/h44knebSue84a6VWj2UmiS2Bmg
f4OdT52C2VKDtaufq5be2El6C8yt6sSepJewjWLWruIyZuVvIN0IUoDHjhj+1K9f2drV4k1OiAyS
ADUkZgIbgCgopTeIzD9iogYKiwr4zyfHsQOvg7JEWcU9jQPImKNFoh19nsr3weHHMmVA2Vj1G3Lx
5yZ4/fY0LBdAQ1q3jebEVjwQaiQZF6hl//WV2birSnpz+HW/Td6SnIprByCtr98z+6mv1TuNAyQx
RiY9/RmICbUJ5quA2YiZySuOhr80TcJml736RVrdrN1IrGux8kEigvE5JbwKplFAZJtC7QIVEGSu
aMTIjSxJlEiN/2HKm2DxUdc+NuFwQ4uirRtRQUU+y4msrmQC9zYscX+PNomkbNCMkU7eEOT1fQ7l
CiTq4ggJGkV1CholVuNMUTF444Oqb4MYm9UxgF8ZxxmHX6RS5Dds7KZYOXxu49UeurxwwCU7icSy
qN3A2LQ117nYYVTWs03ZS9AuS2/AFUggWQPtRFwvkPCfMoRtngQJsDc32/EvjtD/fsLfNcNDygZV
3N9SU/ke0di4anUeBquZdL1FtU8La/yhnC7MxlRKIkQFZt6wqsjbfsbcCHaoDmgoM42SncSypwN9
M8XxkNb1vfZfbukrseXx/rWLpkOvxxgEfyE34OL5U7wRQslJTApMTxmwJPhxnn20EVaxbhGdV0F1
6IDMSZC3bUDE9u2WVpg8WM1gcqRXbeYTU28q+PPDyGqH5m8mROdnYLbOuoterxKDrIsThfmfWTeJ
5XcqabE94UeMcpV9CLPzhqL6otChBpNx9w/HWs2nZArG3v52OL3qGq8NynEPhIp8R6jUEMS+9tHk
oz5CKlqZhaOpHde0heCaZukENrCjCKxO3ok+Y2tG05wY1rasuKn8DRyZlxehDdFJ2dGFM/LoW81G
NUbb+uWYwH63zvVLV30xHFYwuOqfAcIydLisHEagNv3vpiJXDJ7BZdEpGyDg2A3Pg0EXzA9brgFN
ppMbGFVtv7/0xdlQANHUmfx3xIsPU1C4QHqWTuOfwKnJ8T6QeUeqZCR0ckoWRvqzppjxgynGgCz5
2IYOddQ6CcuFu8ljDGx2PmdQQBZdOT+Gumft34xhlf4fLF21kyq0k/+oW4vvMBQIKljedI+k/2+B
I0kfbr6e3DtRrGYbiJZaciWjV8z/OLILWr131Py2u27lfNXH2rY8qH/5aYBRSuSckGPoem+EXNiS
9EORO+Igremz01H7FsCg4nD4JzQm00th56t0ZhFoNVWqQ8AyOYp6aEDGYcQpayUWu5ImzuGG6aJj
LG5A7oGnbxQgdIKa7mIsxwcB3w8EQ4qK/seIqYSvra6UEjJH34CXRWvmtRB7Hj/8TXooyPxYOhKX
cguxWPU2q3sjJ3xeAS76nC3dJPwyBhdzmSBmPF8rKzeH5yaD+PaPz1jPgwov0wwuN52zms4qnKEi
+uDZ2j6ybyfyeHQCgpeERp6A6BY9MKIPJ8P0JpOAhxnWmHtg3xI9yTt4aSGXbRIoImvtp4etFvMR
TrW/TaTNnl3HB81v3d1A7moW78yzxbtLpIMwhDFgxoCCruPStQ2sb9mMkgd6pjNQPfK3srQaBcD7
Ir4weoD0XrBm4sw20XTkF3AWQCsPaHGQxfM5pcq/KseWixnlSVTDhC8hST0oefsAeeXewrxJ/eif
jaupXA4pp+VOILc40UwrFcCdKmXJEAcQNVKz/3QEOmcmDNNMN/FSwQmiAxN+og36Xa5U7PoXhejx
eQsxUrsoqXWeD1c1IzWqQSGDtcjEoRnt3h96XjelNPNvEWNjIydKXaZb3JEgUQcBuWVE29VrvrCK
cTfyJFM586yoPQHkwhRkUyCxK2Q77pPauU7gKCI3v/N2KoPjs+pFvhyVajvU8+cDOj5xAJaB5P9b
aOQ6rG6TlftPKG7QD6LNGrCBwHXH99wrUsYj6VVo2SKIxK+8wrgnEkZK4w/HYoXDnfuPTQGAKT+6
/4VY0jiUu1XhDmvon5M8aI798ZjdXhOB0GB8CxjJsguInbBVKHb4AIKWNF6igQaNsqt0r2TrJj7l
+J61bUU+ocRKXq5amfyJ4k6Y7hNrYgFEgW0Odr28eJL4fLJnYpKnnDon3z9IjRFy0d89SXkMfXqi
OAZzMslXOK9/e38pOyu/jFIpyQe99NCq2RWGeOvLCZVYlg6Y+FpqEpcWd05Xv9OwzKpmU2Gmcmtd
VuEz8lq2WwAiVh6kldgtYPjw2rLagrRjg5kl1cH+A4uMm2yllruO2IBN0Kwfl+7itQeqwqwk5iG1
JnrwGGuY9yVN0/FkGXyUnUjYXkfR8lbcMAWgVi3MVpq9QV/LN9a6SgKq4fcUalTvgZRGeHYw0C6A
MYhCKLam8Du7yWenaJVECGjU3DLQwVOyYapE+S17lGJ6WA9ixYmVAAN6wx8b9USulaJ6/x6B9cP7
CtHDIFwfXdb+8eybPdSlHFOUzalVa/cgNELylZuyREJ9bjxkXzv3CtsNc0TK8iTh0i4Ftlk64yHJ
8nRxCghXH/71pN+vRZgjtesDd7PFy18qZSWrttBB0lmTlwfU0WtkV/P/+mAm1+GP/Ap3RQyjksgV
FlA8M5NXuj3dKD5QozZUqhIEcIu/CV8SvtY1PNCSD/904QdrsUUnowPgKB19M3gofSlLX7d1UTXr
byRu8zfUOewrKfXt970FNZ7yJ/BspxC7vs8vGlb4XIzMCSSlFPvQ5/uwwS/qHlvPxlB3SRK3Mp3x
46V9gOuzjequvipHVZbbGM3vXoYdl8r1n2Hma0Kr0Vqm6NKKznJl1q+cgBhZ8V7d/+Ktc4FIt73A
4LdiIYZwjP06aQcKvX747w43fz2KRirFW0xDpPuXKFk3lZtoybGDM74bwEjWZs1l6sbctNdULtc9
pyP5Ss1AWxesslnQs+4EwpiJA1y70JMP/IQwIOG8z638J56CewVec8/cQHRGuLpv6gjkWCYr/3TY
L3YfciCnFVRuehdjS2DpeAfMA580mgJHJJluASpQQhbk43W1+bPPRoyc2ARECrjtSA7s7ZhzeXfX
XC7Hp2dPCUl+FrGVknLj75ceNenfEMFus2GlQgXB64+tCYyxdO4jrQzkMpRa9fsdHzBpOEydmHfF
mWDbd0qrxHMo8Fx0ZFSk3OUgekVRuqawfpmWazf/kragUPADKIeDr+9yKVF0w0mxMBHL3aNQKXC8
WRYLRQK3PQYLF8ZHx4kwePFlkUA48NpnRH+AnKAnW7wvqwlwP5lv8raDsb8QY5PMdXTP0WKuK7Qw
el8GCpuoACZeAcG+vFleXfbnQw2z+uK6jXNyC4bZWRaWxWduxcYwMnGkdW2iXzwgXtjs31M3xRej
YjgvF9/zAuyWQc4qIryMDUW4HzGLOWSaExlU7vnPabALxKStgL5q9ySdkS2Uno6JZXOAxvOY7wwU
OmbCOxMdEKcS/joGjOBj049L+gN78zDVji3NTsnrfqN4PubMQDfZvpRyCTpfMAa96gXPA3pBxGxk
f9QebUI94HEnHtN16B+/fUtmwoJgHcJ037D9NTfIpLCYy7Ii+5fnY9lFukMqm9YQSQX4YhZ/5kmw
UqC07xUInuMlm+GQGeIwaI9hGLqZGJtYvWz/mtHHkszPBsPsckkSd2xuEjbWqMH/Fs0mHScO5L+u
x1eEcbRKcAfPQgTJF38sODq/fmOGl5qVSS/lKtnpp6czMmsbw757MhnucBqkOnV8mrz5CNLzgT3C
CqHh6P34TeJ1z9YrDnS5cphnlKXsHgpDZxaSubJX78samBFsU3RkxjBR6w+h/5R6Ld6iYcNONuen
F+g5shrAYiMi1BAmvI39d3Ayd0dPDOHrLzsps2+Ma1MXhaHtlMAafwrWzx8l8vWOUXzhl8UUpst+
FTnUvFIZiooZOyHcPLpt1YgFnxe4VcaCH5LBxJLZZ8rXwKlnHiUEd6Ssb3vyxObGo5qzd1l+KyVo
0belz0bPvJ5HsQ5fqd+9lJCiTX048XkMsD4l5dTgDHedwDmLb76KcoGskjzxyG6lRJWPXyAYIRiC
WkaG0mN5r3H5blqwzQkQ1f+8+pT60fBD89UmzezUNuuwWeQl/7ulvGI7hIByBt3+iub3eCKszyKs
guOHwceAvs0QIZWldFV+3DDSyUnKTpvK7kCnC8Z6V5fAFIFal0c92PATFhNsyyugJ3Bj4sFlHRL9
K0bI1RJbexr2nb6ZdGKA2+bZ3WC9NulWiIsSUN9VjBWcLJuSjanZ4nDz5xxHrMdODpj/oD276HmF
qkyISJE5D8QzErltW31qgR0vIrFT2EpU0v5vyECRR9xsEmuVPfiitwfeyXxh1Ps0nCV8+qRfnH/i
JfybWmQ9Xz2lv8wcRH7hZWsTDyXg9QmtQH6nAatJGCwBFIkn3PFrABYMp+AEP8dsNU3fGTNFxHou
NYmwIGyes2azHZN6ppcEKYhQSDay9RJ6LWbs1bcarcAxnOeCjQ5XiXcSErIEqMetwk1vakQ5WC6R
qrcSkyi5BpHgD9TKHy2ELaIvj7DSHH/1J2QqhcHZW2poSC9JSgZ88WyU6+kF9L1EjhuxL0AHBlTX
n227xWfyvVymFzN6lpv9LlmoVnU1HzTBEtBYyryMo/vSUUSxOQNH3D5OsxxmyWLMX2yyM6oS9C+M
Cg6hkpme1IojLdodIQMfY89ypzg41qacZgGpiVt9WjlFAfUxGaUd+C1cP/wIWs0BVHlYvRLV4fHo
BjpxsfyfKpyQprwjvrYCvpQeD3BIuU5Zld3UcZjX9LpGNScslwYLZpS7OYEkJUbuigbq/Qvjyk3G
GKsQuDWIULRnQc2IhRkr70DpgJWmREL46tZE206M/fHiFJjclxRx1/nhg4CeNWZQf6yeeoV0aaFX
1KX0cDRBfjtEMcP2S+C7N3PtVLcEYAxFeiFSQe0Cpea/SVtTo3P57PqXfN8ri3yVo/9nX0a7M5mX
UdB0FY4edkUny5q+WeClVDFv/46LqTtyk4Vkf4Pr1DfJW+g+kNjeLCgFN6Lg6aMLTrsl/6EKkqB4
VgLDX9ZZ+RCNIMLwuwoh4TJFQURnA0LmvgOwp06vBc+N9kKz9FWZ4iMJ2j3RRpk2/A/E6zNqmxFt
thjVIUsqHswP5dad2jBkntzoLKQz9DLIT11KisV0dYxTRTUkvhqgFbVvt6HjYty0emE+cGjpdqQl
7GByya/h7+gFqLHirlj2LTLRoVB6MOF/h/poRVrrddVRYScw6r3oSvrFOmKt0UZnYVl0gwGTV1rB
cvQla39RsyYWkbpKhqngKrPL89TY6PxpZ7IJIACOW7rbpssYTCRhP09gQ5GmMqtWMXfj71kQurSG
FPCzg/drTdukUT5TpCtzeuHBs+UvHomMhe34dX4EC8ZUuhLOa9H80QuZHrrfHTm+0UxSe14ElmMF
JNqi1PEnrf6WKh9DoA9XQdZB2N9gwoRQNFt0ykmA3e0sA0Hibn0lWXDPQRfFTzsByNJJqlbqIPph
PPRyAnsz8tqo1kmInbhIfuDyQmagjc5KPT5x+DcvU1VyTMPLW8qDRNIOJymBgMaiIHtP//R7I+NB
LYT2Chv2r71uLNS/aqqBVr9U1T3JA997txzG1VxNFsua71Uv5m5+EXQM7DqtdVGT86iIeqFxaWPz
7JBbHso2+82WTiwfupHN/ZOWQnI2OFza1PUffpDCx1hKNj+bNjpvlmxX+w2X2VEZ0cyd7/OUEuKf
Sfl1+sZ8pXXoc3V/yPpuhqMCwE/9oZNzL9aiBTRCeerimX1Dr75LaYn7lsOpVW9gRtPmv2x6au3G
ArgpKsGvVbd7ok//Tufrag7EwY28EWemcdNopdPwarRIFVwVWpsma9AyZaq7Oi2cZfA6suoiyjks
MovyQG+RSX5HMiQ6FUA82WUIzbS6EBZ+XF8hE76rLSHhlQQxEeFlaMs/C1XRr3n04bFHUR8IAdkj
kmoU1O/Yqe+yrX4WWrT7LCp8h/U51c/tlKqA+2P5U1rtq1rCuGcBEZlj9Rvln6aPxXLnA3Ey+SQx
y86YDBIfIwi1kbcvnYRkmvDlbPjQVUlqxsRniAomLOLBp/O0wBo6kWjvdea4CnymMgFory7NNk46
wkPpQhwrTrrh/5YzHPfKYpJ9P+qcSsUcdKNfNlO4FDkIZ7E19yA8MWkq54J/9kdGS23MhgFqANKP
H+iBx2na1CIOfJ0+4eXNhS4WmDGpOZjUoj2jVdp1QEvOXowZkV6NqhrdXcNad1oztQ3/1kA18PD7
JcPONJq4v7AMtse8CNcCFZ8ttGsJLjcLT/qg2rqeiQ1OsIbONPKLagMjaL++if8wbaw43ziozO+d
VqZffONwvZPwNEhi68/8EeiVju5ap3zHMxOkEqNCmxPIQs7I8GeVjXcX8EWtqCJF9O/0SXX0PPCL
YWEl0Xs9mN0+HfwkBh4lUWxNFOTbZVtU1NfpgbhwIwqbZh2N0dau38wpTt7EXz9etp6VuCMyEeF9
s77yheSt/RuV4BFfv8inQ8aMKpWnWPyt/igX/vuaQn0hBwFw8d64LfcNkgwhnYtA+oDVgucnNZoq
28b2uLK0iyZHNXX7qgoDEQW4Y4pkr/vg/d3NA/xTQgnJu7sL/sn8Q/x0lVkSAxckasTh3X+8zm/P
i76kiiwRDjF+2dPy8dF+SUmzJAlHk7mvSwebLonR9AAvoxbsxo9mgMCyLvNebQGfu5Lacd275pjP
VSobcSlIxr10xzzP9tKEfy93dvg1Z44ldl4EpDn8fiIbaBRikf9f8lSZd23lFhNyeg0rlAunLYu8
X3G/TWZUTHntFg7T6wOgLP9IFwXTAClW5kPxc8N0NHWQjLI4XFQVVq1I9Z/J7g4eHwa5+fjXdsAM
OnwvT360jVgD870BRt8rbqndbs1+EcouBB3Uxeb4GZhxNDe/l1mci0CJpMkrfbjYDVYsiFWHl9DM
ApkrZMc8GL/BeISdjxBadN5jeoBzUgBuEMjnMvBGKq63DX1pLe5iGjxCZrzqw7zrcQjnkXR2qRGc
5xZgzcUJQL7DVQoGdFhOgHe4yoy1tRMMaTqmGmV9w6mJ1PJ412rCvwbar8oVuC4+MFR/lAoSup8h
QODiFSi1qjOZ9a9DV6g9RaWyBGOCZpg2VISey5dm2DBZfRSY0CYyGJsKxuAhdd1WeOmP2RItgQC/
fsiyyBkA7zAFEDA5FGJV9zTG8cu5ay2J7hRWqaBR7xt4DsZisCBtcxRJngN58O6r3pyb3dIwIc+5
MDD3EkxiFnvoqsbuTzFSzV325IJNeq/dVoUlCC2s9939jPUOldy/cXI2B4eSUjAUcQGr2T9Hsv+l
CSIZSLiRDCYJSopgLzeEpw0JhmtzFn/FakbLGscLyQz0G10rV7lkKEgxslfY5onYjZCC/q7gBypo
QRag6UjJy2oSqnXd/OyOpy5HfcQM6PHwOpLJ0EUEF5YFCayXeP+PDo61b8SxeZOnmvQZYoR82A5F
QC6Ug4U8h3Dlx522z3Oel3JtADBj4IyCF7lrMlA4s1OhWefoEx7CMAT/N663c4SGG4a5ZAN4Kd/n
fYfd+pIYhBKvJKwFal//6g9l/VmbUMIi3ylfBpe65OIADAEVuUL0ofI8/NvOS+vWVaaNRSD8anYm
xLRvkz75lFDfHU6kGp5rm2rMMwC2QEiKTBQXctP+cuBWJztTzvPCJUD9d8zyweNbvpQSL22/7u0k
ac/3wj59jlkgwzHJnwWY41Nk4mrvs8sTDXTeOzn9sD0nWE0sTkXmzuxpPI3/e4bmuP6Kw2oxTjLK
ukPuupo2210SY1gwMrJ0M74ue1dpNc1MFonjmzdnxge87ydP63vM/lI3WeJTA/JlL80Hx7sDV9Tz
st512npErIxMmQ8eCk6/22yMV2nySeZUizAdFM5a8nMvAFt5UxIdpLL6TzxuNmDTc7BItKadGLNi
mXh5m26QvTRPTlYd732JJ7wEBa1E6aBwhdycHPYRD58Sr5cNb81SMcMPZTZqbDiyVwshHZmqBHUS
Gw30SENjP7EXx47Ko2ET2R4nLDQHD7MByviChBcXckh8fuuqiFWP64I4RsNiQk29Cizk55U5cfSo
eniFRPdyOKfeT9e9fLY1b7S8I8QJrdQHhNNnYDbpm3ZECS/Xmv+F10He6z3HDJN3u89BsRSM8+l6
RnLdIEYnLKNXteN2m97C0igqhGBYrtirxzuy9B4m1/Gtl76IFcWIVCF2NrMdijhwqEuo6k7snWbx
WvSUO9X6+WaKtKOjV9g6+gLGhBsSGVwcjfyWRTGajeBn4wbGNsfNNUyn3Nlj7gSG1tSU60iBezJ2
73pKCNsf/oPTax4tAVS73AzYybvnSPGiLxuEsxTsvJRIOFiE711h56SPfmKiZsxwZeQiV3b2s75y
pdXc+YqXqtm6mNBrKaOTJqkcCuPuqy0CBRKrZuEU2MD071kC5C1z0y0/OvuKBsxC5pmiZtnF00ug
a/oHKjzJ47veK87hlKoFv98xoS8Om6Zyi9HKeYkOchNiGLhd4Oz8v2aDx/KIpUf4DT+DwN5VNrSo
gmDoOyXJ+lx9bvTnBEmykz3gSbzVEOcT5QbKQPMB/jEebH7Op3dwQ8ur5n6y9m+PyZbhBrwBjFb6
UOdnaErjno+haUgtWmIZ9Ui8/fpdFENnuv95Re+lx/chrsm6+RnlcUUtjGlylPU/LN/HPReMVt9+
ffPpcjs//u+g69G8VuJNWWJ0DXapXnz8RnAfsk1ZZcjxV2D9KCNgz3OS8cVpAO2d4y63o1OeMMfo
a4/E8FF4bIqUqfA3gFqJNLJbOu/qDzKNGSyuZc63nD0gG1/y1ZOh2HdMu2EmBwM3tlURj0U4CFqO
tMxgPGYGxYt4bAjFiEw0D48X6RBXjL5khabeZmVmglDAf6wg/VK+L4k2wG17HXVgBRw5nGeVBw07
DyeQqXATAPUU08R7YR/rFxAtld1cYgWEtBA0piwXSzP6jobHQ6ehZCAKf4LqiR+gkh9yV3Z3NOx8
VZTr9xNDHva8cA8zemSOsCY7lEqlE1dgCofjrz3E78ADWdO96UOwoEBPuqhPhphqAjWwKkCgfTcx
GiH+MZEjOiyqIc74xOoPSHQ1D6jkD2F3QAY1r9e15Kfjiz8yblIGBlfc7R1MYJ1hjCfYUptsqVJX
Y8YjjBvbJtANl3hXMtSyPyLMDvlahxj+aZfo29FqQq5azC3lxDM9AOvCb0Zjda1RQ0L0MmMsrgm+
bTJMBkmQCQkGbFPB0AEij2xZJNGGKrkxCurlKa3LLs9zNYmUlaTXVWq9BAnjeGYDlmNa/+L+/jFx
Uyv74k3GvyYwiCWrrmj8MeF5f3JlT4NtO6iJSD/fR+8V3LM2FyWmpaVmWTxZ3y/ZkgpQvAwc0fS7
R6ad36rPbAIjMyCUo7dnqHAxW8u9NgGkS/ODuRtE53MJ9ZNCFpJIUl8edIsDKrsmGJNycVZLfHp3
+VSk1uvTOvM/yapqjF5b9sfPTDC+eJvZ47k6Y5pNDqHIKdpjnoQ7uCRIrKB6rLjSN6DStKP9mf5v
zwbzcuL+ga83Dm/rjpILrOB+jT3/GCEQv11n1gZjsi0CbbiaOXWbDKq1lHUrcN9/V2SG29GdSejo
Gwo8m2nMxnCDGyT9fYp61mxVKnaylthqFdCyzIlbgNqz9xKULicv+ya7m2HcP/yA4KvRYcUyMmAd
NQxaK4sUTBByOZFd1w0G8XxFxPFg3g+IrzZ0pwR++Y9qp8fSuOvbxmPrhJ5Wx//fn0ZPGHaI/YsG
cqUKsF57I85gg3Q9IdHwbmRcPJ9Rwot6eS7p0K0tiE58fcVGAgk3touomkcJtMtvLmdIhIcc4dWt
m8EqEFNLe85wzVq5AMldQYK+BiAQnHhKNqFDZY7JokYWTVblaNxD1CFMYMuyOIc7jcrGMobSYh0/
RdoF5m62reWq9Nail9LJwE8jckSeoOpRXDPqLTzFNej4FXtDeGCHp4q9StqMXItVwAV4QUMl7RvY
tM1UqydJaRIkhIOPe0CMR5wdpa3M2QKGJXkzUFPPxHfVqXjaMOql4MfuTDL2ym98+MwN7p+IaEdv
bXxLqshyy1S8sp1o2d6bp89+DCimu+bPL4LsKNZd7uG6wVpSpH8yRMAeOmf572cjtoj+LMpZo7BY
wPH3if5n+g8XrrjmgVYGGt09UfRQt+KRNhhmQX8LTkAMjsyZLTMrUXaqGgQarmxi2/6bkHHQwLA+
Inz+DCn0kRkk76fMwRaxKol1Jf4PozfscR1FCg9dSPNu0YvKZHZsZheME8VFJQSNB0OMdImEne1M
2jdTNdW9f6X59wRIRVdQx8XEXSa4mcKHAQ4ZlhZzvf4Sz7gdT3y/JV/nvNqOdcYs6nY192LvwheP
nmiSSAe11v3AboKrnPMTlol25/lmFCKgupj4ymxqz6mwcNH6a5jhI18blgk63LOHoxlwNwcvcWor
2iaXZxQHbVQ18OzpaL/4xlJOuPE7ED73wuSWI73MTBDtcPS66H2bhZ44WwsQS8JKeQvweSMRJbf3
ozPEyFUX0Y5y1XV8JQvcJJA7eRn1K7zorOAZnTmF5OqQueSHjUgJZ6OrCVq+y1dyqgh27ffZeJ/r
7xUf3KX2ajtsqyu3eODGvLfFZcR6Jo2OTlza3JepnM1CzEb9XJYQLlxaU5egwJVVBSHsE6GiZmkr
wZDfnT5BCUCjuAacyXMC/Fg+NjYKJU2T4L8zWT46cdEDjn8s/+VVrlr80XiWRM7YCbRMGomliMTg
qbPGrEAhCkTIiwl51jaT3VfpGHDvaawxo00+zHc1K/s8+2Akf5hpu8ixZCkRo5Rf2B6FclZeCAFH
87vTtk5siXECpAYwOJJre7ZMFwePgdCQ1Gvet9lIcOPHAZuNnyYWEkSUK0unV+gILCwVIqpgSwys
75AyJGxVWYK1zJtSMUQMf28OoNCllQlKE9fdaoYRx2nQLqNZNXarcH8mUP42y/ebj7dzWS+blYnC
h2+ukq5k+mCmK5Gm1hygM1sj4ZCZSZhRstH8xL8DUQLLfUDcE+usXwIR1czr4fe17eEt2NoaYXoL
OVtPQi21fpL5XtQttFE9zPpO6Ny2leyG8Ptz+rTLTsq5HImxJrCfOcuJ2H/F+zn0PQ8xNToS7z29
IXnDqXh94w0LvFcbxVh0rJVs2JcnItJyq5yW1pK+Uqu7xBzDDnk5u4Q339cYn/sz0iCXtuyY6ZBg
oFrmZE7c0A5zp1ZSUvPAulosOPfBrF2mu9IbBOifLU7OsXlHUMF+IDqT9gTEuq2PSn2O15Tf7Gdo
oDbSVOtJqaD0fTIfEeMjgi1BJOaK7NGvwWRjoZquaMxjKw9vuDJE2Z7aZiCg/UEIk2QmqQepVxzc
6KcVp9EsUx23RyDEMza2ZOlmjhXAzgV1cCchbyUjhX9sNE7xgbvAh6m8sX2UQPkSaqLiG2uMw+XJ
Z247buiVvLIIUNQjOkg2usP6Xdks5V/F3V1zYcYlnOFef4Mkj3Lzp7aio6J118b1NnIvzmbFyvcW
7q99h1TWaABiu4INkLn47d8EuX4IXL+xOn6+QneBQUnsCzcPcTwbvFYDZcCrNEBe+fv6KffmsaSG
1BW72uIgGEN7iTVNbhYQDXZXrV4GilB/Z2+hdR6MYmMHvnoD1ZgQukIIczsgWBrWTEWHdEt/DdkW
blPJLMewEZVEh8QOx1WigGmblugixgAGy4sMlgsfULqfWsxZtD2OGgZFTNAA+EyWSTs1vhNtl00S
fZQ9LS5rQarR0xLnhXiEN1539Va1EyAw1V3u2INGwpl2cw32h7BdDnkut5Wa9Dbn+KH6Vb1tvjCO
sPATX6IrGQ1CinZRTADhlkyINqca4yeL8sWYZZV+/enwYurwan+9VtJ1hEf0Dojxfmk9MrudB1/s
IKVL9lt4WDkhW5aQEIqhunE9fTk8HNc/FVpa065ur+eheOxESzHMNm2z83qr2bkbKVXs1gmRBQ3N
BdpHxbbUAV9GYtC0outBiyTuKc0Eo8vJaTt8qGtok8PZLRBrcbYCGwzWH5VtQcI54w0hBE0ixXfC
l4uI2UWNt34kDh/fLFU2vdRuFFwu7dDD7Xzjq4fciEsFA92k7RiCWrtNC7CznjTDUjvtADaz6/ae
IvjS0Ql3cJg1jx+DCKhJlKQFoD5ExKb+6Kb77yuF5Uh3y6Mz/bqFfEhamU43i1yOmWh1pJq2fo1H
X1QZp0zHdWhhltgA3wg/BB0LZBwtdFgBCZvqxWntt5MoQmtQQ2A24DMDJ+QbvIBhTJQXo8g6uHDA
azmMIUr4hS9X2jhEjj5hnRL0BnzCQB8XIBACD2mEd0zOMOd2SvOB6x4lXzEQ1HOSByGLqxjJn/OT
2SVJwWeNBMnnlbSmIh4CJfonJh942yH5CwdDQy4l3qjWeYfCfuHMZUnzUYXBbCxJrCV7bTTXXYTU
gXYnX4nApF5soAsUOAuK1cMPS8zdfLAj74dpSVO9tsMiP1tnTWE/twFZYOTbj11qG1uZrwtwdJwD
Z5L2oczVsLh9FOaIYddyAqT1zReFfAaSnxsscLeQKYsuniNjBet/olFR+K5NuR+Qa8ee/muOjkUz
ZSM4tf9eHrbNEVOaUFhcM87ZpU1me6dG0n8VNIQjO0tByPNAPNz7S0LzV/i8CPTTUjn8PKQ1WzwW
7DfBDZBOugw/YfJ30T/kF+8Rt6+cLEKYX9qgKgwVlH9aLq0OW65UJDkazkpw/f4hdSlD4EUdxv+g
ZxG6vxwm7P3u6bGQa6bwGcW8HcOSJ/gnpQBdeinKHfABE1EiMik2ksEhnt4Plai411Ozra4T6mNg
Z6o/F6Ol0EiT02ZQ7x9IQB8x5nuKrXk8CJEIu1yzeTt+YbtPh0nuVion6cj4Ii5ttAsMraUUPOYa
6/nYDowakgDyg3OKGV6Uf11NI4wR43BHAVX4B7bb32tIdBlVCdhYCdHmApxSocHUEJ3pB/cYDygp
pRSnqFf5nBL1sry4bPV9u33WxhBJRx8rmRijGfvqtW0HvvboW0RAIsM6swUbzbtAO9zO8aARu/+Y
A+aiu6OSaHLXxSv294fDWmPBlDivLkFsRy/5nDVVSijlsqy2z6h061CmYRO8/LgevO6kz/gSq8hJ
sD23w7f7U9t0ipUj3RQVECGk6AFP3fh9l+Ke8LQ0K9BThxkaISDSIl0tZ0N5rV2Z3Y06oUFGMRyi
+9FfFypq3N9/nEwsE3eknZAZskvs+x+sQoUhHZMlMpj/RQb/H5oEvuTeTn38veqBrUYYa0OdKb0E
4U2RrrbY0o63UgZuuI9nvqCcyXlCYHXwBEzBuLukL2/PAY8zbJEegCCtDCG3Kh/++DIgPOybzN1t
Ub3ChZu4lSTQnTdAfKcA/3hrTPUjPChaj8ELdk03JTgSkeoKh5/z/B3cxDohdtjX79R+c1CmVk+7
8jEZm6g70UYqunnN/E5WVJuEJpz//41vDmOCYnrQqW2jCtielDhU8uZLj81NBI+fnH0ZlLUH4vD2
7z4NId7R7at1MfYz1aMBJ2/UkvwIE1c1sGmEIDFdGB5y/1DQyBgLiAPy2R0KBvoK+B/XNo6PBdVK
R/eNfhaHxw/jWFh537mKZThd6ijZd1H8GOUzL0Zj/gdSsCcsk3gatCOKS0Gq5DZLlJHdX3jHC6Li
H3qHPyxy1plvFXV2a+2fqfhOytLYlX5Lpel/m+QiYIViIk2Z489SvnZLTVCpSdXd35Xc1w5kqtqu
rtnLIeRr7xpHiIlzuCre14/uxyiIV4zvCVYYEoCHkO8xoe/24RFIw67Lb9WRLb0NmuwBjfG4NZFU
OD+Goa5OXDg6MKGsAkv3/HlTFTkUBWkRYEJFE/j/4DUQArVmd/+EVBe4tRDkO3xFNDtPF8e9sF8X
RtJ/NeLZ8HA5ZLOATOJlPqFeOJRNwzOnN+HdFQWLVaIWUUouanekNQf0uOKIy/geuubLolvyx5o3
9Km6IgMr3i76+whCguAptSrT/T9Od8EKf3S4N6A6G1R4Ls6lXqdWf2lebdS61Gc/I+ASF2DwUo++
yt6qeL5SmnywKM8aRpa5avV9jVDFu4Xsvz5h6XYCwOZ3UI/wEjPqpQi/+ccqZRVqGG/dSZjQgGoN
0tPZWNpGyXBOVfMfktpOyh0kDCTvIa4JwmrtK7EUwfmH0ZaTLcqi9f3ZftlEZ7e789YkKmvMY7O+
7xYCKah/DYLZvF6p+HxvTuovLKs4UGQYsKa/sdTyDFa7sZJ3o5zPscv37l8RXsU5L5ephVpBLovh
aXAdromsONYvrMt2uFPteiUWHyKegkSkDPs4k8TVYzeuqLtLIzeG3too85jlqsEE1gkYWfYfNyPZ
sPzQAcizL57jkT7ssTetEbrlekbmYlOK8NpgpeS0JxU2XJikyafNQhveOrWMK7gcZZX4IaPf4GXV
bAZBF4zJIBUfUC/YSqxcdRiFsBP0v3VZQO3WvtzoE5WLwzAuOFhvz7K7IgxdC2HhVcJKFhOoj6TL
7r+dPwSDk8Oe0yhCbVFDFwOK7hZgd03F82xfkbnkEKtW8mcR3GpPmWNFWOKH8MBIVJ2Kcnw2UfI8
YU+yW9OO7JiQlFCpauBKIRz59VQl13tlrUc7zjRcbrcalO6iSX/Dtm4YRttXE6RKZpVpNSTK+L3f
quF5jSpDSUN6aoVI5/w1uxdsJ7QhNRqaPOJ8oXuG1IjVqHPM2so0a1bPYMws5nEvEqeJ48cj6czJ
bAxgpy5mzeMoMRG4h2t80D9pAjS+Cfp5B7pK4ps8ga04dCQFlNKSx8t/7utvMhi2MW/Ou1AzoEzY
GwUarN2xSPGiqbAn7Qwxw7hiJ79AwYnFC8gX3ayIAPYST7feuycGcO4ktPw9tZRAYkkDXstCf9wF
MCWG8iegb7tWpXluhrCYLPdgKOmoOH2xP+HmtirqcmTd1qTrwHQXue0gYz5hFQGGG8MFdhFk8pgK
AR74OVarrMtPOFkyVrj+awfVouN/vdQ3g5wTq61mmq+bS1cMZm3u35NNZr5dTdyK2YTYDn2uhoIC
vTIJG1F+MS8cY2Zzh3oJ8Mhhm1JvCBtm9LZyQKE5+OFxGau0ViHmZ2KggMcJVE1shqgq9vz15dDd
kXVo7tWRKIh7DeR7/rUo5Q4yfEiFATd9zT9gIOhNfhYgSXEDvbC7Jl6NXWRR2dFUSDWdZDEEs6w/
zkPI5UdW5ACszHjDv044ozmIID/eRw7j4ct2rRgQ6TrbO/3OadmWW/vlpQXswutl8XP4ZfZx1T+u
9+EPhbvDSy2JWr0PvlJKLc0/Zv+Oy/bFpUQCEYWqXnw4azYEKNYO4g3d4uGUJoYqA+Z1L1+USSgX
3qynHPAj/zCCCyGDAOLUi+zd8uutbI6VagdWWf704yYPOX5s/zg5bG/M9f08alKrCDtz6Sgw923w
soBA28t6iNikSt1bebvGDamG9lDDmbBmQHU3S5LRQcOj442bGGVJTWm7PiEkHCqOjRmpJhSPeEgz
Ef1MO8f16Y9mEYL7ajyl3bU6y6Vp5as/A9hiqhMNLWbk/i0v6wpfJw3amZkGrHBQNR40G8aZ21BY
46zoDZdOhjnrXjCSvbfeDtyMIeTbMRPucz+WPIEBixp7+oVB3xtbqoxtj+qP7HixdBHigUtyUubp
QxfP2N1CygtmfYLseLkUdFu2H4DTJnkr9TeyXMGQSSzxQusgKUVC4g0XL2iaG+K8dk10BDGb94XH
mhQWCDw5rn8A3TmCJRMYNQv8Ra707BiL4zzuXWrpjymUmft77CQE73HZqO53tFATMJcBdLw076Yd
1G7LAFzAHSkPKopJuMAMpORW+tqXKGO1n5yegX+08I92kRaFSwHIunoehqMUuENYJlADfUBP26At
XDJOTS59qx1rWKR7jvsVgwvBvsnDQU3795IzM4hOujg5GleWel7y/I0U6U6fr9cdksp+732XSi9h
97molBVzus1ykGwY9VV7GLnXo7diw0fvhhV88lETuHhfOYcyhfHk5WoP8qj/MrdY8sYSmp+eze2k
S6EOvohQEZ/b2ThyW9kbb4VweHSKYp9Rap2vNR2xK/8ReyNm6T8Mosl4EwKkHhv/6baaNDp0nSpI
2gKv/ABDKQFvdX8WeuuJY0V1V5k5u2mu+Azrqd5iZKjj9wUVYU5/SB9zOKFoLiC9L+qrm9v+0w7u
f7AicmjjlUH/qct0t0IGT3vBBkX59rPbA1n6uxw0vq+9DGLBysdvalx/Usb/omk2Po2wGvalDJdI
DYX6I1O9RWA4h1epFyFLCP5V5blfZUwa/9JTAyHRcBvEODbuBqgEBDM3eN6CKVW6be6+/F5ehk+W
llOBlPUJNVyGwYWe7lcPnJrlrfpvmjph0PRzsaxOr36FQAXfUaVdL4SlfddI2Kl8HqdkbHYWel99
0lr/fvLsdi1IrqvV6gfGyj3XthvW2aPLtcznJrQXT/T0X8G8wCFSFH8OW9zWHu5EBDFeVZhb2FUk
aRVVmaeNIPs3TqnMp8x5+JSqBNkv0/Vobs05RVTZyjquR5WVcxDF4iS5pfZnFFP91slkEQkiRrbu
PMnuGp0uTXGm3yHyC10MMMeRFNFN3tR9gzReeD1vlNfZcsEKIb7jFN9QfQg7F4fjDKKLrQpcoZEo
Dmn4Jfk9kQt3vDYDM7Ed9Pq/PsfL1WFtW6itzebZik/rYMxVUc7v5ZQvIi0mWLL93VMTgoQzD2aL
p0/2RDmngaV5809gJzaWBkeh7T1AmtSTlBjYCHBHHnSa6ysogbk9oVvtq/aanqOMzUDtNPzxYvCq
sLWo7RFyhAgG4V6QQq6Pav4SyFbIldXEJhO/f/NUmvSLhxqdM+0EZxY0gHsfeW+XFQ6F3SXu1Dwt
lQ2haEGO7c+R8i+5VdTkRfjJtH19hGzMgpRrBFZsvEAeY9eQ9rRxYeGRi135Kn8+3DBsVy60IlxF
1bQ8fGKY1v6qVKlD9qghCkGO6Z8MndI1/o4MeB403pA+Mo9kkDPG9/ZSTkR+qdwE7kriWaFxR/Kn
LDSQtx3zKR0QToYw9Ujq9WjioooPqWqYIpqYKqc41n/uyzFC5Kuwb2wfD9vpA11Js0ySAaNbBmRu
FoVBjs3RuPrbWd4h945dISZKV1Rx6E+eM8ssb+RZII2yitOXS/O8pTezVWbDEvss+2iboUQOfCuo
olFzHK0jFX/1JqCWrAWqE1HOX1UtKiMs5OA9IhLh5X2QnaN0WpS+FEV6BYI4Tpw3ihnCvWiXBTpX
mEMEswh34OSpngsQ80kJsheyf47Kf9Vzhvtu2qzG1Ht7ygFPTxlorrH3+LKEun12ZgD33QoN57J7
58FvYM3bG425XFfNfAAQjR4MlcnVepX9TBy/DcaNOd/BxaAORa2aFR5HVKymQDa6LQ7bSWWu6t3J
jgiTEsXcmnHayTo4EPoJUDYyIdzO7WNDpemuTVZqT/wLWt9nwCr6x8jP1efhv7w3fG/Big5JY4Qw
pdGqdM31g+oHSk1Q1l8FJfQHXktFhWxCkFLuhWkTNTaYD8PtH2fUNnEO0xm3FrqAx8/+nacUnbCm
NfdPXADdunsw1x05fqrw4h842hHP7xbxvpejgvnHR6F4v4/WCJWeHD10nWOvR43PrSR0LylTrlh+
8sQSuV2pBHUmUKgYULbnq9b4QPNyHjeb0jJVLjyCHK287HEDq8WWbI0z7AQnTubMbGI4QbxvlHpx
ybTk6IzsqFWdSKErJQhqYFwbnX4zT29E0yiL/ffdlQlEE77/0USA5kbuXylg2Rp1/HMu8F/rKHVB
JO8CYSvKV3TFCZTLSgTInmw3aw22sWV/rCyS3bIG1GUdxWxGGAqN8/iWiSNCGh9kS1u/dgsCmqq4
ERxQrQkBzGEbbH9w4IYWjYXIUBqpJuRzm1otyELz1GEgLifNg0BofI9cYPzjOd1JRmrddzr22JDU
sDbBkARwGo1Ny/yM7MflnvmfOLYv9ByUY8tR9MWxc3bm+xKwii/ENAy+pOIXPDX0zEO0pxF0scEq
vE4PPbejRQB9jn71fHY9Ca+PSRSD6I4UGd65IWjKpMB+YYVQsGaGR8ncqVMxUQx3Rc02I/TuKAFd
idGDqLy5r84+QZ4vOxfh9ea+YH91acryUEd5A+QNfjOMZw0CmQEG6418y2SftKK1tY4GDxKLYf6P
iwuU2Wrg4928tbD/VDGSg8kDdlqKHuBR7RXEiFHFWXktZ0cwLuG8jUS3bePHUMG6st201aGZ6YOs
O3/faS3fvzb1IthGNA5YTBjnM+YBebzduGH3wxn0f55rQC5IZClnKIEBE6cD6ORYvXGIGCiFNDW0
mz7QVZ0aqtJAaCx2k3e9tyGsXJV26xBEQfPMbOeoXStTxDH5oEwaN2Jrsu/p0HKZG6vSkqQhSXc6
iFt6m2fZRycgIWeD8+QcfS7x7MVUPHFk2oU84SuK6sVGKDPMtvKNowRb2mK7y7MSI8CPB9RjAcfK
Gm2usjZx9RTy1va57zeVo0KODkBZ90RQ1S5idjc4w0rfgKvgbzML3yJLQYXEjagISBE3mGpv2IHL
mpLR6IydqHbD27Dlp+sWB8vkiBISf3Tf6gJuQAbpvd9bEl0z13/hvdsolZT8bHnAdDkvLqCUs4P+
2f6qJ4oURSYawKscSjBgrw+nT324ZObDReeLue6RoM6m/B4A9QiUb/7c4S95bnS599AwkCPdsoXz
esxJwKz3oN254bGrIb5Gv7+BD3vGYvxFHQFqFKUyAtf6tpbnd0cudsPFRPOO3aO4gVQZJVmb4OAA
nk6HKCOz+4zpbT5cjkeDFcJS2cLjE1YHbj92Yc9x6V02qos8Os7pdtvB+alRq1/4DToOqmHWIw4t
zUuP2vCfAzTA4BYuipsBEB0wUfkL5DlIpV8QSsKoum1nUFZ7D6EffMzqFXQnDQWqz4dVVM9trxox
KtKIfavqGK2DGyH7fXxD+C28fU9sUaNSKqbqXvZt52hPTbrgRf0ke7zYIJgB4B90beZ4eZ2EB6Ax
TYO/XOtFUV1hFya10uxVb3GvCswSYRxYoUQPxGzIiYtywHJBek+UEFesPa+2wQXP58knbSd6lGyu
Dy/P/OnUBBw2Bm3bvZ0wpfw5lNB4vDFRnK6FnjTHnzQA2YtWgP/4GFkwXQbTRwIO9EO9don4J2+j
Q+umtCa5rWmQiO3+rdcrHN7YhzQfhF04czvEgLvzHRIAX/PL5p/0bS4kHS28w2kTAJ/kE3oKw9Ka
MZP/8Fzd+nP/MqBillLafr/HEBJinoYP3IowFWeTjLCC4osDUyXjkhPkV8GDvzLJJX1xnQIslgax
SQG0WEiyIttOFStcbCuwS4NvzNT34PDoxMHVGl4Bjl9ZfdBtluNWlgIzEGVb1ZGtPmPWBwCQKg7p
uW6tSqgMVkE3reO5qVaZCRb4RhzE30UO/R0UEt6RcYU0cSjiBYt3hD+p87eK3sFYjD0w62VLnNz0
huN2tRvPVezhGoOSxn5Ld0wqjq359n7QCCWRagCjqhEnyIwvN6bWHKO9p0FaNpWJLmWe2FA9JX4W
N3Z9/u4fvxWO/K7wMlkTa+rWoxMPn6Wnf/+cJbwxfRn6hwyK0Vkf1v2tUkjjOM4tmCFjddNHPZFz
b1ov2cK6iu1F1ZP6xG+Z6BF63rUuhUqwT+ajoX356zmG3yKjOklTU3s58QgvRZid8lS6t9M/4c2y
XO1iVQKWgIXebdXLaW+6NnO+UkOPk4UCJMcRnPggiPSS9ME8LJaXr/xYuzcQfT/4W+XgdrfAkyak
HSOP7wrXoXenMJWFEK/JRaB+AMIjqcML+16YMtQK29U9WIxEHWx+asAbHcoD6XmvdvlRN7yHaoUK
jpCP4DmFhnD0otNKrOKlSyk/BtHqdBjhhxaAfbA8GadE6z49yChLxnoolBgLPHrjxIOoF/Z7Pizu
W+D44zA7/Hos59WDjiATFiW5K6VxbUuELQCP5JCBEXrQnqi0hbhWVRszhPidwYwHbP9lVuZShS02
yy7w2ecEB8wv2rpA2Grq4izkpUHrgIS04xGqarZMM+hjDt24EJ9kGDF4W5YCVf0nILRiX59WMkUr
or+jbLnUwxx8BIBFtLsmvkt6cxwJhMCuLaEytm6jA66Z6d6QeBcYTKaBBbf4/NvfdUfN14R011C9
6EWv5ZW29fcPCLBFvxOllTCp7/mSZ3eoeT6iNF+acDR9Fi9CIaSc5donkMxUXewP072jNqZV0ZFD
wCj1RN9zwQziitkA3WBsRM1iWfasnT2VJDQHmCYyWLxSBNH36ikRkn/FrNYX6sYyUZYH8g8QXhQz
t4pwOG0Hkl17m3AqjPD/g7d/evsM27iYjQ3pvIuAKfe/nw6ogolKJnbzGs03BybacXSPai2an6Cw
+aErbVOWQ1lA+l4BrFG9UO3UGQeqV5ENPn3gBcMb07nHcGqYlWrTxnxgeG3FCje1qOU83tNh2EUl
45iIMWrsDBaAXxciKiqWywdDosYtklzCLWAbuy8ERedVbWVNBWqczy6ZzOWdoqmbkZvQYv6trMUg
nNiicEG0Iqx5eDdic/aw1c48fn/hGdJN/E/YJ61vw0UM6ZDGw7OSzRa1Nq3ABew4sXjJfzS0Ydug
nafhdAOTuowpL6Ggjg9rhP9JDq9JfTLvLRzuaWF3CpkgRIvhjaXJfOJ8gDZXmrULgwqlG4EmdcB3
4b56s2jMlWVgZVvNIHe0QMFIrJMrIYFee2d/rwubRgNeDrZJv1y5TJ5b3kHqtsm/xlnrHx59WyrQ
yZNetCEugp0ZFE2Z8jrSB3huGVUHkIx1k7l/n9XCVjWTJiR7k8adRe5z63X+covD+SQTA/o083D4
HS9tEhSFXFL3aB1b0N1ytLc5esug3TIe5vUlFsWOR0HL1yorc+tMqfQgTbHkEMjEZf/6creW3HJB
Ym9OkACrZLsT1qSMLhk6TpEXjQ1dax5ZBqPl0oWh7DowUxqojj5otEYSUJP9n1r8ClZ7IxYybCwr
mblXjYKFiEqtTzKiXpFy62fXa8tWMVc4T59fV8ExmB98lX/fhVs0Bmyw0j8r1CpwcHnAOfmriOA0
UXIs3NnQiHM4PlJwIAl9GJ+cKccXE09Ju5yQIbQwl8FBXZA7Sin/mujJSrN+gh7qIurka+3suunt
C8fR/cQnaJhxSt077dvSpMvyPUtY37H/W0KoMdfrN1wYX4Qaqti0ppifokcFytJ8XeXHE/fIxgK2
T1BuyzFtZAKoYUxE6J3yHWRXjcZrt+LlCF3U+jZIXbwZIj3RhZRMkKTdmI+KmnTY21S/wIvM3uTk
ELH678yyd8OrReEs1Mj9EK/sbQre553CnkmgFYFtgVPdPG+vh/3U2XKj7+CNYyb6U+7Krvwnchei
O2/gSDRFHyM2YjY+eRnlRUUmlVEG6Zgxf88leULx5JFkXq3tZUU0A51FCr4S1xEXKgztcJpOYPew
pl6GQ6Krsk+YZ8avcXhNEvxP7FdYZU6RONeFyHZaO7yDFOtuF1Zek7cgBWMVl2R2dwAtVnijHvZn
X1DskQ3DzCGYuDJSg2flOVweg5ws+8ur/67V1enl3iCp0j17uhmLBOAv/lTcLSVx2XBPjhiw+ref
H+d5HyZH6QRBqqm08MxjXn2rkpTFnjj3f0oV/nADWb2o7E9eLs3eos86GiEgkh1pSoY0zXWkwTAM
HjFDFhICi/UjUd4JJPTGROzGRyx79Q0ltPmg6lpi2aIQLbG7g8e8R5J0dPFq2RmnALTRERnrRiln
xqOw0VhaS/Cb8Ll4tcBV2KYw+44oQy/2VmnglGNUtVydlePyS49EYc62SOV4KzRluoRQv/7PRZPR
D2u/Z8jTvSK7PUAbXfSvzZT9v67sAO9v7IaxxtqaDMH/m93Lpwf/sFoC5MqWjKYl7ydKfBHsYpoc
aYR70PvFncMaobThmG2OpK98bTwjWZHIruQi1tOp4UElAiEgQxtp+ZAH3t0sqvF8Q0Xv3cKHS8mX
Sdl9f6KJBr0OvR23aHY2f8Noszew2O/RBHmczHpFHhp8xfWinvOrdy4wnXXcorcmSRayc8K7Fs/m
OCn4LWpkq761nrQO+asWe29zgT1/oNPsLHHuPHUTX9KdIL7O1jbAEqZhKM7T6ys0jaLqW8GrhTk/
8lddAwWTQXWhfGTQuBoyI0tWcv3xcUYwnZL5m7OZOYGNDlnYB3qV6HoiMpt3LGl5Mxjmeeu5pI0W
lXv3dQ0n+wxKn6iU6qceJbxLWy8ZkjufChdrcf+wpwWE9lBcxRC1QPNB06XIUyjxOxU2lwn/DtWJ
Uz/8hMu3ff6AOccGdMiR/Tw70PosRqUQw1SRdoxdTZAdgCm3Tebsdrow/QaDKuFOIJDxp+mOu1uH
5bdJHI8VZcp9tLj41FgQaTce8XHknfLX+UAA21Qc6MtlyAOb46V/V4S2GQ+bNaHmHqI9/cL30yB0
7BsFU1tBzSmyf7p3PZlpCQNuSdW6xqn8Xw52GGe+7N89sU4+kbkZrC8+LxC1YPQyMIhJz+CsBIhJ
FO2mc0PJ+8flrfsmdd85RXXOIAvmYLlwmBpiFFP8AeB6Z+tO1Z/P2+wns26KITmCutb9oV0oU4E5
Yxp7JwN4tz/c8FqaLroEXayBGFq8rMDyHgDY7gPLQ/KBQ+704e90muoW4a/P5kZjwhr1FkypAXTo
10sHm2V8nrs+aUQt3NXsYiBBH3QHu4rITSamNElOfS4LCsvQxN1TyZNVr6EfgyaGaKyuOP5SUU2I
SDbz5ouCGRhOHSgtILlDycvUfdMdR1AbIyrndm3tM+X35vRwpc9qofKAa4wQERO89p10lA7Jabj0
eUGKY0TJFJyoGdLzJXoZ7qEdKmEypCQoHInmwoWFmLulUjvCvlRRVMaq0usrhFy5qInuFw/oZMxI
awgO1c6qx3MOqqpL2aVD+YEHmc6xCLDcpC5TYjh63NPOrUdzJ/YCok0EPs7AplB7Ezejy68i2ej5
53Ih28BBUg48f0+eguV8+YNeT16UD7aNSub9yl1eZFWiB8noRInyvyqAa5Wf1C5hoHWdeo/VMCNP
CtfcIiciUqvLpNscgfK4aRsYT46J7qIMcUBzAd7V+6oQMANnPdIyovQfiIm8pRJe0G22deryX/XS
EJaZXiWARaSVeAokSpCGTLCTd//58Ohbehf6JHNBXa9Tpq4R6vqD3zIQ2b/gd4U8S+gtIX+sEQzv
YWYoT8ijpTQR6q1tDCmQUUmkQ9AWLFPFh/sGTo7xc18kG8nrplJD+i6tut7AxahxWWSTEreBppbz
Z30fDbtNeVhMKPxDaF49lMPd+RV9dr0xKRHAAXGP6WKkIchunnATrYc9ddyVM3ju1W6EvtXi/8Lv
Cd1SwRGGKfzzJhOk6SnQal7HcfNSgESHb/cGFHgsyQKde6mMIOuKLt6N/2Hd0ZAj9TX1JBpSJjtm
XPe93OEaal+DPG7UDjEHmpIATy4qgRv7/lJVfKIX2pLmzdSmrbVSOcQ9849+/VOqzlAXy26q62D5
xZNoAhQid+N8Nyt51eWAGbwFNY7u1LKdZFbEch493vk8FTl7idkgXE4LYcK5+JxFai1l+C+QmJyv
3kwRgwnRyz8Q1zN86q4H/Qq09fEk6KHCIk0dUZI3ZZd8M2zPpA4hF72xB8Waql+h9yWfegQbWNNg
n42R/hEGIs1C8EuYpEqmxCEaP4XQkAd843ZJ0GlGZC/a514eFlKBcN0zGSW1Uc01v//1PpZ/Also
nSaaeuB0r5fQ0dpYhJyHMpwZJbscJdNrptWOznXhowgP2o3lkt0P8Ewq7oFJbVtiILuu/3t+/PCP
ZarpRllNhLeqP7CRXx1YebAbMGVTMxGYkdSuJySK8UKYCdGZvwbPPPeVAovhXsxMtVCJ+lQ3cuQl
yN9mYOXn7jofXjgZSCOmrDF3E4NS3QVGN3wE+/BB/iTqyWyD6tgi0N0ifqiHrvvHWrf9AdNUhCdg
dxAZCTvJhojZrSURqggN5gjo6YEbEd27UHn6yvCZe2Y0QdjMSIzSuYLReRLGFYLvspL7lehWnsJz
zkiXsH3lqPhbdh4IEcDLWxuUS4LcTLaj6fyKRDwXL0Q6yXno/wRY/X4+4eOqoPtKJOSoK/qbvh9P
jHnxJGp9DE9f7gmfGCphqtzeCwFARe7J0Km6ZEE5DMKYTdafS5oDVLgoPDHHYw4BdHk6xDwM25Uc
7FIVVR2psGLPepY6HfIw2y/SCc1RONrrzE4qM6PLFRVgvkHL41Jw8mxB5J9h84V8OoeGp623YD5u
pZTeKzen6875h341yl+RhecdU8vxAv6x3WlXlQoSeHTyuuKKMMAnAOssnoLCx0dmdjdZBVoXRbz+
Boo4hKDZxACxH3GLsoKiUI6DqTjgguRAEKQF0emFeXUNt+LW4Zcn/KVJIIrv78JrcaHjLYhyViCI
6PtR2UN0A9NkQ9yanGDQX3iRjfAl6oDGw8HTwg9KQ+NdJxvZTprmDO5MrhwbCmGcmQq/hbOKKAqj
np5Uq7EGwtNXf50176So4RiuQaBs0wO/3kThmdZA9CcVftPDjFA1Am0xLAcC+6LFxKNv32RnxlC5
ypDWWJGrIOz1xGtP5LM70YiKAazG6Fq4IwjnLbVAtzC2CHum4TwvvgPB6rehbH+EgHCA3ug3/LyX
Jzp4xt8jBc7sSGLwgLh5PCeOZoEuyRcP+upq5fRacVKUJH4c9l52nlZfy25E5G2vdSBoh9liIC45
Mx0y/ba/ogigciLMUiq9S0oiGJ/B9AvQO3XrHfZidzmXthrEhqQUANLk7ar46iOk4Dbvryq+nKyy
5aLHJE7pImmCy6TTlGleDAgC2tBHpBXuHB84tH5tDHZbgPl3pKKJsQBJf3U2T9D4bwW4m4MXL9HK
saMd7bbCsDemER12TV0Rh3QYYY/dk+MiEsHzMErE7xk7N3pmZodqhctaQE9KgpN8gEp1knAxd5+a
WdMKg4xA4pf7gbHaaGVi3E20xtTaKJMst3W+Q4EQne9HdOGgkg9QGaz6g9peLDzi1stepxhmrxRD
Uv9ZIZHiyoHKG3qSTo8AudfGfuN17ofy0VoX+F2PBmCp2t2ecyoC94OshBd2TgLcrpz0ASQQa9d9
roy7hyukd4VKqE8/PQHHiwAwawCc7CT7dvnJH4qu9soy7G9khsa0ihRrThpa+gz4DduC6gU8mVSg
tN4KdGds6/VIFPkegvhNGyh9Oo2RCJz1zCF22Gvd7+UseIrPq5tEoBU9RRDo2+aBNt4NPXZesPXg
gsKMLLxTMJrs0DNJ7GPEvWFWCpAPIXlZD3+N5FyU0oRX2zNM3mfINPH3644JWLKARtwsnfhCoOPp
3BsEoE8+CXV14I2SAmt4VA27RB8LH2WgBIWwOj9h/56nPuvktisfKNE9B7riXQqHxoHKw26UHATE
mwRilv9on3RaHeMGXLtU4N7R6o3uIt7y6gIRtu00BH4/+sELEEJahRyuQAK9ciUhabhkVpipLrbf
XQEhL0R2K/Tx2ASwnsQLNwIZCWaPTnnQxnsl9TaLp4JxdjtdLvyzwzM2Nu0X1e3vFn1xMZbWOHr8
c8LFZYOcDHGVSthBiboIEHBAPQpdFurw6J4WLaYhVFOteCZe42oSjwTbgO7+HetkZryKlUq/Uip6
KzCxtg+N9MyP/ww504Ers+P50+KrkjhjwdXTCnTrrmP8JwBo2/1+4y5liy9aF67ZxfDEoKEG6BPS
1YLDyDwYEhFC7v/ec/xy4k+kFIWrtql7CtWDjdxY2EpZ5BZz23Lxya8nA5oFM69OeDdl8b3ZNwUY
su/AUa4+mwXcFa1eW3TBEAWjzDgCyfypV/ao7WFCBs9EyszyMCoenCr+fXfs3hGlBufdHmRBG1U+
41YD1TDDv/TbABldT2ymhmSNkuuG/X1i8fLMjkGFZRaOYqgaAj9UuVGH1uNdnYGvP0gMUweumryb
q0vn8yEEUb8NCfmbni3oLXIriAyNBBbbD/7hjEkNXhJbX56jfgXuS+XUtFgiuj+KSM4pSOtb+RjD
aN3fenoiZI+iGg7+XNOt2NDualWr9mgRs9ZP7EZBGvg5rDxrmBzoyOweRSWtpuO9fuyybntOtn5a
QRtXw5VjBZX+GzbWaetZU7JjxuCgBMbjmn41u2yec4Dy54mavqjiDrMtVMdiyEbwuS8zHz1H9z5n
FaBBkT4hRBVZCswq279Vav9ljeSZO/v16G7m5yseoCtkiX+PM9i8byVtweyu7T8wOsoR1MP2jHY7
c5naXVGY0nnHO9EvgFuODxI5jNfHu+zy+BBYsEbN5UI9TV4s2oOBjKeNVXxiMuGjG2mdPhy31epZ
aUuQ8Qs+lK5hcQWQjEVHZ+cut0HkdljOm2qolqaRkNxqkojJawK189JNwpmR7M0lfLYahE/fKRwF
iJPUC3rOtAQo5ZADdxsHAVtem4p8cu3lCFhxldCC52Sh1ol5G+LSydsZ6UjWXRqKsJa5rwBoNnRM
9ciyKNXwMyBPaQLBV5W6mB5vTy0WIH4KUj1NAGpMUeqfAwJ5X3VobaTYTDOIsNdY3XSbt8CsbNKL
LCUaUvj9jOhZWwQ7YgnjTNgm9gaPCwc7nRvaZgNq05ndLrn9HlrOmfYK6Lf2qmfyhB5WeHBQDGtv
zrzk7pGunux6wWzFZHCo1ugWZUQmd+IRhLN3CrUGKF73nCsBgbECrTz5BdSUerjdzcIRJ4BJWwvD
kCgsNzP1Dw+Jr198jSYHYSosWTZEUmoYEgg5WYcSwTcr4eyErEOYvmSTNxYd6GUO9uTXDv8C9gnP
5Q3ARb1YBbIhI6TEzadiRmOl4V+IMVIw1AFdvq44U9NvET9/vFJMRULyfFyf6wrw87biq40I+s7b
nDPiSXFmqUPdGtrjuLWmU1wIIsbC8pjGIO1nkuL5UxWtDFLnDc9489OaZRFj1h14NacWaGXDhTm2
VDVpIMOsXFZtTajIz0Il2sOyaGMXi0JNRaKqBtqyw/A/Zz0T0QSYAumBug3Ex45BV6mIZilNJFpS
ZZXiMQihIdgVH/Yqxb1H5xlKZe2j9SXdIVqyoFb+fS1QLa6c3XgZ/jVKB7rNap2jMyek3GUyH9ZX
rWvL2zDHMvYhFlhNATg1GPbFv8DY3bxtp+XKUiCYjIoQMppgAReNKmXLGybGQfY+lyJoTobk0+aD
x4TP0u1HkBskB5wQF59Bh75Tv+A5hfwkduqmC34Y1nKItl+B9u5uY0Y+JWMTXx2fDcblIiO7RLjf
DopfIyQG8PV42rTnzR6XJYDWwlZUSMQV/xP9INIQgMXx25ERyMhlanQFFgHwwTXhZ88VWMjrXVzO
TwA1mw6+o6iCTlxU1mzymwH+lNz8aVIESAW3vHaCONV0DSmpxiAx2oFyEgSeXQEixPi5e5wUlnFk
4GjLfTooYkfSS5UbGewrXtx1mT2xzIR6lkDd5YgJVlMVQ9dtzoEDfJzAJpraB/UG/u6IVTGgKWki
dpDY97xJMZqb4IUSmEgZPLzs0GQUL48Jf4K7XIHS+uodmU2bmNYFTda0lHLO3V+Gw8cv27hWoz5g
7donvJMKCL27Q/AsfqpKC/U3gmWe6sEU00npaK7wTFUOczNW4auyXDFLljWV358a3/kZgaPZbiHH
Tp4T1XpPfK3wbvqyoVFpl9Ll0f2A0hJUv0xLrLLhN4GRpurWQDjx1mPSRGaczsmgpLoiSfEcwJx2
bZx37dT4PZXcdVRdbJfxksTABeNjDODAJtHDcTWijx636nYfZrGriwtiKLw3ajQPReDUFriVjUNl
qbOgIY49G48FXijuM2C7q5UEjcpl3CS0oaqvNkVl0oQ7K8QOx6oRMVNZl7LkRGy9AxCruygpQUT6
jfOBcV4umLzNfq6Yl01hT/frdw0UIdZqw2B5W86NQmuq20QvbzYGkBXIbQbT5ewsIrNi5VGs5spt
KMI2irWAEwaxmvJ2ldSyLT9Q9W5XWahyqlHBWWtcl63hQo7brFPQ2Jl0WUfbLMwuoQQRuzcHpilb
zi3M1cpy6FV6eCmbrdfhyOrb7n90rm0302ArVXH96dAphP+6k8Qs5kpAHxFaWWCl0CE3P2fiaQUq
C31FxN47E74ZWw2/GBB1Pqk5OAeTdw5HtwR/MSVFbaEGijajLyODdywEUmXYefz/vBlqKj0GQ34d
1QH7o1+9dDApr3N8UETOetPMwWats9txHzVEdsjB24nHe6cqJeJSejL7IE7IWNvu10JAw/7KAq2U
ecHwnoL4/P31S1pyyerFBSH0OXNlMGI1Sxa1AL6hf59EPrEWmnQ3LVctL5rmblVzssaR8hDb005q
eJjx7t2rZ36VojKQLFQEmyn6v5s4uq/QGcZuhhEhFdzpndqQln/iAeN3fbSlXG7cLH3ALa6nF//L
esfGJcInpi958FFujjN5frodszk64+swgj3HYVyqTv06TJL3Y89AKSwxCNeAt6YcSKxZlb5E6m35
rBlD02349lTInm6gMoshrZwPQeu04vLgHbPP+SMFQvhglwlVnQCNvkD2RxcsuPm82D4u1kh1kyG5
ODLMkFk34qdvjRvi64UUxrklTcMqjoXVz5+RG8ZNxntBJR6UQrHtwME/TdVbKHkrywPrTw+bkXOg
B7jtzDy76YeF0i3/ow33Q4/WbIcTvY4au+ikDb9OCAPjfheaBv3wz9gaHVD4sA2G8kpLHZvH7HyC
ShwJym+mPoWJZluFKaoHdoFlZgSbdoDInFzAlcb4A8HXRY8509vCq1ypimtF5GHoYpc5lVVB6jbt
TDP96nrH2O5NCOG91E8pmxv5jP1A1d9OGv7CdD2J7v2mxXaFYpyiGgVDzMJ1nfDwm2l3xwnnxowF
FupuB9WqfPauW8BxpZyqPJxW6ACOGGm0ueN+rDjsI8d1PBK+wW5G1ErcKypIxEMMv5Ad9PRxiNtg
Rr+4kPaTKg8eZaadDzUzLKhGLkVfTGrB6Hw0M4V5lLNM0gv1B/i9oZA6+FytVl15uo4QUmVRVzlx
QbRdtdmvWe0GUfb67bnrWtVR3KqhbZPZrmpmoLkzMbHIWcDc/ABjSGPodCy/b5R1Gs5gDSI6rOxU
coW06vg4SDJDZmZB6uet3MCikSCs7FMUdX7ji72C9zFHiWw7jg9IFOvHGGGiDe8G2uzxXLABO1/e
jG1upRTQRlM3ERFucvCDgQ7Jq0+fYSkxGIV6BPKjszdQ3DK1e8DjZZQpJ9HnnoWOjdBzH7RaprkZ
hu6ZkiFNqAqxSWTHvDsNjaHX4No3zPzBRPiEuxS6GKz0Z2M7aiyHBw7S/z0fPwRjQgKTTevlz3fE
C2aufTcaz/sokThK1zEbyVOoX1F5wzhEemhuxhuHvjmruH8hRWToCf3gWiLKc2dy8HQ+4PH5OOZI
KNZco07l08Kh75m0kmVZSY588FnSfR7DZWXTTsBvbXDtQ6rSgvHalrhOenlpLVPB54Ip5zMpBe69
OvTvJSKcs8i2KIqVyQkbyRUaY0KxnbbW5riUCvqRwCbBqPNPJLYcbTmQeRjN3zqwrnyQLwsmydbX
0gyBRjlK5tJnC8lApqoh7XsYRHmrdhZYTVEkxdM/reb3tkG8K3rDBPXuqAjNWB2pHFY7YUtc7Zv8
/qKVoMZl2zFvYIMpsgGMhl8jaBA/+F0DJcHPX0496ghtW4pz12bMJ2Yg5mGrPuTzBBpZ9HYARJCR
x1Dl3YQiuMV915QxWRFLVNzSkLPE7N9EwEzhsX2E2fulNWxpSarBW4rVuD3p91VPoJBaCPJ0OW0M
msfcmim4a3NbhGy2vD1p/scVIw3//ZiKe3Be5R1N9MZCVy+HeBpzguE/ApziMMSoKoGBPao3lYRK
4bI2hN7fjeFfcxazj0WYAuyN1ZR9VtqYuwIAyw6EmhlN5QP47uX4W2VP3lFqPRa1ArSPC46Ff5YB
bk+X2K5ElmgQApETtvSqrAIH989qreaFW9h1zYKmSz+ZwM7LxllxTTOX+p88OAU+qyMcOOrR9DQm
8vvO1B433Wb7HGlQ0FneHG0h+3J1ZS5PohJrn7xsQIggw49SUT50Qu/8KOrajBps34YcRo+YIdCn
5A/o99m3Gc87dHocUncbX38E74Nt1EHogYVEL8HSd0kJ6v/Hev4RMQpdEn0EwDlWYUdj620/foNq
qdxJMiVkLsHa2TdkQK6Yz/IShqbLBr/URTbrr3p5s1Bt5Mx8/ec2BhojSoYeJhhsEX6RLkwNqw1d
J3sC3sMTlTNED/HLDSrllS9EOk+h3+m1TIB1tUV9CSCwVdoUpkKgdON2siPeth7oKgyld1c7wH3w
DiSguNxry85xsPFfToC0uqqqw1Aw3tYBkL4f+9L5VKsmM9JydaeONZ+T01cZl8q04A5UizL0JZFR
ykvD56ADhYq3S1mzWsoWIwAdPlhyOt0o0fRtnhuHf+Ra2KYP8mC4w9VyjhTmboGRxUwkLlxxHES+
kcV3RuWX/E1wDntiaIypw1IQGEipT82qPsrpOfEBFwqmmbtsefO/s+OsGQRmcUlzx0YLgJv4iqKc
2HQ8L+Qkz80+CWj8rHfDNHMLWazp0NYN+EsLPmZZLo6LRQ4ct2OTpOKWT9TDRUdsqwu5kuQzOYdO
/iRAPpBoJLr4pBjzp/qHJm+D7MWSwpybAdx6WGaO/BPM03Yl+T0gQIBa3F6fvwypbooIehIZOQ+a
h9wqjHD/g3GO22dkVqOmFT3vZPyFtR4Kkh8aBKFdn6fGES//JH1oLr/QUy/3RQ0UCMDYP6k7xPBZ
KQ2ucWiTNoNE7EXP91N8wTsoBv3GK+nCEAl0KwTSe4aWb66VKhXHhOE1+GHvplA8RzrpA4pRs2Xp
dsQkHp+gHpXgmiuvHAVgZTTkxv30yf05HcEGV3K4jUUa2kBCvSMvlk3Hi9M5+DCLhZ6t+pIvNYR3
ys0dYQ5UBF/ExBoHk/OzTIO4aK9B2UkhqDhMvtvcQ20doVP02uX029o0tpFvNeVmLSWLv5w0dBR/
wCVdt7jpYYSUjsoPZBdQeO5U0QcgY7LRjEazrMwLMenrccYDOk2PK3XPAj7yT7E4A8o/1LgqiEAn
JObq9VyjhVXmvio7Jhod9gP59fqibatxeuQa6PER1SAkvPC89iXD9TXdl3uAyKsAywlbtzSvohjz
EKBWnFt98/2wL5HRGgsmhpmPDas24fmqTXAnmt+SKksuw3CZCBQKvH3fhNFyykZMLAwUP/gg5Lpt
d6at6bDX081OpE6zMfkzv1nbpK5Mm9ibdnII4EQlT3l/hOXjTKkffR91mEivE5A7+x1Q1NwHbnkH
kLjte+MGMRfhYZVtYQBlQQ646QuYKJgVcdGIkM22dThsSRihWTQ3AmfSONlyGNXB0wyloXw4vjrZ
dmnDZC9/gXuED/cnSpdPiRA16UG6GBVmuIRbhEtWfLZ9Zsz1iFKZCmG2YByR0kLzYd++muATkvb5
z6l2YIjkPsPmLEKzR6NEJqGL0hanKwgO1+cxwnWWZUIViQ0uCGhYFsIZRpsMMk1ysWKHtPsmnUzK
RLVY6rP8DJf1pYv4qOuaY0zZlTx5ogbNNuKJNfeta+cbuLTkN1CHDRTdqpKXxvRX7wn8Bs7v0RvB
aP5HC8ViWkH/m/adsZ9Az5ZNNq7PwIDCSEEb4kTFlR5hMXFwo+E9lHWRbsnn4WN53nUSOfbLNokE
ozvg3d0Ne1KrVTVJpb4zpLEU4oDE5Xbbnq+/qMwP/DYOz2nGNcrEsuFZe6wupgZ/F8q93VQdunSX
6EryHskQLsB4cn1Ee0qbNlR9AM7BWQ3bdVjJGpwnSLDLUrDCBUlHk4MyXBlicqZPiSXmBMyTmriw
uwdlZF/+Cm/MmsXJsUQe5DvzoSnKZaoHkY4uZqqYO4kLV3glGqxu2vo4/wAMK/t4/z9rqOeXIDuZ
ZmvWKxRQhgQoV+KksBpTDEk4q/g3uwUQJ3JWCDcGPm7VT0IOXSz5pWQ4SyouSylCkc5OlW2WYpuw
hLjlSVJlJ4meDmUisx5iVl2WQmz6EfbRo8cMmINxdNpfbabgLcNbq706VUaLovgLoqKLXCzPbb12
inaHvrxZ4UHRXx+FgHl+//+iYz4kz3BL4B1wkeHlX9LXqjlGEKjX7DZx20g7+tEU2jdRzda3zLUL
+sl879296+L5WJ5Txyvme1ZNGj0LDRwBNo4ItTkNwQSs8vBsfaj90eD3ddkTWnvf4EpGRVOQOyhU
bWGSDwWLWyYeM+oWPOkQNRiyHB/5Ap7jap3as856X4jhUH+4DFcOQMy4sRG9vEcRltQmQHssNlQ3
yNzBaI5/mdDHFGkEr+ErQ+1zhiqZA9MFf6LcLIypxwsTKaMWCfi0kFdA8yiPbdBIqdGS5Qj8Re5H
RQLSKvzSHKBB+VzMMSGFkmSXkjC1yUmNnLLT736AC69X8DrXoz4Yk750dJzxGFlAXSav+BRB8yDM
GVB33KJ/Gpluqbt5PNs+9ZjgdiTSDDV8mv8j7+s1ga5dfx9XiahSb5vt8ooWnSvwWI0vp53gPz/4
/DynDFRNL3/kTL2yyY4OhzfojT3ZSLaXQTQsH3ODVBzg1rzRW8mY2Ywh/2NY+PzXQMB8DIwrwgAB
cTFfAntLypaJbcXXdGZD+6tUMmaH/KMh5opXJeKY+/7GEg5u48a8Kd5yMo2U8j3jyTzxjNhAIrZQ
JJCVSxWXG3xzFI2Xx9QWqsVSiQf1UtQZIHTe1PNOaDPfZ12KZSbC5FBnnZC8YjQDvUnHLGN+tnzs
tiuODd3I15k0PocUAqzCmjYS6WVXxKCWMCfXDTWzmM+UTEFE+bzd6WY7APcD7GgolzUxF74EhkTt
1bGsKDSv55vzZ5E/TNPeiNwz8XqrzN0Ba/1saFSFMnwyghAglPECSukUnqabR1K/Jr2LcnpgRtiL
oZB0GjOUhbzFaHe/YXP4bPpUX+qx1PFQFTmBoflJCj43yv0T8+wstCyChtK0FI0mL6V5dNIp7gYA
Z+fPNUxPxskjppLfDq+I9QcJoBx9km2Z1xSLwtOgkRicyj8Qo/XB0D6qn/+bxyyiKz9TO3cXuwUY
1UmNnwH12eDTONbB3LBVkxB7WpTLRYiiEJ/T0K+iXfERpoeOTKx4Q1cvKbpW8FZN/pDxQDdzFKnX
OEAkwYb0JDlxlp19Gf9bKzD/ryrtfw8HWLlZ2HXeJ5RW6r/7V/D6WGp12XWy9dhMDSWR57m/5PUA
vQKzqSnyHxri3QwdaR+T779hykGsjGG+XsKPqYm4hW4IUe5T1LgIlHkFdfQvitb0w2DWY5rq32Fm
5GXdVIL+BLmF8QdBsmzM0o4Hw+KdnfoSPdhU64Mfzj1q5aUDv6q3NdvxYAcrQcfvzRTarYuQQtWj
qqEuKt6XhaSRa3THoVXiO/7PnPE4bgliOw3u+Qp/qBDaPk5LwCbnLP4vADGzb7vXbt0NK5FHr2yi
VuxCGiZThGMtkOVBo3o8mddwVi9ZB6UMkiFwj/hL4xK3z7tyrGoXG7XyX7jJ6KQqeVQ8XBYmsJJ0
1N2v/0YhhekW4zf8ZKlJf6+3aVdY1ksD6iBtKAUVuUP6H4GJlCBFbrJ7k2Ki/tnRJuBKS1mLlay1
y8E5cSFAYKbUke2tVpbzJ8MlFfuDj4dH/Vwk7rKRL987mZLYOp1G9oVtrrKQXgpIsxpYzJl5j2RH
WmojTzVr5kFcTcOTuuk15YvQFMqZ2ZpYy8qxgIYxE/MUNv72bl4FgZ5X5NxGYK05Ljk09hFJ/pQo
MyJAWLR9BomMke2tKMSj3GE9mM31ZMGAOaSaqX2KDKZcCdJkAHOwAGNyH8RbMZqc/LVIRjS0zrW2
MePQaOQO6GUEJD6qKr/3jrrdWfOqJlgcakWs4YPh2Fyt07CkKkR5Uw9+4zOHE+t5UNlbiva/jReq
clTHdYcPmeGf6Hi0Su85c9Fh2qwiD61jKEIvFnU4j1whlCTIsq4rICCKOtaBHNY9qYWjbMjNmZna
mqLWwSrBVDNAaslf9XL7c1RzgK5vaN0JKRWUifiMOEgJTs4BDLobCufxNrOa5yJgegdfouzoFbWJ
mpQOtsEihtf5lVdFlQ2VXtE/8D5JnCZ4JKwlTGsm8VPmUZ7zgzvAjY0x4Dhik/HB1WRObsc0DBvT
cKZmeniHpIWBG7H6EigflTWVGK8TBlVe9q4rQjiQP7eoWdkSspfL5LSd0zgOsKvGcKbDkC4qTRc5
zrXnkYII4L3o75UVcj8aCSXQAPLm+2J1Va1EUrHhNZhWEwtE8LHlDnqqnBMCmVe9O7BtlSZ0bpKp
u3CtoDIYOqBZIso1yQAytwyjfOKluAFz6SP0dIFtFGV595b+v7HBcQI+jstdJvvj1nDY/9+J6w2l
2sYxSk5GLYA8Vkkyt7ul1h78/tNfZfJ0VraKTErdnMeKUF/RYRhxLuZgqISqFW5CjVkSdHogIr6b
YPT1Xpwc5zM9mCvG/gIhMZzBo91ERGhnwj3qgHI6yX9x2TmuKKGP/4aNAESo9cwMvvOEbLaQ/jjd
Y8dYeJnsnMjPQrYtegQ8XXS6v9ff/qSXDOOVM3gfk/vkLWlh0TncnNlLkBXWCmrCXrsp4za7MGnl
3zHx6qPcG4/3N5q9R4YGLqwFUcx2uSYhIco8cbNVBxqZSb4cNIO7nalNqUUp+5o/L55BpsAhtH5H
DwEoUCbWnD4WYnyi5+72TQuRAa/kywsfuG+kt2a07CsBVy/JijkmxE+pO1EHoZPjUyGu/Cz1tHLo
henLnCdXBk0ro814FZ2Ldr1Z81py/GBsRVdmjaC554KzrW5jTg9yl9Ub/AcsrCXv/EYufM5sJf3P
+lPlU4qMPhZaeu4Mddqxttaj1NbG/fuR4f0GyGb9MB5NKSB3CvKhrOY4LiUHrNGdLlNS8c6pRhqH
qVMr9LVxeGVtyPD3O8YkQfJYGS5YRzKyivPc93HekcA60BrT6sUR2NquuggQfg1ioxBOSnBrUYPh
GmWTBNrjI0HqK+/iuJG2zmTN7Cx+97C2LHu1TNbRp+4caQSfEh4UxARGeZZvss9vr/RgKGxQmuBn
X81Y5kPd27tZ48BT2Qp1viUBu7cvELRvNnUjdy7eUctyCijYBmg6l3d4wV9aEHWQeH0Eg9jSwXs0
MY6m9g8dTC/YACnat+HxUAZ4NiZ47ofD5w1OuEbKV8jPlXiDDCr0BVzpCWFY47sOmvksYGH31XcY
kapVgUUMXjVzIm8zhP9/XiVFdeGXdr8miymRHA0pWgFAq9jnWSoBqIWQaC2AjjCua/BjCUrdUGF3
cMeH0Q/faboNkOMz8UMCN5OHvl+eu2q2/HgClDjwd54mhahCaisl78ZsfLaR2ogOSjCvUMCnSda0
JB9O6pI54tEJtfk5+5kKjuV8Uov43Mi1z6WPoJmO8kSObaznRRPbL8DiBYbDCe5QtH7Gtkg43Ylt
DaqYA1WclRNUAw2eD6MzAi4qbECji36PiFb4uz1sh9LRREGCSvH/rUxiXazhleF0R9q3UyEw7VLB
CJFsJTaMm/ZsXqU/MlyEZCCxfMQIoQytk26N6XlhtP/3/X9Lfrf8fz4a6BZbLV4qUCPixkvD541e
JrS7SJytNYrD1qB6yoi5bTeBzIwQdgWczBRBCg2cuphRodhrtUITM2Vd7MQK1uruaPm6OgkO0VAI
KBbRQHRjtvVrolOX/G+4bkhReUIRVmxK85SRy/8XbRAQx9JixflvzQ01xVWgbycTnF+uvDq8yRdr
toRwVfbyYYRFB1t6SyHf3QXTxRtUEOgcxp9adUFL6t/aG1RrC+Ds1cUMpy9zlb1zqhOm6g+RvM/Q
35JtFGvIz55iRyPm8kwTdmYAA3hnvvvdnK+1uI3O53U6M5A2HpXgXe8vsSemYUE/2lPs89ZKvMmN
KXTlPkn0ZfOKsAdyHO5dq7vLrZAdU23xslU+zCgkNPEG8FoDuXkKWMMNL82BIqBvWzL9TMLSjhBC
ku2rOfiNBrb2RwcW3AfHF+PsNXNoB2peI0Y+dX4HNR2GnZnDevrkxSVm3A5Znc2DI9MSkNsbayNP
5q4Crh6R0HgNSaMEFErjJiaxa6rzoFH8CSsgsN0+a1g8qhIIVrN5m6Jt7Ti3B0KTYO/7WeNLqYGm
uZUpnhudRlS9bDHqmveDHUVA94oNu+0FOpG8MOhlSIeO9FZc1N6fUqrKraHfv0afe8QyBJv1KrYK
wJd2uUqNIQIdKK4n+bV8xpvXuAjjEX6RNvm1T1zlUfSrY3PzlB34oiYWjxTxi1saj3GK9Q9p9fkB
MdETSIUKmtTsomM9gzzAqbd4d3smR3ZaKWo5nQ0c9jQxqvYM9FtsG9qY+GXcqkm3HKCKn9pOQ3RA
jMW5IYfolYXBEp4mDWLrsmX0uEnfv7QZ7pvA/vGS0b/C3UyokLkO17s+wDv5nyqdNmoKWt10m1On
eaEVNP5u+UzAI/O1cAWcJQXQB1XItnVUzBbGa0wRMw81SoFcD4uBJ2b6jwiT8aX09aAFWHSwoAEo
trDMASXDjKHLfr/P1EwY3UbhW604T8x/AkYdhrsprM5kFDyCZY8b7TW5nGPPqAk+2OPjLYKtIYWc
GNCHnc6rcJcPyEO8YHX74WXbSPhjiBKjnSQBBm8zpHnjjpU6JCEWshuFnqr4JFRpRUteYrgQ+IlI
BrCES+ffG3x4gTmzoxPtpc1+829NGeGbY4Zs4hcZo47dAaYWEC0A7zCA/nOUsZRLdVV6kz5DwuYn
CDiTf+GDLyEskZTlAQQ+S0NVnOs58a4ONR8X221BYCRh3RtbrjVhkejGqeozkO0fhfLTsjtnnN/Q
teidkqWfhRHLv+ySs9MFrEHXT4hufASvoZNmTfweu8oSpBCD4IlRxYgRDh5yCYt6zBjJs1N67Qao
GmaJy94oHqJR57TGsNW2IkYJOECppPus/HPyjjSTErmPhX7qQH+rSmKO4jW7srmj07mJhBUmqDdI
BTzpsO9NuRYTORariZsDPEOLNVunAhp07KMZX6WR97/xdS/Y2O8/ENIAy/2lIuUlpXhIpU75/7uP
2KkhclZSEyhdhnaw/jMZBm7POwk4pOwWBZ7pgPBz+6REXFjubLETJ+RdXzpINBB36ZZ9OQU0Byc3
INKRdn166ur0KOveQ0dYvSHBOIinwbAua9QoBmg8AQrSsFh+BEAdAg0jH7mSzBOPuSAv4QUcHn6v
smhzslczWEkgDg2iRSAFMmGEqVR6mRIFiVTMe4r9f6IE341XbXdD/hMtd2tRZUIcCCcFBDq9Xqj7
vEoLx25YMz//gsM5SQLb2bXkSpts9dW3MP9RiygzSVu+OYrEioGomQVLBHbb7OV/BxHwv8epW4J6
Bq62JIlDC37ZPfL+DRcEEfcSB/Dw1x715THZfevl/bXRFKFEF40SuLBbLOP4AE48j1gaDqbIgQb+
kn+4WMECu8CBx2741Oab3duM4Zu0FhyXVNXgWPg5RDUvLzuVz36AyNjQuUOBP9kqTvelkr8chjKm
XppbBS/9ry7G4cIEuX+bGcLhSrTbvgfqJZci/GRnMukm6Mk9WdC/4U99g1xA8LjaLxom5IHoraMh
iYJF+2tu04E+ghSqnT/rMXa3cnUOpW4g1JeIZbrRG7mehwalukZX0Vtb1m2iJrQnVNqHUDmz3wDS
LMGqxuVXWppiGN3cHzQPFPEfpJUgzr+PJXHe83A/oDuL4ybfXeO9k3V6WmVEPm08ty3STSkFyNCV
qENTZrAxS2gXuMzMXOLV7+5EDe+0YL8XliVOoOwaNyshWjBcktAnSFrwXfwaHS2SDOmheylq1bHm
8LIQIA3oahVC5IKCeC3R7OBBTBAlAeUVY2wkKyWvrfNA4+OI8qjT//HNhjfDI+oWzj/XN+ZjRkJ8
u2ngsnCjCv6PmNR9+yqK4+Fu8NS1xsS8UHkjoEUofPXdH8eDezTUXyEHuPs5fp7BT0QJzpHMH/wW
lc9Yx1DXxF3+rjw8iENHk/lU7byYrOMycsg23/CrocrJYlMMnhB0k1j4C7+7tPGFOgmAMDaoRqPV
RdNb8WL46HFOFj+v/vyE9F6ril3ywZKv39c9d2Z0fbN+Z/2mpyWwExhtZx8yByGPSwHCObGREUp4
raEyC+f4wFajP2A/aWARnGB8yKF6UWQMk6xFxofHUtMImoqvHmpNUFsm1fnAdkNHTxpwYJNEpDhX
tt8oKdZj4eqZ2FfehSYUzI8KEa4ELwHTf3l6JxIhiQIYhLQ5y8pnO0Z/QtaOWOs4mG0Ltq/QaPja
a4zMRKxbFWym161nX0v8dzr6tX0qs9tUcPo7j1nf/pHlN6C8FCT30Mi89j2/Abo9tsymItQ894xv
Yow5WYaDDl77a2dQoEg0cbOjjDJJmRMAtb1sfD44xxL8DSHwR+5dz+vR1rlz3IeIe72O2xgjR06k
na7mevWBnrQDWopkb5IxOaeNrCQQRARdd7qUo5QYcytjttp0r/sdhjy8Y1eOZA9bZphnxo48xSHX
+pD73xShw0RebdhzW5jgMEowbo0CSIFev2/wApLdzCtFtSpTPxSo2fJ7T+8H1GzY/Nf3DVEtSys2
tcahDCryB+KcF+PC5nj+r9zlsU6h1TagFI5B9pdwkDTNJI/jlUGMyINq5C4Gw1RE3HWIV/c1YYx+
YW14rzQQei/wD4u4pSBoaaiOnDdNz88VMH+R08o88wpaipDjvdIJOMHAX11BOmnfjqRmD6kuRPHE
mF4py/lXcGdHkrQrpH3X1XTKLTPnxD73K0DjbtOn3+Rb3nmd4RLQ5/bAm9TMvxmQwQgChcE6d3hZ
jUvmglmKKcw8L6aEVNi3l0nbjEGIk7HFZ9m7t7tLEwtrd+V/b6vNU09YCvHtWcZ1jjepUofMl+7m
hQOm1pYPhgqlBEPCaVuE1HHgFYX6q+VEQcnEj8Swh1Gqw/4XpeDAIlHalYCyIQXiJxpUdyTLnD60
PT7Glw7HyJmiA5xICkKDBGQjihqYR7cio0mIRJENhbY1FQEeIvvIYt2StnwtZX0eKlAIwGjvlg4l
HjfMc+hoUVUu+lMfntunxQlVko/cniyPz4RkxWBdVOF2DGAD6beFvsteFX/MCPD5fLxZaF6pO+WM
yX0Mcy4XUkZGV6MqSQd1NG/pUNrHhyDxAVXIDTeYBuwUBjW/GVuhZwIq8jZEXuLcprvA3TD4DnPu
wPURaiQDLIMEWdL6PCTNEK5CETekn2l+eyCmNirbj7NYfxFwI0nvnmt3DzX/2ClazNkZiwAbhWjW
TkOBFNmgNHpdgzpTYHMcEy/iUjLsJWmHYHW9UW/iHnF7IRD4CHgIFIndzfhzKyKHMQ8D4frfzhVH
RQ04wLJQUKjuHy0IaAI7FeVNUzvFlfB18LGVFZqqBHCp5XrxHnDj+FHnHW7Y2+Aet9cwAKdAsgJG
ySAiZzYk7h8WUStuklaKQoQSZfjvU/GSe8ytO6nzdP/oi2MdqF/USRZeGLGI8iYZv5lEUp32gML3
Y8gK7Qf7+TJV/kOsQBpgzbc+prB8WnyJLPsujID5qQocavSNb6Yh+WHOeXQiArgMeHfhg02oIkcC
Fg7QFhPJ6SdfXWa7kXza4KdN/2+O7zDMDx4K3sY+nzbPWbsnC3A0u0UQM18liP2jO1zXu53FsnZv
4RzTEFax1lMUnPaiBl0ozlWK57FDs5f0d+rD63z4jaSp4fgRIsSL80LMUqx+LcJg5oXzeVxKLMGl
X+vb/3D3VG3hm1I2X1MpwOxSBLOHxNTWpWKWP4wAVc1Ez38TWF8YP2Axa/7OtMOowoy21FSswp5K
t37O2r1HcEi9WwHKJ4LCigQzZgDtJzTrp2OLbvWLw6zeJZPOk1NVuJoBmODukW6GQ5lkQF+88YC9
tXatDuyIKQuVZP9cb7NUa5AvGQnjDHGrmHJlz/zYNQZp5WRbfu9BMh/8l5HhWwCE6AoZg6SGMe3g
CRHB6hG55II4eAYeKMH8BT0oPWRALHCCHUizBZNa72HF/GY220dOGZsoQiGlYc8gxZOkl+id/QrQ
fH6lwYhKFd2qiVfUegRQCHz7Cd8hSgBZp+41GflxZnJQTlwyojyHmRbtPEoAi4UaHH3qLUf61DDN
rBQ4dzYIe9u/9oJhL3crTJm0itcqWUA9QnaEUyrd/WH5mgpTX1O7moPH8Zdpzmgl1mmiTLUV42F4
gO7VnO5voQWCZVY1Zzw3N0jguNL+7RYpEzXc6ybuZ4Pf8l338Z48KpTSLdOAJ5zRmxPf8usYh0fM
eHiVU0yCocQEPqg3TUrWO3Dxy0TCj7RtHaxwoG6FMHq/y2D8oIU83YfAjCnashpAERhf7CLoYoCb
6Bk7P7l+15fQxevdbAir9+Dia8iwXWz1C+xHG6UtPbyb/2V2IE0eaThR9WhJ1UmChVwiKPaCpgRE
Ypy+xF0cPEk9S1PzyuqOUcF8uY7uBFofHxrDGpH+9TRPVluMV0GXHWeZMSfuHu6P18HK4+sSC3aC
azYOmFljpdMM0z5b0uLJ/xzqspGj/GShsEkOO9kQrbERTy/lp90lpxs1zGiTpsWqsLtQVJV6NiVy
DhbfJbXwOvZRn9VUTBbXUNCBvDYEidtKXyddJhSY29tKGMYGgc8sZN0ia42v7rp1DmY4Ujo4J0GA
1eDdbYMMMWv6/FMYTigkb16wFxLC/3hg97Yt7WGdeLp2YzEqcOcf7usD9NTV1ImcsX7p1kgyAuUS
RapIguxIbUBfaFdxBU2odnAKuHf5cj+x9MlvzvvwetDS7jGuKKCk9TadXRr9ZTV8P0hrinFOfLZU
lg1Eb3Bp/KQWctIvHtcSk30etgjszfmFdEuvnqNn7/GcZn02TrEKXW6BZ0oEKt/Wky0xYndnrYnr
HEp7xcZKipV1TIhOfUrF+S7HRL7DHa0ZZBulBESP42TEgQF6z3o5cjAYFQYDpY97EYAiC2rIWoIh
1615tbGe224eceHlspSTX8029I6JVYf1GmrsDUzbOy98jSlfTTGYL+5oad4Lwfu42nvK3zi8VZzp
cWz/Cp/LMezjHuh2gXZuCkdMlUwDna1iXeAw33hXyUj2upk/vi87fTtkVxXnepWAorAVDF73o+F+
F9YJ5aN1K/VzHws39vdDph/hNxOhY4xkNRGafMGhzG83cVvM1EtQhUill8ltLlbRQ3TsA+UVPOEH
Q4CE4azf3C7Ry0oCcL/2++Ju9ilyKYnpa02nB8GxCpXmRlArZVbAP2jNfzgalOkdZgaWgpibs2hM
mjtzcrzNEAI4T53UP7u6zPf5zHsLSfU2NTP3BUEEiCl9C4BKlxzuNh9I0szNKeMY+kJj+0OeJ1BB
PeSPR0H5+y5GNn+8IYkSctPY1/ZfSa6jsyJIEGb3ZIyxAOwJ2y2snHoWqWKrCSGSn57NTGzdlhzr
4dz6eqSG007HYLOXFr4sx2RPEyBB/wFpkmMuEb55sZMnWRwjcu9TGwX1brPDq1B9zcSc61c1mZhU
79CdQBRp08j8qNsvs9BsjvBbMVY2EMiSbTCuaMvsIBnZjGfP1RgWE2eWnQGrntwCW+IdV0Yt4ICX
cLvl7h7f22xyYkK7Q95m9uKb0coxFQpSWti4Dp2FeEJOet4qAOt6CZAsjXvlZhDsVDWugRk+0xV8
MDTi8eiQwAU6ycUfft0gg1aDyYXIWdh8vhj2H5MMrSFfzAMKB+VWt4Hc9K3+Z7qTQimbcV0Iv7+Z
VHBuB76oIuRN7ud7qiCzTWBx+mmCX2zAiXWprHf7fkuWjhhqsEsmjDmUVwt+Twl07fFoU+n1fe3R
E3qsUcn2K58q/0eyTaIfF5OlwDIO4S+wguULDtVE5JH2qE9F/vhWK55BKE/kUgxrl6zbv/ilB5Vr
rQsNyfqO2h/Gi2OwRJU7I55ADmT/hCxSoIQ4mS+w+ASpFyicp+Q7hpWCSqWpTLUbVmSVT7BrfUOU
KKgpa00SUZi0AKuM8ALYYtaNlfkuQBd/IKf+glbbVhGqJLS1q/beriaOK9iTvxuVWjXCJNguNdbY
Nr+0arEj7ICH0W0j5tsA00i1lY8+MXSHVaTKi2qBVIn6vpjXo72fAhd0M9FOaaN9RCiz7QkmbmoY
P1tP79gzpBVYCM+L5MV02sWs48z9GhVmqD27/dNvtBsNx7AL7zhSEEO9Td00MEQe4n8cB3+jz7Mb
hchqWlEJivPjbeOm3H/9ICee6bOWgCbhBiO/sV1OVx6nW4J+bZhCWKzKKSSzCpYai4p65CuoLrfX
+qY7CLeb7fO0lffyEZwqFC9hpzeJ+Fc5LdcLO1coJNrGO3u6CDEZ0rMyI9HJlZlFkuR35DTCHd6V
60CtHkzpBTQ2qccmAsalgAaX7YMKnPHwe8Xu0nfV7z5OmO0m1g0GjCnf24OHjqDwzeIJmwrJ/mbC
j60AGKkTSu0GqrLq/MdQLq4BKgzuI4SznQKGAbTyqiw/tLgPg8LVt+hpdJ0W5aABsJA5VSGOHfzp
m2WxDiSZdRm5WU3/F0N5Qu4URYE6bjEGTX6XSLWbAml1uRNTPtPkvszWrcGMYFLsxNhM/Mpf89jg
/FCPiWZvp4FSe3pslOvr3ySLit1mwHXhggu0SthvZMwNJziG/6oAIEENZdIhoMMACZ6ype9F8Kky
NH9HO/rTqtKYLqCVxIy3xepTXxmwAw2c3Ifpr8aLgU4CnPEm8Gjhw5z8WSU07sbyfjxq4gpoUT/e
AeKykwql4gtLK5EilzPcJv2bj59Tvzr6IUtqxQcap46LN7e9+bQqoayRjqWvnd11e81fZVxrDaG/
szPmUy+ukk83rq/CF9tgnB+XME1ro8/LBkCkp80sgM1RZ7ISCDzIGsv3RDeiWtkSK3YbQoLQgosi
yniwKCmVbU0nu6+HJ0dzu0h6VgXBaMV0OhSIcLldcb0Sb8P6TqYkb7fuS0RENtVIogV7m+Acg9JA
ZjBztpF33xG8F1GMLmvarQgOtMz01WxijWPQNLN3PrLzxF5Fq06v3pYwUsgKvIdbGr1zqmIugSpQ
7D4xmoT+hKphYSxSZTnAUw2W1KJy9zW0JDTvnVKet6Dk5nC03MtttiVdH+4zM0aIAAuiXEfCKFBh
DLVxjjh+OPKcHHKm1M1CIzGFamuJM7tMTbTiKrpzhnPmcoztT2c0R9gBvWr5cAw7brgusPiSBLtU
zUerg9ySmfR7A3suO8XAlWXcdBtX1ogRhOd6qOZMzGgEpJusbmgq6eAY+T2lB2z8UOPCvzwCz8jC
1fGiuxhNTMk1CHOJnNeTpydB7HWvhsbrVu20iEY0p8GhbYxMxmq1TLigPnIxLZMGGidAvLEuoRmO
0k1fzPtc4a7h0kV0gBgG0NMhnHeAxtOBURLIjKK/3momCdmh2eLA1NKomIeaiCVum1rXmkGRLSvj
VpbVlwAJrQ/PkLbZsFPznyAPQOT8DLIAT1IdVzbVQzI7LYcbqcIqavgfPh4xm9T7JZ2YxqPmILu9
iZwL1vAsnWnDd/ZPbvaiXTDrcnZCTbyCEbPTj3FGWjZFV/LOpCl8n5s2tFT7ZUcdgKMDxb3fQsvG
nauhJUkhrx3ApEvxBCzG0+/eFAYdQyDUJ3uJDwjgPwQjWvND3mi+t245y6ummKr0DBWnYT6l2xp6
hQ/tV9t5BaTaPC5fvI5CxtudDt2Z8pycN4SuhNVAFW3G6wSlYtEi5xat8P9Tvo4I+4jTyzHzMOfQ
7a83wa5g+g1cHk0h+wVZUWYN1huW+gDHrj46NpE7c7Oxz+5I/Gt++EAwa/ckWpT7Qm2VT3TjF18a
/qgpS3tcNTMarcX/elRl+hfma2KoSsfypZ/6c/8xQ5mF0iYl2pRLXPdjh/bUmFPyIetHHWAK9fKA
EnMiXu/jHdH+Nwnq2BBy62uMMxkqf85p3u7N9Yg6Bg9E9vZCg+q0QgJxJpuvtHhi4gpCqni74RuM
/FrvmM3pi2LipPe7y0U/0s/Gk5IkuQP5oCX90O/Sua4EU4MK6adFmaENQ7uVRrRNgjamR9nvdlRR
jXi3sYMqS8TXj2DOnEiH62EL8MhrxEsVGqeWETKOyP/1aTzjwMxrt4GEdQ/YJgXNo89xPxu3OjgL
e0Zmc73zAPF/zivm97YQgvZf/ZCUGS3FgmTJOkMAcPADxy4XKycTPTLM2mdWkK/QDNeuZ0QQo6Vg
QXcX7iZJilzyAL1rfL3uxENS57fNs1pSZUuIU65bFwaJcaM15YgyIfnF40Ckt8DjTT4XzlR5f092
l9HxYHe0X+EfKaQGHobctLXiXVtOKe3uZF3qF1Qb0RSQ+d4TpYE0u3ymePX9ZAg3x/NRAdSbZK1H
SuiNcz1aKlDFizX2G6B30lfml5hL5vLg1IKql9va11Q4o07kWHL3/7WXU4Rgv+HyIrcJi+20cGe7
CfR0Dl01NEu0hZI9eYaJaj8rGvjKU6+QTjegRe0Lkc1CZLalrurNnKSTboHnwADdI2HKwffW9s2z
ciBXQwMwWq2ifTnWndV7VBqz/KyLBuxUX6ntb0Ou0LoNktkjvAtg1wjQHHpp8+SCm6aphtS8o9Rk
ASnVfiLq9HgRGPiJLGw8h9BeXmtn4ZP4PCTe2WqHeBdZfpQu+e4B2k68axGUbHcbXLTbQUhLZe6N
YpefBegkeDV/A/FX6Z3rZ3iSATQ7EUGZc6jL7uUgPvc1/TSithcqOx2iR6adiCn7zaTbiNA+SYAh
B57o0DuoNul7WtdKw0kdp3ykajlakXcaR8AU8kMRlXUENoCnB+3U2Op8RaOXbudQUrixOzDqH7bk
G0JqP3pBdr1DQT+uvJQ5zZRk5Nh1L1vL7uSWOC+9HV2/K+ODEZJeVC5Y1nT6bljpLAk0IGobti3f
uA6IoRINBVJu3n3CtHMhXwVbqsa80yDyir7olThbeQ2vl9VpW9NLcN2rgHeWJU5OkmXvhz94khrZ
FbNrJOf1tHRRA2sIVeFHdK8L26FhTH7+A37iJsQmE5km76fJcLzggpRz0cICSEbSZY8oyGpuExBS
jmX/p2ALLX2yBhxtkh+Yj1dRWiQo9lv51DjtNTWutcB+SqZ2TJT+9zXrSXPZSohx16EMGdDrOhyN
5tJld0CgSTIKI32emgAn1XrpJrAIv19CPRvYzURiL58RnElaOFJIiPRPW0LcWqiOd/JsvvKUxew5
RMac3M3aLoikcCtzHsPKqd64TLQVV5ecIX125ihWDOjHrm1nrg1QbTsqn++kJb5NC2BaHtct3O1u
RS6wXnsbLuCBpWvblsvDvaj0bnPShLgEBsBfKFiIjnWdwF+DySAPIl1/+eoqddGDcaPOTgN3EqqX
egT3//y45fqBX082BmHHvQn0eiu6oxx/nEbQvYwdC21piSFJtgeT/Ddpv2AoPW1xWxcCelTTsSnB
6MxpmVnaK1bXmLPIMZw8Qn+OaGcSLW1Jw49xGPWR14uje5D3AB6MG+5vnVkivenaWdoiJ8Byak/8
+34HqIAtJB2zma9JRlPDLTyv6sn9pCR3sVn2XO8tFOXRtm6rPZ8BlEccybQDloLK3LUJDOLlxSsk
X/Ial6LEMHi5drTOTdybcMZZ6k5+nvlyrtsD/QITUOraV00g4XaLu5uNBw4A51cofC2ly6znYvTX
Og5iov3TbWsK2B0TikCZPtDcTSkFws3GcClD1mPG+3qdwnvOkTCiC11MZyrdkqZXDVIdnx/vMwba
hucoR+XY9WAgpRcHBaw1hYBjPpiq+DeYhlEsVnflHU3rcqothmShkYU5FWd6zHhXjhzY5lVIkXjl
w5HPvMljQl3k+czgaWQzlMJIyde39R8YE86HejsuoKvX1jbbgeKbokgEEZDclgYJrYU28LfgSUBw
L4M0AkRbG/Ya22BuS92WfmwredWkUC3asvtVBDzoQOlRY3ESjqD1Logomxz6CqHKmAErqYKYxnW6
3bqoJTgH5buELiT2+u2+s2uLdyTy0D7kyUDLC7a3ugzidK4aZ/sVyUBqUPviLCduBgTsaym1rHBn
LuukceBmDiESBd3EDsf1R+apv4jPCXPAkZmoiiXl1N52mtQGn8dQ63ahdsIdz+BhHSeWqpPsckjb
v8i26DY50SO9TEiyFwSrvacWx7ulvVMDPafs6aEVbGtCPHmFyT208eSoNtArzJaN7UStHsMakfDJ
BxICmUqE3RRHqvdZSBlxDD2jChHMCEItVEvnux/GTVAZhCPQS+mj4RbQ2IzGbK3j7i7a4k06xiFr
COBTQ6Y/wKK7aldnhHFizlyQgkuuUfTz/5a76eZw49ncYQ04htkM+gp9s8lHi+uIFEdVttMUCscj
gw1+0eribsPKGddEN7//euqVAUy3/nTH68S6Qpsozo2c6mIKQWsrIDzalB21j4VWzFoHUiySr11k
Pz8F1OphWvzJrFtQCUX6VclkVu0WBHJ8XeZRVjfpQjrD2JvyvM+vUz3wdfq2eqrP/xs5U3fSq4yQ
pt48vNh4y0ue0WBSxkzPuY+M62nA5CxG5cB9jPyhVKE6N587ZFUffpA3OjbU1Fri/S6fJL4dB25g
Sd9MvKUknjhUUzCbTnb+Jl0HfesKtS2zw4GPK/eYC4hhymXXvvhfpATeq/JEGZc9+itxUvi2Sb2Q
10Zh7IZIFvMPcoHFco9KXkT6rN5u3/kq9hEAbo9w5eV/7s+0BNsrdy5hzKvgB1M/SWauoZZzIhIj
ppMG2QOHx2kleBRTM33BDLMLLv/MW6G4l1YVZgJdQXmci+/INJBmQLW7LiRTM03t0DkznQCv+WRU
z1WBR87wjCuc6xNdoMNa8qGobcdr/m3sWXiierwqslApSmT6pwZUiTZEErJsMIIxGoy/HFOgy/nB
W4lKkKSOwHY6C49cqJu3r74h8BNc1KYKjMtqrhoWLA/E2IvxAdTTT2hsB77dX/I/egJnM+wHnr4v
RaGgTwLL5Vz6pPz6fH/sh6wSs04VSPKsa+iiKV2iGnNFcDODBSx/+KPMVVKuFDsx0sURWk7BV9xK
9K3JIFtkLPQ85TDxhAqSnft4cbBmalyoZhZ0+pPOJA+mCERixBDY5CWnHpOp0hlELKDwNAx34+rR
GB9af9QvALHk94oDnoJ+bgpHWd9P6aH3+9mlZDtpytKy+pQ4x33rUNCY6FDKINLF5nNF7pvQXvsb
4eL7/W4CCBxsV6MzzaqYyNDSdNVZwH/GHaJW1BG1l0bRNAPddGBjwGAfl36BCLvaVsbc1163F/10
Iv5GCh6l/y5HWFsrijHAMdBfnYMQUxYXl/fKqEUPYxS1ZDegQpZIiMcRZvEYAYNUWUCVicDOV4eZ
6uiw2TuKdrUrwIZCv2zA13BSQ42hcmpR5DK8zlgYI6H/6h5auFctvoXBN1Chrbxv44jvhTvpRhz7
enzIO4ilJl/RH1xdxd7R/rhV+7UvDBUCsrWfJwB5Xy++OCvnxOtuJChH4CAo3R1VjArj+s0C7eDH
AHnEIn5LifFkAy+7JVOspwYmD5fCrDgBWhGgDP9JmXc4jnw9XF3NU0YOC+DE5EYN3IkeBFkqTq35
su9sL3ytlsAu8djACXtSI9XWnwfnt6fZU9cU0ZoY88nKxzGGqECG0nfTqgxPyDyx5rU3vc13sxlw
vAznCqi+CIVxGS6+hjn4By4O/QvdehHX6oL8NbgbB30jiZGNT8snKpDQ9sA7UIZCXHu3w88mtLGO
wQ87s5KgS/ci69SCFPPRi37hpKelX4/rmSzjJGkFP7hEkhJPPEmXG0ZEitIwuTpCRK8chh8qdDKa
nzkb/6OwrgO8NNKQ1eS6WPpD5GFH7uOmzLq2OQnKjhOE7/0UK5T4wWIvGYWHI46BwRoU+DIOBDWn
NpzyfuATPW3ifRxSULLos7eJuFZlt5ilBDXqpApQFCUZQ+8m94uLiONPdVZyGZNUMpE2JiV6NWlK
cjMvdEpxu8lYs6EkQQX8w32Y4XEEEcXEn8uk5BYMdroOfR2SmFuMNXxiS1SaVFgw6qbho1P9hOTs
4FKbqgDot2XLOQw1yTtJtSYQrozKhKs9BahOOUtTd1OsGG0EQnlajUxBLLhNWtQlkaw3cgN/TBaN
Vcf2tOExguhRyVlAgUqttF5HJXVhmo0LKCogK8SvjZ6FohagqqaCayDlfPw5AcJl6ey6M0SWkPzi
fKrg8aI5B3XeOLoTAJyZjbW0J5Ccll4CHMx4ksBNYj+CvKHeqFgmgDWWo2OK5ydi03rkdge/bj8X
PkqTz0IE8yjo9W1LXA8ZLq9B5Y3rghPNgBV7kM4nqcX9khFxWPA/ZXf/F2zzzsp0xhT+M9tc6FmY
RiTc0DnM9fVij8Ji8IgCfhOsz8F6lyC39tgPDrNibSNA3BX4EJZaqxohfWap7s3bmizOBiImyaHc
zMuz5D+dhiSrSNAdDhX0SJ5ZBBQr1u4AxVjeBkRpCpOXYdK4Lu0LyL69zg0l/cAof7KhK5XBDfOp
zATCfUPmJnMeRkKrZRyggh+gEty4zEIOiDzA19sfQuZJPGaverfARms2EGnJ+uV5Aqtj2QL9xM9D
QPh8GdumXL1Hxn35RSvtgm6MM11g8csAHhCpBc1MpWh3BNfBSVpDURMiZeH9FvIeGZ+xXFHGbwfG
7ygWYdpW1WCJ9tQMfMbgL1gQBFItK8xTDas4JpcIBMlqpJ8CZLwnxUKEJrRwffM9B6LI5XvDBN5T
KnyLYW+V092VrC81Q0n2vIPQPY5taszON/B+NNioE0jyvorTLFhNat5X2+J0y0ozR9bssamC2U+O
BsB5/4NTRbUKWEXvLf58GcNJcqESSHegxd8VtSiLb/qTcqPzPw/LHzfXSuXak3MtY0d4KNq+nyjX
Y44KgQf+hAbdfylc8ptg6juJ6Fcuey7nVj3LAhpMMyqzoOBm933u4SOM5a6jYGOVwy/VFII5ApkT
Ljl7P5EzdjlQ+KNp7K6oRug6yR9VAQ75LGN8BXiUeoT3E4UF5Y2BWpEjTKlngFhZfqom1/uReBnO
Agv7atVumLMk2DD6qsGvLDBDXz2IgumbvHFHq5EU7L1bsvHSe2LvWpth/gIfysMtIyt727ZB+rBR
G0aj05lD2z2S9NvXTVQjmADd08J6GpYu2tU9ZyYAptAVuz4XUEl76Bs3+PI9O+Cx1cU+cS8Kv881
wgSBLwanYriaNXJbNHw4hj8h+yc2CVMxKVMmflPixF5W8wJFCy7sCtYz2TiD/Nm6+AtqDhYVAGpW
un684ih3OKcgBjn9DrtrwmdZWkdS7ERPYGZDdQBkPVB5BGh3s1umrU/g8sa4URQMzafvcoDarDQk
cUfdDiKGG8Q5VhRTXx6ZNtrXXA0oat8qJcpmag5aVxE3aK+7F2zWdespowc8YxBgoc5S6XpfLejA
v8PsGGEUr9hhhobrmpn/bNE4N1EkqP37FuW/lyEwYVt+ZUQE2wCIayINXx22smQAvdfvFdy0/PMb
sEI/YtCA1NfriJpdVNFnqcqOZP+AIVEjlQl/Ma+imGy43wHGO6csiRGGEGZ2OUfuqX4s2dJVxuL9
7fakx6GZl+3Ep10lck0+9NdDLz7wXJs30n1WdpJE5cVLIseNJoah4EyjrRKQBCQDTFgHGiLDsy/k
nu6+LJAQmlgeWNxHARAQ/P63lghmHj7doW0dOesXh0Z6UBKb5A2nawKpC8MlocZdfwimeouZ0fJB
A7YiR87m4lhQwMb+KxuoGwLJvPogsN7kQpDqRatq+kCXcqP97BZy4kV0UgDDt+Wm6IYF2uLSooJ8
pQe66J5+UBvnbg983Jho5vO5sut+3QM221aYxL0DDcfREX+Eb/pPdOQhhtBcPVxS+RgapjHujdBw
VeCIv9ZrQVSmh1aF6A73X6bia0VtluF9yeYX/Hxdgf+Eo+J837+aAKxADbFBtB3OIa1+iN7UHJK6
TXj7bxv95F+OMq/aZiPN1ONuvmRk5NjwbPq84DXqgoUzhGGnUFE/TYE8LUfBlsBoXkMRhHKnTUOS
G4Yal4ao40u0YZoDri+kGFuderaXQFma/ArnqMApZz91pjk+G++YQoCvgNz6B3O2+vzQPmzb8FtZ
OZ9e3hnHaWd0ZxFQOWqIEk+QGxTF0tq44fCyEEzAWbHjGTVUcn9dNOvk7WKBBmsln+BEWFueqtfS
JdUQb9oYQW4/TRdE7QE+hPplwMJG8uXz0ADN0YcU2KQ4Qj3cjIOmuMaPWHm9Txz/CeIjkV247on7
uPgx3/CqYzdMUWm0DX2VUReIWIg3vq5sFBzUPq9xS8pg9+VRyGo/rU1QEcr3I/T5yQCrjterQEie
CAafjok8yp7rPwoxwJg0GXX6qen0DLah45sfKEhbpqU21gHY459Z1ozQGuTAC5RtTMZ5nDDZ/QpG
u1q5oS7wBuaxhgp6ytUgrGe7DTF+9s38PL4sV9R8JaCUIXJNdc70230gs0Sk6RMSTNGVqfjza6pk
GZQwHV6HDgLZZuj6Beic3wBlSIyJtp4xeU7DophrISGrIf/+1zo3ceO//8XdtMrSfkH7ent0z74D
ApzGreVzikSdQpUq1Q3+HIZKZskvGxGK9/z37iu2Pg71DjyHtRO+VpT4RxthQReGTqmNuXQej7lV
Eo/F21nWbHtZ9V47ZgiPKQ0vlcvhXWC4MU+IxgJvK7TLlSemtCSP2QAKiGBl896YSVCbEXXBKItq
sKOYDJ8GmRUMT8f65nj/XTXSebshKMDIw4WNsjsDqtj8kpZed5z9uXQDXzZJpZKzyk9IJvMaf5Od
C6WpZ8tWavwxIfUUHJVOQRGbjCSUOzD924WpB0+H9znoikUaQrw8wOFy+XpLomnwily2sDd43Ef4
jTQPa3SIS9kfYBqMY2j3WXtaYABhS2Jo4L2gYTqN8F27mUmLkTmP5QlSC2WnYgu1QE5FgxP8Qndf
GWpZqhTYvuiwVFLXMgzmJre07III0LFhQkPSh+QqYo7FYexTX1DGI+v637HIgxs9+CqEcrlIXPpq
W0jkI3MXmHEtVOiDkigtH7Lkvbc7O/fc6jRKcUxrtqVe7G6Ao2LfMvBog3Zo2qi7YVWzpdEGudsr
CVrSBXh2gwhpma9b+Bbd9sScRbhKy/Mhfba/NS9ruaj4xvThQzTr449fbylLiwJ3/A9kA1aE8nY7
XWt8NQ977mlX1RpnSLpftJFumgmz7ZT3FUKa+DlyOEXO0Q/Q/dHBUlZlTSG+ijLyX1d7Du26pV9N
tEmjP8CqYBEoPE5cziE9smlSVz8wct7+4BiZU1R0NSB85QT0nthUUhH+MNQzVPihdy3oWg+YRAcc
Z38WHFnsEz5LalkE10+hgHEp7pJa1a/5XSccPyFA5zprT+z/cH/9OZRG6W0urxHnDBsJvRp9Mzkf
fUoFRE4t/n19wzG/0SlXKxYYujLRj0YTiyi9qwjRGQArkqGGsRA8o5J8SUCwPdaN4ATlQ9WyBKtX
Qa61Yj2iSjciF3B59PieqZslqmQo43AJnoycJwUSu3u42OD875/p/2a3jcApbyRSTF/zoL3IGypF
HraF7fsiZxlBuQtYYUe9l9Ynv09nL/gEQq+hutuQ1zJchQEcAZeJC2kDioTIhwtc31+1gguU0gqQ
XHAQokxsKxOkItejAVVe6u74HTnCpRXeL7z2wMGStV4WJJ2yBYuxQjrLG9vzHN2yBvsxcoe48nAj
Zt373u99coN1J1M6u/Ko8xhY7WkH8Q7r5G2wm0NqFPwUt5bL3bCM9n5U3j9J0uewOKC6PfOfSlUJ
4zjt4DCUHQNSWhx9JISYFNEniHgF6JgGTNEeOHySK66RPoMqFiw7s1LtSgiPQAORnEpq9ibDRj9D
EF8iHrRuU00OhBjeWrI6bLC4FFq+7Hy779v+EXwVFQqvvLE7Xxrubu+4ZsAr7C3J22RjLSOss3sv
Rh94Lk1Zj8/LO3xjXG9HrsAN7tItBRkysLZcdzszzJCo0otC5bHaqCcW85qPaRc9W1r/8QFcRf8B
qEmEzo6syzyGBfqK7rZAxB5/qyG7P6YXqOrDI7XhfKo+2BXefqvBRZ16/a4GFfnghZgMaX0ChzvS
9jGOkKnFsX6R+c/WM2G9k/5ryHMLN9adld9dImBbxXkLPJQ8uT/keLWhr0s2MUktFoDN5DXYst8X
9VJRyGPSstYCbJt7b3T9ylNJGAvb6UDRLF4IhaLpi9GkZY4vo6KyQeDcedEyPPxbhuATnRkFlLEE
W+PI4K51eRjPdvqA+lIAd/oMFo6FcdTzfT/ITsWiHUil0kshJVQyd0HZqXNggDx/MLIa3BEcokmh
qb0y+BFJSwan/8/xr9Z3dUiazIZOm+mB1g7Jo7Ay32yTWeM/1ciQ/wbSQHztqACff55NSxXkqoNp
0fQdqHC9f+Rl0BMEImDpfK9l7ehIm7R7sZ/GFtcq3rEwRze4y9pEkXSAI6xEaoCmXpLaiVWOXkWS
lYpw6GVaiXWAePh6PIYMUtWyWFS/EiWb+r1ey0m3bnVHLR21JbNa3g6EdgZa8BKvoWpZe1hG9LT2
bWN3gEPbMHh13sfG/oxH//oJGSwDeFEmeav6bWZj8X9T++hPCFvow2M2Far8C5hBoYJgL0KeJTM1
B7TZ57bxs58zfiGlvhC3OW67G0agl+GYghw0HOkQDsHGeLFHUQAtKj3NP1WsadObUO/shtYrQN3V
y2QYS+PS19FXbpBMHuF9pRxHuFkYS3PQmXmEgF+LadYTKKuMvgH0Sr9lfrE9irVH75U4slf20PpP
yydlHqhbBJljsrFHc+nyYGTR036EwYsjyFi17UUaSEnXGa4rP0XXo0SFn5qy0AlDAPwicHywci1T
mZUJ9B1LVGRiBtD0Zv7cuTMn+GtCMmqPXDV4M4zOsWdm4785L1STCpQ8e8BmAcqV+zX1mVReU18J
247do2NnM6pq/vCMYUQTu5pYtOQV/TqMbQVw+ZX1DaBsXOT/chmWyl75k2VkLlCbtvhavXtF0fbl
c0ri3QVrSVsLUix3y/8u3pzE1D6YmbaplaiJIeoCP68b56VRpSuk/S7OKCdMr48m2/XkLOJEFlgf
wYJqC37vC2g2DYmY8HU8OxTHows3OBjYnCGsXuEbS8W3LYwlPxx4sYSnR/pdo3pJAkVpoC3y97mm
TCf5TK+g8kuAI3l1BxTzY909/FmVXzdOCQB5HxVSUJ5sr8oD4j96yzw7Me5il+avPTtR+b4AnSBB
GnIrbIVq5ob9jClSyS6gWaIGsFgWQW4BCRQmlHLe0rH8cX75zYCpvcNI0nKiFIDXHkmP/aU7G+h9
qe1k1EEGN6ZTDOzuv3WQG4kgN4V9B6hREMhoU9ohasyG+r3a5538J6W7iahTNOZessB56VZCa6nn
m8PDSq4yz4RTAcjkAgSPiAhIiucLC+nUDWnb4CLGTfD4iLX+HAPh7JwxiceBWGyNQbhIjxKU/xyQ
btxzRZYn17WKJXOayfB9T+4GfMmwxnmymgxnGZ8AjijlHiNDrf8tkIWiFpLe356Z4whC1EEsMXp4
BtGVWpcx2riR/5KX4xNeQHBEicad3GwCU24wyZa08YjSgwkAi6L8UNxYQY5cr6D2NX/88W53pSIf
UMjvQ87HCsmJkniqp4894A2bD1WaaGI37chmr0WoU0RWYL4iW42xvqYmf4Xr1SYQiRXRcNEIPwBZ
i/5DeYBmj+2Rk68LCiVCjoEp+RnsSemRT+nMR2Qmc6Tc7kJ83C+Pl+s4dfIIJ6og91kPa1HfJ1hm
OM5tSb51aul471jqH58aP46P2dA4J8ckZdc30J+buUHaLPb3a5qstBowMxoatzh7lvHNYliuF7jl
qLK5xq+3IcO1dnP3a8Nv5+PYaExiIu4yp5PrZ0eXS7EuqkWKYRFppSO6gbUHpebSuYqrS847VoAn
Nx4f2Rbve5OdRd2r3A+wD9cIfVKw9n88c9FElH/Z5eOjk7lRmJS3sjeOLEchxhobqWkxuJY3niyS
CRhmORMEHZuGWPc1IY2QcIGZy5sttgdLKwc5cY0vOjO8xnlSOJYasrxXRSyPjGVk2kzgd+bCwV4e
2tTpG22w3LhyODDQrLNn8E88ySzdY+LK3+J1J4mGL/c1wz9SLeUf2dG22+4iGDHClv6WgE+n0jn4
SZJEZHmGNNzRVhXg5kWmkkwjSma78TpAdJba6milldm+QSTQ9RrYpA0CajjvwqH6jG0rrckHYNqI
dORx0uyV/U2o3B+RwNbfRBHZxChk/VwGirieMotpKdu86VS6S9iKlaKXBIGvxEPEMvGNhq0mK+yN
hOZNDD/4oJW9rQ8crFzHt6KaM08CXu94fqFycv3iYwEytUp7C4I2/Uwbo/CWO4JHkl/E5KbSXqQR
c1/f/7y2BP8OYMZy2ZDcCCgGiVtMs+65vBJoPPiZ5vLJ5ayXwpeJTcmg3ZM19g45MM0oOnLgfqK1
s5plX7rH1JMv4/eAmTB2DBtRLBK/fwPs6bGWOHu+AxCAjm5yExHtU3VQaMGRtTcd3W5fINa+D9p3
nMTW8tkdvJE/4ZuIo/s68a77nSOFkiNXqed38AGbwmuTf/plOawUVTLcLniO6EkK5cNWiK2xNkUw
V4LlTfj+e7jsheOKss7Ws5g2ugH5UT5Gj6oSOBm5VH39HvgpBJq8eSLzOovCfUL/ldTPzBM3rhge
EprDLMpQHrXZ4PzPJl9vnmUESFlBedmwGrYn0RCcVV1f1bTub7OQ3Kw5bF979skTTo9hIRBypFyI
xkBGrVeNdHEH8dvQIxP2k72jBwnhjPU/Gd79xjNEUQaaThIJD6EcQY23s9MvCe/dpvSlvT5MPNW4
Jkq3v1Kv+0Y/u+Et5J8NrM8b2Ppk+FXHCJC6RbwkRnc37mu2xYOTsKSro3G7a7LKijlir3Ql4bnp
cweDGQtdCgunQqFwzb79QPfm/pq42PsLT+64MGmAI/8PcdWdSNrt1Y40xy/q50dWOH8R/IM9TjwT
J3K4sB8fs+w5NChaefiWW4WQYmM+jLgmOdLvzKLotHW7HMk+yyVVYSsp3qULnpwR+cGseH2NQbE4
bkdfG6pr3grqAzHS4Nxka0z3dWmsDXKTyiLturRZ9c2i5XSnQrWjcb3Rb668Ikiq0WPeY41sG47r
oc76Tl+cJDj4yIu8VYgmnbvc1JJ9CBhIEv42IgABvRKXHrI0cKMirKL9joCBriddUZGxyTUHIgud
/n+7jVRMTlDDIZQWbH5269ZwwR0bcBWwtjLEqvNuNTYjo+Tz2OtoN3iEyGP5Z54/uXTJxz1tXxv2
4S2YTd3LLvPzdj99LSLF6kNopbzXct+Sjd07ja0QpSTrUK6kZEtpE4SoVkGKj8DXnWs1ikFNDmEe
DsJngMITID63wSHUdeg7HhybZlmLwO9ELuCI2aNe0t/3uBqnun/u12j58tqQpCNz8B2J1ap67xyz
5TuF1NyXgFv/dgkxKZrTTJRldMSGHY/6GPutA1RL5GqLtyObymDkmQq7Nr3RrxFEPsJF32Pbi+6d
Vl5ZYuEn3AD/D3rCzhYEAiWUV9aQ5v8rkAYHInWdHNhguRFdke4kfVE7GuNhjAPDexktchRa0lEL
K5uIT0PE0ZMa6NqRLIAUWn6dfNYBpeLc2CGQs8y0B4X3Fx1k0d6GiydwhRFwcfmxmbZUal8jk91c
jLba1ZSqN60sssjfciBXnsikzq6UWf/f8Us/Nd/IN65qgravzg6322kVix1MEEWmsNuAW9XeeIyn
HXLu5Y47wmFQ0jdHipBbRO7QuLOWIRDawf2MdNEG14+EHPZRRa7eFiNSvQVbOuXVvaAehtO3Yyfk
QlNJ62VlWOOD1cbNJQV6Ba95Yog/4gUozv/81FtsZYDyUCw8X9Gw5H+oyC4HJV3M+dryfzhTu8yl
IzlkoBG0Q4eGk4Pl2h/9N1KlmRY/VUIyHaKl5ehCF3Pi2iWiy8NXsN+tsmak5pnv2jHurNm4y/Jv
fN93iFsNFj2X6pLXEhLVbnm/n8xx33YrhEGFYfeqTFvf+C5mikaOtQj7A0jlTFlJ94DgM4A2mSfw
cmViWJswOv9VQLrIU81p/2nb6BCayhD1TqxeXehpzvIHbdUw49oCe7lzxHnBcKxKhs8oBv69NJBH
QE87cUourbwHnzaM4fZzozRHn+s5mGRruxOi7yEvJ+Jq0meodeQ0D5IkuvpyoBKeKaUKsQ49ZhQu
b9RwIeA+iyuJLYPhPiSC+ppw+O08mXBrnccl0q+udQBxVRVnJVYpbNjH9tAkZP6Arg11M++vT4kY
cfZa003PT6VSHpRqCn1AsfkL04t4jr0xi/IOLws1RSVQxJNT5lrb/6DAoxyI3W1kQULIshPI3HIJ
H0x9PghF+TktD+/zG5coLR9wNZ9gB0ncoULL3qMqhG4R4fIuXWTGD7iRmp/m3g3Tob4zoAVuUs3g
HAOMh4AB2zCK8Kfo1kO9N2WgLh5+aUU+vnuR+RVnudGBOvMD/YLcDio639/A5RUzmxtSBbJjL5wv
53DUeK1xbGR/+Sh5TxXRs+DHHADq74zjGqnhm46Jx2RErsn26RAyL636/Ri3KwBJrHbHbAszYZIR
w7UL6rACNk0a9w4bDROjokiO/esW8yPg9Zsb690uPHKZf9gtoTVILs+v3hyUBPMpiw3H066SyTrt
yMOWPM2Ko2TLu08s+yIK2RmKap62R+tfYujpprj7jQfbXbLnpjNgnEuxWXNaAFzhD0mYBRJiMggV
biwOlW/TJaa4QDFe0RkC3y8+ChzbW8+HCdvb/16mYV77ZoElnM210vAg6IQOynJ1zSBi3shMt3bk
o9S6IYcDAoa8tdt9au+Ubdq3geCQbKoBTnWu9rzt6PIEP4HRtEa5qjIhr7IWIGufCMWfxT+9mVcf
vs7Z2NgkI5C17aQEvnr5+t+Xzc4cNDb6VxPuwJJkYK6HHLt9FpitflJbwAewaTzkyayPK7z6FXVZ
9U1roICgRAGuiV0jzeascHaAAmEfdGDc/07nCi00wTaeXcazTK/5fzV3AIVi1He/gamlhHr68wgj
vzTxMaF0ZcpARaLLgbifRfmgQJzwD0+PxpyemEsYKVipDnw2KYvMs5z/SRydhr+W8abRPOAcfFG/
SZ5U/xsQbypg8Btufud+P/gyzPWr/NOd6Tss/MNyzOGpJaRoo3WeCaLNKV5e777AEZTkaXzmUUwr
iz5lJKiDhV6HwrZH4u1AL+Y+0RNO82drGZp4qAnwsA/vLNXDnNfEVP7sja1OT2uHGfTi+ErPJDIq
Fl07W7lTDk/tzOWMv9Oa+NXtOdCtyhL+D0F6KA+4x8djxwJ21IsfYyQzur04hvlJ7zSPIus6t92r
EC/LhSqEfFblAB53W7E17MC3yGeG4KNJdkBaTpIfFFy5qwCPAaCk9Yfj3s75IPVaFO4xNL+vCQA2
EaLofMDzNckv1VTlkF6KZqWZFW2tgauCiBwO6kDZSrKa4MUT2KfV1aBLcrh6SUJcOiw2rWR/wONt
KraUFT04edEhYPjSrI4a+GKgWTlYpy5HdMcalAPrY4UG5ItazuPlLCeamgjiZyRp6uzHYG1lBaiz
H4k6q5I18IriHYTauL4AHJ2M/2q0V78vIISMFSpBko9Ty0+M0mBiuEuk1/MHrrSkEuuCVV3PNHNW
z81QW13RvD4iSsyqGrT1+pWDb/IRcuuv9rBr0y4PkI29oZ/37WECV4Qjgh/j8W68+GVFGJDGpX5h
Z03BYL0He+QkoKeJooEXtQ2QxDB4IR45L7J1Ao+Wp4/UwHoJvyn6QhtcFzDA/Olx93m4fxtOtBbP
q2ije0LSyd6HiP4KxMzhAIzi8al9d+fwJS3OwW+JWP6+sHlh8Yf6AmGKQokyuxgdRGNgFYgJs4Nn
6IaGslr63GTeWIii3poBH+dz3x+IJU02xE+nPJ93hSe1CnAYhO9xJ7vweSYtbGFvJz6ndFlN+q5p
VuGqTVfLLJcQ4TApKctRsxcWq4HgLT3pLx39dizchZ2g4tWP/tdui4dcT35obp7lyYPfV7QzGaT8
Dp2tS8PweCeohuDrhoT9S7twC9zCuZvSM5pNx27EL0aFyzWu8KF22rZH6DO4LDEmhchSDIpzoIVJ
sFCLBuztj3YhuKz7Q9P60dVOmbJnVm4AboQzoziIiojXcempNZ4evzccF2fISMLnKGsHacNqcPnf
o/hyENWDB+FvxOLWYIti1dQXA8TGXwv6DAm8DrdMv+qZkqVLU+E6sMLEYeQ6qEpbdxiJfwMHAaEG
1rXdhNhkPbKnJYrY+kTEci1b5Fa69ixTx4mMIL8aRpTOG5POHYKKLnDyNI9FXWFTH+kXjub9iEu8
7pDLdx+3kZXCW7ICNUPGIBtbGyRb75zXALbXDjLh7xcNy4z1GqRApMX5XjHFvC015cEUGcPgZi/H
zrsAst1xmrhwS+t4eHX/mSK193mqi7veCGxvvnFtVF86DUl+W8hP+OLncgLPyI2UAHAT5Tl6llAN
6q5V+dIfx+/iXgzgQYofb8IovjJL5apg/rN2fHf2HVzWRDuZTsvEQ1FB4+9xngO+Ffnyna3i1zdw
pRLPJk5+8c7AlxXpqpoCsfcwnMkGfpiV7y9M54bqtVMe6QCCZ64w4X0wjtC5d5SVydFGWH4AXxv1
HgjU7128l15osmfeFa2YQN5v6tgXjOiJGXl4v8JOim01X5YNouNrit+35qRJ2Q7F5YWWNjzNVPsc
wSkfQfVxEVwX2t81A9uwXid6tI566WYuy0DIMID/mHp8u0V2uYlkPHjCFjhVNSwrSnj8qA/qTXXP
iIVsbHf7w2nwOXGNUiC894gw2GiORRj8jNaR9W5ODn2M7JLnd0o83pjtF1xsZrx8xBaXo7t8Fvkg
KJXGnStDkhNflwLV1oZjX366ncMBS7l+T75HxsYrttTrQf7w97nz0VEqojlEgOlHNxHmd22F6Vjv
yETUlDw1RWX3rmUCqJVY6a7kMq6zGBYK3TeB18zP/KuAvwt5gVtSshNNLsmqczWwDyPnhaKmXa5/
oZv4UcyN6gedL04KxtxpbP8of1Vb8EBk1DOfNmtv+uRQF4A0QZ9N5ClisCueKOgzUP0httbcoUuf
F7/bxUO7ht2xJRWjfd853eZHx3HuiDzJVcV+asqd24oelrbM1gA3hJpsLlz9iPz9ij1vexp9wW44
2gtMV55zbPWMH3EXVf0E3s63oGxEjva2kP/nY6sy+a8/v5Zu2VhciQWczh56jSmXFDUsnYgeL1J4
DgUUXV784gqrk1p5kJxArOVmfqGF45JKEoUrj/l5bc8Ao5yaxtVWVgt6OvTv/Ei+1S48++Ha0K5j
xJD+48YITo7IbN31s3yl8OcaVwnjODAD4PIzrXg8CAkgy41SQYnaZpAm+Dbm99z7UPLMhj+ymlKv
YGcmUQx/I99Zxsb/gTnltcScT5tfW2BwlbLNcpo7INNM92pQkM5Ut+ZsVmdY4YS1bi65vXytHUEr
7qYybiC/5jPYd0pfh/JxhT8gg2T0g2JWC42nZbhm3Ow5BKxGfWpihDtxzsRWLJ/wVMpw020OgIMq
yIq2h4/13I3T5IMvQArL8MUfelzlrJDSyTzvrcD1fzvyZpmQTW42q1xgKAL+qiFw0EYP98Z63hP4
yaKSpQ8uxKeSLDt50S1DQZzJOXeefEXIQXWvzFxPecaX4s6rjhCl0lH20z4pnRCtm670wqSPIXYB
p9c+00egloNfcLGFCwbTWoiTVsaOe/1PixrVyezC90cMtxTCT4CasRH5S+1Cd0d5h7QHC49oTEQb
IsQOlAZkOR/zfFkNMFjChrvOH6k6aDd1rdM/aBhZC69yfT5XEPyashMXzLmzyviWwfWRYDpNH9r1
eBLAsAFDownbA8AktXZGRuxLNoL+SCZCEnURbJDe/Z0ooQtdIvu901pQ5We2L/dWeUgIQzGn4cc1
O0/+nKz/Bw7q1v9o+ackjgW3/eqeQ81B4j0bSspsOUPQMUmNKwcWqU74xPQPbJm4KZl8Hu9SWeQP
MktSh+QzJeGGZej3V98zwrMp/tq0HpX3noFCXw4kP01nSY9jyRvLkQYBg0NpN6E1PP0lm2FuVZtp
2plBkjju8V56a4bQAt8fcHO7e6UbEAL2OyIBRU9bZZBbtsrDD9R9lO7JCU1sMG5gB6E1KW4F3nDT
uMWrlDqCoYzYLePkWs9eAQgxypiIEgEvBEc45hqRVeTCA+8NhNCAPNDV49IBnrUpExMysLqRsgYZ
+uaJhVcsiRA5MdfnsiIAWe7ZqOXbt7JJzNG6RHEcFZ0r5jur+5UNOpYUYrF9QzGR8g3R0xevhLOO
jz1IqE884GQYhXq1bQ+HSr1qL5wTNHmhM4geiSJDBauJG+07C48de72Oh2+CdTABtrM54sh+4TXk
4UvNa/1Np0wycMyqqqeZhEzB7A4b/b7BO5ye4lnX+eSuhDmfeyZEodGWNsxd+VH3AoK5p+pDFduI
LuMmXuYpN874i3z02EHN+v8yiCPbY/oPjg1ey//Fej1qmgJwEP+mc0ZPEdOcay5Wr/f09J2UHTi8
UPad4jVRJpb4ylUxm0xbVrQMa49NlSqRvat8ySu8lrfVvg5xecD4EmL8Lv+qneWdtva25Og4apY8
FfD9KQ6uxi1hEAfHzk8vnitM+BknCPplXtDIwB7F1EOIwbRW5WaC0QMYI28jWPLCkdOG+TWbafnc
efe8tn6tymtj9cg8r2Gau6BiNeBxTBrjC1Ezr+Qv2TXUwOEbMKxb/QU94/14Z+YWRLIqrW7HqWW/
iNMcS3c0skV1eoYS4pwgSA9A0JREhvw302CVuse7e0TQv/3b2Wnwv9Wq0fnlhM52W5iRlCQn2HR/
QvcwINS/6ZZXHg1ZBnDn40BQDRE7TiSEACc+IpefyPNBu68FxBY5sajxqJOkiH+eNaz6KjOg1IkR
b76HlaD0HD/pCwxTlKI4rTOiFb6p2U7rQR4AwIYc70gpc8hqQAniLsz1fdNmqEitnJ5Ju74pkv3z
LiHBCZ9W6GGHPMqqahvOoAuih/h+B1BhbWart6JJOH9bP0ElFmjijDqbwGZ7RYEPgzb/8gyabSny
tziOvb+SFqfK/cjVKzz3i2ntCEq3nbBhEpKPOpKrm2lVbtzvf1Bzl9QyTdXJlbA4Gu2zqaC8Wju/
BZK3E+cC9qM9BJ7mRvsBfxubydQY0JpBt81ei8PVbMlYr16P7jyiCYZNr6KTEdngw8lYVBLhoXd1
uFMeqemvbLqlkS9kfSw/A2rHYrIlA4l/K3ykMx2Qu2lFeP/BmAvOEMfJB8vPalZ8WqDUbQYQyo6t
HaQ/W7hCRKh8ZYU4TQtBSHAdeRsQj4/+ngBlW3vr13QsPGP2OPqZ7Bcj26CUgFkIXRGykxubF3hZ
7xcNryxhsDVwxRL//Q4TCnMKzqjlEcU99wzTt4UQdBqsy2Ptq+rG2CuGPx/KKzkEZULpKGcU4Hgk
j0qkGoV7SxV2Rfbgj8xsTAyRt0nTl7UF5s2H6bI9vjdpF1U5671sHywRFO1Ox21pLyRthEKWRCr4
qoa7/5LIOqnSH2XTAOYGKMqiuOyAs6kjv2sleynUNNJXpdPD6mzYFeRpioZDK8HnwvYG/l4rDaBH
tdgWnewCcrX5TqyTnpGcISoxjHbXGhjQ+JrDp3z7plTtA331UwNrxVpOSHAK2R5ygFsuEwId0Vm4
8bLi5iJO1Ajk5Dc1jXrw7HFLmJ5xD0Y6hMPHDHHD3lFXZ9C4QZY31aXIXRd6KJTfMGFCgUhvEAVc
q8XK+2LSxHcSt3EWnAWWUpSUUF4AmtJs266AnXMk7Mfyrnzp5gao1ws03JMGLY+qgQLY8Gd1QaWU
Q+wtd9OKCywony8jHlp3P+8oBO4WEQF054tSJNIPcdSO4ch9y+IDJKHlIrSFIRmqXX+AzP7NXisV
KFirhigEh7KZfoAS5ezUvGASDtn6s+MLjmD0JW6ExlZyVT5JBhyv6zcnQ6HfLRF2wXr6x48LkTcD
OrBQqI+3A481hv8aF8ROanpWuTMdQvLX5u057aKglwkeqfQ0r+lmCmVB/wznNdVlePcASUzVPRwF
Obv5Jaa4HD8kVnTJJa2f+kGJRagfTJeFu/2gE0W4G+kAc/A6nR1pQRPtno+DiS6Z/WszisCOGgLo
VKLAFiokPxYUap3bnEpuVkM3SH9TJZMNHiKoeGYh9Lt6k0hQio91bWGHa+kskGbV5qi+RwkJ0sRw
9VBLSaWdEH55rTbfhn3aovdOyOI+YUBxF+OLMrcZMd74Xy3VgC0NwxMpSf9NXeSnKv2rEuUhLDrs
6ZChFeq5S1349PQyDizd0dI2Tl0PCz7g1bN2fO2Tf8oXGvTu7QGym0wBXDdKxZ5EBs2Ho7bQBBoE
Vv2f8sICBcp0rHZvEeNVTnK4uYU59oa1ie6VAEySK5MDw37f1dAb40qRndTvC9C8tbVjr9cw1n9x
zJWQLgXOHXNXpX1bl3j4vnaaWBROikyLfMDDBCOi6B0SrtYp6rGTLLQsBprZiBbDFOzlJRPafu3T
zApJbOaJgsdnH7JoxcXxxWQWJSpTajnjt+keOWTVfHqyeui2LTOU4HMHdbi5v65zCPGfZy+q/VgF
qWld7tf8ax+lTWHpqP4Fpl/vCU8n1VHG7lGojgvaqIygG699DtSrcbJNh2dFUH1Gig8USH7BQo/j
cTJgLPb3IpE2OXQKSND4GwLdaIEEqpBHjaAgBhlkicAl4uGTgzl0imlCEMyjm4W43jRSOz1UFkic
fzWhnAuTCCUDfBVXKLcgXQg7ZiGa+QvQInmXLGFXGxx48yeFhP/uIwBYZdbSGEQ+vR/st/TCQ2jN
kQz2qNIGOOKNPEVmV200eMkfLd6CVcdITHHtwgMhvlcu3dzHCVa9XbFtloH0MOGn5tSfi8go9par
YUIev1SBpjMIus7NcXIri+8xd/Qs6xpVgFWqSHojgCYJkCmuIXlhKAD+oYtUP7tP2waEVEbGl8E5
y7QlJ/4W5GXcJycPIAFQ4Xg4y3LJvY+m97+Pb1nFSLqoh5YxdlYpoM2GnB/RhPizlU1lhTcUzM4n
wZBQXv9MlzzQ8XCJ/X0z1NgiLM0p7nCZG6vIQNc97kluB71dIqguXJBsXUvSbkRcw0Dk19uXEhgy
NgfOkZB8CMTLIAkYMg1pojU/Q2J+o9lvhA3DwWiSB5iGUXGzSSizuKeCYP3BdsnStkQJCRPUH8il
1TBkca05KgxIJA0+x0EIvToU8lCJw+SYii90W51hYKCegAJxL+6nslSUGCepHmWncc62AZI2z/Dk
8ZGIDxSupuwZo2mukK4rJe+9bGQrSFnqhS6erd838J+/N3hT/SxR9fXVdisjPbrU0buaSuzMqzC2
YN57qsUiN33IN3BEpeImWn3JjLOrPAlQ1/aPCp3pKrzLBfUS67fo46YCydVgIkbxy0bQUYGYbqF+
BE76VG2DPKYXOFrFb53ZIeSbebo4iS6DeUFSVjwEUgEl1q3CcVg0vCsj1t5tV5ArfIx2zsV9i/Xb
77hTmB7MZwas6EIBFOf5F31TkRBIPnz5bALX01b/kC2riUlS0aTMOTQIeQoqSkE9WXOhbkEC8Ozb
IpXLf4h1lZ0W/mQvC5A27u9HTQFSsLvq4+n5xBxQG/og0ceFHL+tmkFRmpQxxjM0nwnveh9u6i9n
iQrFSXb5dTC0JIZXyxVivrKp8beegK7KD16Lpgi8CpR2YAby7ABSfb7x0pDSCxulO7AbzaNQ5XV5
66/YPYVqFsA1ecGrOa5Okqa6q1Hy79hWfQPJM13yL+36bZlhK4eKsmVlyIj5UqbbUEkn22zQ6dQP
OLrw6j+GTrQcLSk7bQbBtAFIF6hMq1QgyKX69A698w9J61hZz/wrU+0jWZJdAoNNUMVwl3Az8rG8
0HeH9E+exI9EiMT8fBPMKeFgFettb1fxLSLcfHA2z+LZo+Z+M/qK58lGBDHeuTqFZncZduFb0YQp
tycT8IVN8XQ7WwTEzivRegELjJz5NlweJrMoD1yWEQMqlPl+S9Er4ejzyeEB/PxoMeoZTG4F7oKa
Dj9OCF/LuFUVY17g1N0kBnOZgBtUD0Zk1qUidtVuwFDuBwRRDmJr7AZY2pUhrALaJ0oO20dmRY3v
Ma1Ivlz2w9oPnMDoZP1p0oN9T7p2757chHNKWgF/WCqI+5LUJUEh9wMVOr0zkfFZ04F/3aMmcF9a
QBXaP+UTXU65zfSDGzpmG2NY1X0llJbRk0MzYfxcVok1HDu/rGCCTxta7F9p405kgraxx+fFprVg
A1DiI4JgA1hU9R6ieG2BirUUyP3HzJNiS0/py7dqyZDi372awEYmAYfxFzH/JG0HYw4HHtiWBSyi
FNnFA97UioyzM8CjcboSBLYy7WT7K73j3xqYSyKBakM6pnELdR52jwDqjbx8nFhF3EDwjorHjpG8
ADQ/2YG7NE5lgsZSGenuQzOCPnBYVkYLkUyaVatzOJPo1hWltvN/9m/UiSGOMlHe2Azg3RnyXUrg
YWMXO72HvEWDL5sjAbAOeiacADPHBmzsdxEHkL8hlh95wWQ8fS2uLK/z9FDz9KGL8x/jD61UQsS1
gjOTko7idkiQRbH0cYGe5TMGhIxaiX5Dnj/hPL0dtemb8IQwOxeT14vg8BpMGoCyOVnca7JRSYOZ
IeeldlPkU9rNU5QvOHf8BCXHoqk6iwiZbTqHosTc8v+U8UUpSP6LGKcu/CatJZZhDDyOvckq1Tmb
8qvUyY3cHiI5O08ehVGr9La1dGeQlPFjECm1hMxqt4u5TDH5wRKUIwr/5LNogFakxFVG2Ne0hs1U
dwqvmIGqMN6YJsAFPXDukywMEdLjSvncsbvTyk/VpvWecR9mkgeEMMH1w7xX4yCxjNyLXG1zlQ/5
P7j7oXApy7keQVcOgl7kEXu49OzS3BcoTFtWipq/nYD56I6Rstv6DwdxpBGBoJxctSp9XSaLdOxt
HCNcfOr4W8AixhOGeZvTiFoWHTolBhjV0bLKJ8aLVa8VsIUYNtpTb6cQL5rrRTZHWKmAons868xe
rFkzhb5TzeJLNgU2JAZc+nnXE8kSHrms9WNMj3eAH1oFVFD/Nm5DauRKIgixzn9STdgszotMummr
wHkgoG8XCwDNUcBiggduzkYuChU/ofYBDj8lDq31/o097a8qvD/FL01P3gQYGUb09hfpx2pxEbIh
3yBTNHwVaeBTau8Wrmh9BA81ke25NxKu97ZNsHuGe9Q+2fXKDT2jRXhvNssLH90E2u9IIoIMsB9x
TfOvSxtiqKVW6tAw4frdaHAOr3sIj87ewv0lxlZ3uFJGpFwz/0gLuCzfHySZc0jtEo/hmIttzCrv
+XfiA19tnFm5fldRRMy/Sgp/vBy3SjsqEeD8QMdEWgqW5n1Kj3YL11OpjZUHb6hEn0PymJ9y20QU
MPRGC4KhEh6ByJbnBUC22gS0TTTdkilLutDJ0/H8I1A83Dt2zYBzUo2KPhpQ+SosD9pTGNvN3l/N
f02sqewBukl7M7xDIh1GvFLESh4zihXKPp6CjD4zMwj0A1BBuJGiZM2nfAYyEiPwLUBooqDlUDj2
RJLbMjKOJeZxdQaAx8H21q6XjIim0TKLd8PPsH+C6uBDo0D5KUayhpDuldczRO8Jk7kaoiwVHdbU
ktDVcanLS0ocD8xF41GGM55r+BMRFHBcack3Jaf6YF/BuetsRY/l73/FjiiaVtmNRp52ZA/AUBMD
fSnIQ6+kuXVTpBkeu+B5bENDLGzJoixWyMXV4z9hvyLIPZri/owrEYQZLTMoC4usIqu3ukeiIIag
+FmUpyG1+m8zAiEg7Y3KPPsEu1/RwqNsAfoizwyCQqQgC2d8DAfYpTJojUQRC8LoYeHsGd3Uoh3w
Ek3kiMnqaQjWfu0cLKTioSwbPfYmufLDn/LhVIN+cexQoCsq8BE8+UEdwCktUo/SgPXMNzxFcyxh
2QcR+UHmT7Phe0ipIE72G47wcL3JRIP21pCFzBkFkffTbBNdLtv5NcwYrPnuPYv4XuVYdjWUdVyq
Ys+K2yjsvd4nLLeMH+EziL1vHKdfyvaMGq2QP2XR+m+GXmIoGN/rwUBZS788uvsHfobk9K21bMVY
fLOVQSP2RcOJEgaySIY07nvGZE6CT0bPRlOvNRY/mcbYjSUlvpGNLotZWAsbaygwRzcn6+KgWZKS
QL/8LgktEXZ9dS/v50jRifui8cMrsaVzjKkdkdZVfaiOkrzFAjT+DR/2VmtOKCh0S6h/rRl4FkU+
VVfapfKjwYYJUC2N+oce+TSlfVp6Z5SQv+DGZd4nOVjoUqAcFCIwAZNR/lgeGWl8T0aMBGQJHNQD
o/DTCh/yG0/RKd7YGoGI4NUGyCWhw6rkz+r1ZiyQR9ap/ImdHKhRwnlKo0e1s2h+pQkFoA4k9S8f
L5DO93S8tw13SFK6Cv2+tOh2WKoUE+0qBpnwPrFM6v4AX/d2ms0jRfsFH5PCGYzDprgTB+kiw+LY
9TeeZ51GuDc7/CeFsa1PxuDBVynS3c9I9TZYrzHd0DJuUK/ZZqXa0IkqPLSgMQjLQ25GI9ctrPzt
32ObE3y5QRgKxC3GWcrLUG88i2EcgdxFRmx01ojltZbyfogvA1d5hLM86hMBYYgbiIffgJQZrTsg
873H9NinN03whCLaOeisvOpoYfQOJrwl1LXHbfuaKYlavG/o9wUWDr7eViIbJ4xgcjxtsW1RE2aC
MifOmP64vkZPL7DyK0RUyEsWEOxD7cD844zajLvYkz16K39Kjsj8BYsrGPSjlzTxTN42+5r8ZY7i
D2VxooTpFgB1y2qCEM+7MwnYukNmmhb4yl/N0qRwFagZZpQgA9P13MirkC56YqggfftgKLzs+jnB
5vWwpOH6gT9arfnGLoC+GVYRqnPK6m0tDI0F3NR+nxd1SuAQ+oyFM+7EaXqz6s2id1eNzTSdAWvb
gyVHB7yuW24uCnqTjmi6PuD16EsU09QrB10y0FwP+uOoHsgHrcpqhs89QCOpkxYfPI5udf5Z5eWs
Trk9+hBLlk1G/sq4asMhFXMqb5dBz1N7JI4iYBIOcZ1/3j7M1ScYllibh8xMUZHlp5EraSrDhdcp
1G+NLpF2mgi9oDr6qoij2i+cdyLOuHP9XdWCD/wVbjdf2abR7iG11QzSjkRsQ3080iMB0U9PhC2f
oklgvJbYf9U9TitruUVJspRrJWhXd0ckhHIyJM8BTsqUKEd45Bx93sXtappvENITfjaT/v5TcPIC
Gb7oOkCFmn4o2vm7t/qsySo//1gw0a6Xs+zHhFrdhXaUvXBLOThLEqKumoQIwg2WwQL73UxDkE90
XcgxcmV7mlUx/4c3XxWDnVRm+PLi2JlvEAboB3ivx7nacjdFsANffoi0qfG8wx37Bl8cYIb4YnTJ
/G3RK721vtC37tpDyTqXj5S5VbhroPAQ1Kc24PITmkpmB8o1Dewe9CM/vjUpMSSgGiG8eiI8tnQW
RbeVpRyPkYf9dHt+UsqA62dO0TE1Itojfk0sSwKsUH/iowEC6RUKpHqiyM4PCV9/mAd98V2zD+G+
aP508ah1tRZB3dj/8dAbHhdccZyPJBWzlbtJaSVKSZ0euanS0ibHW948zEzlhhxW5D9OyxRijLy7
2ovSJtnilcjClPaAnuSgmvovOIWNMalUDifAxLN1WQl6H1XGOAWtEvDcNbF9COyI2do5syijKGbF
cbT7gYoM2o4KXDuNJfMPoketmhOiIvSiLJ5Gqx1sGYxyU7P0mA8AY0hPEwMFWLtE99oXW9/ePdvV
YJhC0LAeqwpsXVrZG7/HdaWqzX4S3GFGhfkoV3jPY++MHQvgdelFJiRmS3I2jbubzX5+hmmZVH2Z
4fZO/0jTL/SQC3D1Hi0UeZtnRyuJXMuanuNQS1F3LiPm/nKO95FyJNfaPb7PBQHsYDB0Rj3fg/3P
x0qygVSKHUIA4nmpTHlIKV5jFpUmlkCpfw4/z9g17yIP9Sd5Y1r7Ssm8t24QPCOLiMkbJWNAqHJg
dh2X89GnVShDsuXQoFfKiguZ1YyaXBWTJLeCEXqvARnNJlZDjP2WG2G2UP6hw4vbe6UJO3DzZBzQ
x/dHBDyaRKoaR4DOzVd9J5nDkQ9lI4ldHy/RvdSDA10g3a0HQ0iNyOVozyp+QQQE5An/H8515h+T
ktPdtHHCswCE+PtcLoPiA49IAQdihCwuCBPRYBG3CO5Ce40h4dN0z4dgFctgqkEA6ZpEikFS8qm5
OJlLmYB5SEpAFjaenFM6XdbLbXwBD/+5PomSaJ0Ecef8Ee5N2h8elJaq1uSIDRcn2QER1WspB1gw
zMHAo96BbDOoMvEda6RFCXYkxjUXA368c2m0XKytIjgXKmtF+2IeYf5BTsLCbdArWu7L+gUQEJjM
o14H2o4PXJE/+wOcbQTMThiRgdRrY0cNFqkxlZKj0U9AFjMQMnCOMXSXwnUX8cnlQV53hUUnfxsZ
9+4IsT1bQuA/mUv80qxdFea4vCgdE++wyfvoOhpXHEETkOt6WdM4RoLZd3q15olAj/ZN+Q3rZiD7
T6b3gjWGG9ePuiLZ/qIN0DaDsatJk2vO/ULBhasJeQp4GuzU9fPDF1uC6unQ8F08vMfcjLt+rUaP
6jMkwNkYR3SBLVGS9xnyqAVk6/wwzGJWZijeEXPAN+dfKAKmdFnrnQIF8cfo1Y+AOTo4NpQyA54l
4YQjbdfh2EPN2fj9G/NzJ7kcikBkWGcN8v9txWqQywyKEChnz9+R/FFChZL2Wath+mTSvKTNfD3m
K/8xqA99MWVOKmNHlK5ArTPHcxh/7+4grbEIZOjCOxACUqcoBHWI3AaScs3kIQ3azCkaTyQl1iJZ
DqHm4+0FVwRCnOrzCjB0/4NOHMA8d43wrQGrnAD7bD+ilxBM/EvKthaj+yP8rBIRmxlgrww/tYrV
Z8ziC3dBHNEIC8DMZY2pEoVEk3/d/oNzqGdCrmIIb5ImNyVlqHP8O5aNHKvDBs45duat+CDsk26B
5hNGcZeWP5fUsAFK9CeZm1IPL2kGRQUtyPACcp5Ni3viXkgiTq7hRpu7x2WrPuwsJgRgQtwZJrlW
ZbK3hYuIUNViVGdf4oB9P2Jbz8SO/+Hr+X0B86XEPY91huHcvusqXS2ZvH+SkhETDCzYuLzaQv/m
OHguujHk08Y2qiPLNrOKXuvE4JwuRSicu7BfkvaYQgVIjN4q5xOyudyx7zzm39tKG4eSb8ITGqqx
Elh1d9DHabbjgSWUsP1YMaksvCT8pRedG9l9kSzwX8vuico3whVTRHewtriptAerSKkKiS9CJLD6
WdHdzNnrAgviJYHSia3cqnn/lpyhHGh6L3z8va1ytzM0aFUGvYm4y+SnqC107Xuj7jWaHlCUcrbI
HdwXc268pwBDvgj47gqcmZz2bbqmp0/x4O3ZG4J8lv7vmULDRNLVCH+qZgiQ0W0D1izE8PS1s0eS
BaSyS+JGk7BskITF4XOfvtweXaougaE4xUCE46nH8jRT2d59igDactQpJHyN07JN71uNQdn2MWNI
iXwK+wnVtMHW0M5n28s0p50lO1cWkM5ocEHXJJ0nzBsdV6/6ilH6+z3cMNSpufnmxu+20M84Xxqj
x8E2G43uwG3Jjrpo9FynouKG/7zuunE1YVjRK4MwvOX2O2n+pwnd8O13IlP7ckV9g7kNn+vUPCpf
SfcQTm/6CbD70I1k6uWNu6NE/AwF+dfR8I4gmIAhmHS0hOU1R3Kk+nJHFrwFXlg0Pr/8PkN/L/tT
pfCdkC43/q/5sLR0rCuQr3REBNz3CrLi8SJ+RBk4NgJD8Oygz16nX9jO/7RTQ89dqKjNx4rATUo6
RzFcZhcdADofnVVzbntpIX9Y3D+/3bv7Lz5cV3YCfO6tJnhZBUOj31Ohg34tHrCMAZqNz+EuOZYM
yyWjqnRmBGsjlI3HL2o6GAYMwKQTBLF8RvA5tWBe+l0eHyJeWdRIx6myZ0xVjTXfjPHq66MVR5KE
onwqv6LgTD5VZeMoRX0OaiTP4vcr2gzY52vBblX5bTVI/Wnw0CflOQBXFFVWVVKk+NjUpaqq87fM
XSh5KEt1mLU+cERjb8H/CiXKWsF9/J75m5MJNBLiGPjTxQ8niDXT09Fkd4aS5In5GjYvPJblu0oc
FN/6V973NiZpwFKDsmE1CD3BNDXvw0SYo+ZlLOp8f9+lAU5wT+H1upc6pEl5Kt9OAlWwAQ4DQJJ0
uMFmSAsFqh9DG3b9xOsPKh+g+eOc7YBgvbUSTr1h61Xd6bSs+XDgKeZbB0OpznxNFZCiZwXR6TH5
DGIjxfsDSFJ1Md1V6+2uhxRikxtUPRWr7FdcHhvNmC8ho3gnmv1nL2qUs7U78iINquKfZ6haXBYi
4gtQBLWnB1QvmVr+R+TVCC50V4MGtBan4c6RqyrXbnctx/tIE936XIRp7d/Q0In49uui2GIrbhEd
VisCqp399Ibqr50yPkJB5PakkhzvOn5a1tr8myGm2FnK1UUAwBcUi34PaU6Jbd7PtFEDLuRuIRfc
1waZNTpTOU6IADiAJylZ0YO15eklpHuz/+AX2qzRUSagC0hYlCjJ6DYmyUhDyiupuzf0Cr9F3XAc
JaGXU/GJsrM9LXfiZ2Tp57vlBMiQG/9YFTIQEw7TirH5FzjEVUs0r8iCq+XoT2Aq93OLqTP4/mqp
irGiKpHkYDZ9aYGPnKjcMnzY0oC57y0Heq1jPvsw7j8V2JjD/IyB4zAsa/3qwOLgCHHP8qj+hUTG
5BTyB0DxJuH1dVUyD8NuL56JTF7zvxWmbNe92GSPtrSpl6d9YYBMwjo3Zju7NlkN+PLG9vyvryIz
qWNkz4Dq7o573NY/PsogrcfGe+VfBs2cMumwMaWlP36MYltb7oK3MfYJ3Rpwh3WNWxEZo0PcyNta
8WD0yXUAULUe0h+uAoo0hsW12YlGoRBsebFYjh71Z/pgJehtRGGuLcnom48szO8lHGY/rW2luwFN
bSNIYZjUCqt3OajYlIpShx8/qMntIgbWSKLQR2JOaA7MzxzHu96FX6qMgv1haqTqeC1IwIOJ0DSC
q/DJcF9ZxGyhAMNUoYzQlcYTb/BEVl9Fzz2YXnLOus5x825SVCHWAr+e5ZX5JoYwYiXx76IosYCG
CIPyVlsXYXJ5QA7G8aHd//V7rgJ0ieFKGbi0O1YOrAV8/3nGiUfTlCaEuBkmEIhh+eKPDV2KMC0m
JomISZpa3GWAcg8eWivKLYEXwmEAk6OaSkblH1KuknBLN9BVcDzj02iQ1hn4kdTq2gZjHR1RfGtm
Xjs0y1i8dAWkxdI/FSVGIDJ0ibbGx5s2RXi8aV5Ai4g4mDvbCuplWbUHDMjIIbrl+LNdNyGGhF/i
AsUf43d+vBQw96oCjG0rRw1ELoehh2v/l7uYSYvVgzx3eewA/b9/XE2MQ9D9k69Vf2vAa+LKH0vE
iyMOoM7UgG3V6/cA5kgQgcb9nZeCvPEOKIYf6owhLgfkl+YqaiapDptG/SzwPUOrTr3A0+jwNowM
hbjqgb7E0aGpjCygly4S0m2G1gcOsul688AqukMBgkFWSTpeNBWeV2iQaC0Vscj4H2BuGaaXcj9w
36aVN11gtWzl2z3aW3zWx37lVD6tIEtTXJ6sBJQpOEKbWxMnyOpcPfpAQOOySLMcwt+U+mT3lHRO
C0CmxK+awUCJ2xieuluNMVKX/k4EsU9qEQYn35a08qkDnTgHv0U/FvhJAcnIsJHe7uG/F6TBNg1b
cN64v86+GLech4SXRLFsBWtRBu/OLEJmzUQFygJyRv1BOLrHtIr8Lex6stnu2glyh+om2xucNuEI
JjM0ouuVCCGzWuCg0Q66aDNG0mLZ7bEzcBMTWZoLc/5J94Z8JlRFVkPTpmesDIB45eiyjxCpOk15
CDn1AUkjCoU2+1ZzC3NK95iuvRZayFxq0SJq+MyHpP8UsxVMsx6e09V04WsaDBkJwodw1yS6DfH3
xW1SMFcJaENmL+n6l4YPpffhsTVUJd4zKzm3Zm+/oiqBxkr1wtrNz6bK7nvhfHYC7llbuTOOewfg
A/t8PfBrNRCidahpeCKhdv7dwNaJiU63B+QbBlGN3y64a1hQK24Mg/Kre+4V4SohS68/hKF1UN7+
YxlR50Z3KfN8EdsEu4tKyhv09ymT06tInzkw+u84Pr/RV8L7mnWgaq6taVheTqzON1RVCRTBGSRV
vv20klL0F4h9Sr3TFGlhwwRjFHxM5z2KPg99xKGmCZJeaClDFDHaOwt2jeWQSKc9QiiZZTM8GEBD
B1z/WzzBgX7U1WnRaKfSD1WUvp4UhHItlmS/d/7g5R3aTaLsgfmEY6yhA115qTQmpkq7tPYd7yOL
/k07JNh7av6ZV6Hs3ei+WloFdFjIK5ShC8tKkvtvNK8Dw6jJQ9NTMg2+YmQXmacDOB3Xb13MiyPs
0HbYQfST/XjhyYSUeg2eQ7UyeG9RXXWPLrnrzCx+H81shouHqU9WYB72gT/CO0wFYNKB8bxU6bLr
xBp5lIro4k+3kOLqZstqhFNp6ZxS171jeYN8e/MPhVgSOrbAhad/JJi0qeIFod7rfAWK1MJvn3zw
6usLKYvApOprpm3QgH8RzocJhHNH2WqY3X3utL/QmODyQ3XU+9FMiq+UZ22KxvrzUnVFYnbF3/sE
o5QRW0Nhoh5G3bL+/3dU/YiThHIzfM8qELdzRrkVbGBHO1j3mims2EV4LwcTVvk5qbSOoYOIzirn
5l99OzBCnbEcfcTOLgwUlnakMZTg3uqsLjyoBlVrGJ9nNPuHJErUNf+5jCvn30ByOZHbW5VxQGOL
TfXbWbLGg6iQ/jQlzIoOzllUbNYRSu07Rv6qvKHxGdWtp+CAr5qe2lRP0Jr/0BY6hVbIecYzANRk
q+kljqRnuDUmkcZ3qoEO0qnilWHLLKYcEIN4GodIqpp2FYWaaM2rCvoiubjSWmRjMg0eYKnf+elO
y9Zrm1nmaZdrIvX6x/72U5kAWDQdsShdOC77ZLi9UsDo6ZSbqFaFeiaaMhy/pnabhlIHfA6r2uGc
Jv5934h3bmvdmLbOtQvU8VuAAws/fzkAmyoCypVBN+Wr4HT/nW8P0McHu2l0aOxWzr7Z6k9LjNkC
Q0Dn7GHjMX5IOSNh59dVZxhlhMxxQi5avplsHRbyhvIeJL8/EOOTCx3U91cp5His2zcdUYGv2e2J
+BlLM6n30HmGj0hVKphyTIrgSST+dE2jOhkRBnxGSCGK8ljretsqsfb6TJKNgha7IXnmyfOJtWtu
+jApDqoOrNb8EjaM90RqM9PKq5rXjbAhj7aUlAf4wefXMZvc9voCjeGQ32sge/V0XuZvYqku9cu0
4ToLLBiOMK3GJ4PWL3gXpuHIzKupz3pcUdh+/fwiC8j3H/07p6KVPYe50a0grRDN11SJr8Sb66p/
IsWV7KpqHwpiVNTScSJiJVPAJHHXJonzOd1Pf2LCFPl3BDixMYNW03eKBguOcEec1UNc2XRhTstb
d316KMgr51O6vVpvcnUUFPnFahMskTSAyt2YEg5e7nPGcJF+FHa02rIfCKhbzrfg77z0MBuS5JS6
dnHhd9htuM9PZBxSReTtoHJt3b/J1AJhWIW8sg4xP107JUqu1i80ye4gmHr8pQ9jNK5NRtcNPPOR
Yvhc9Re8SgY+1In5Dt0y/rigq5DCpFLn1HpsND8Zbyd4KFlZL4sD0ie/GGrurfWIBchXbez5j6oG
2GqEI6gu7LOIXUvLRIy+nxA2Ec0UYvxv4I64fPNLNXZ+CVzhha1elJldrQb/O1SZ6LDVdm70jWzP
rzqT8sGegqJ3LUEHpUpy3J2e8IMoUJr1EDGe6uEaVcBikIUZjiqYBdvszPGVoYdjDASTz5Qylqdd
7+KdRY//eJfQuCvnBVIVSJoSyhoZ9RPZyMuChUgpg8OVxQW05tFVSVGgCh5PXlQU3vWgzkqoDKlV
Czv9/PmnK+cFdqwIg6XGiZHXHzgrtUrmOJtraa2wQGJhxHWT/T7JC9CwDeWNQshpnZH+b0qbUGUw
YiX2RW1ubO2EfZvaxl9VVLr87UdoRAl1tzoc2l6UdOFmC0L/WNjnolw1srAG49huXEAbs2dh8841
vsf97ZHVE8hlnWGFPNAy9d2zJktYnrCuYH26Vhe8mLac5y/POyTp8slNcpBvYPPPWh/ou1Pgpgcs
F4iHW1qbmI9s8GNLAGgY567Y2e1bo9Z2CI2ZFwWNWG6wjTlTGipvZLz2AXXQgkqO5x7OSpX4yha6
jjf76yATloC1CDwZIL8kU3Nfc0mixMVB1isfGhDYhF9df4Xuy7yhFwu83oM/m0qo7OcwUypgyu+l
Dga0JvDJWr6d+z5a1NJIauDpN53Sr//28NQCCffY3gkdbo9/fXsR6ZUEjoSg2RIsiefNl6G47PJd
50XSYc61d6djmMGdV8E19iO70IdJpKn8voy6RsInBB94c5+Qo2n1+pTZiGaIdnokAzqk2nvfERjS
I0GXgimDoK7JeZdxvguEd32dJfrsjFQdetFrC0nffp3QH7FXjSthkgtuHJOo8/a0GkrA87y0yYq3
vn1amTi6oQygqzxlCnxQUlNoBzahEt2U/jgsqWqeU4m9TCsOuR/YxkMJbqTBxNR1o/dzfJty/0Kn
kQnFKl6uyU8Dsapr/sVF0InDttWWW7b+2ysjUBfZcqU5F993aSZoeUAfynPHhAJyxx50PE0VOo2s
/PAPDRyppyjc2Obm09ZL9/HMBBiKIk+fyaQjCJO/0Yz23xf/LWRLDOp+IQE+S6x7v3/eUOBl+KQa
BdmmJsPDhIqaBftMClppEXGaT5FY5K0pq6c4o+1MRWvzm1qnkLjVd/ovSJfN4wnIyk128cq6vMb1
9MBVxLQKhCmGZR6CeEpw8peJ06PawqtNV04OjtgTty+cI9r56OqzL7vxJe5hHiLf6etwN6UGwAe7
S2Gl7m0wbCgXPIba2uGQUEVXDQvT/nXz3QJXK2NYX4ODf3+kPMiRy3PSr1jt918k7slN1gYHZiQl
CxLnNMb4xi7opVloN9wUyMImG3JBvRW4s5a6ZrTX+dTWuLJu8IeB0RkiU/JJWdFnf7nFUvWS4bp4
9UpVfwgRBnwZFyTp3MrxUmzT1WlP9ZposBBGuJ9umt2pPi1NevmeNx+OYJQYDTBvzWx4xhL2eXUG
gEzFutCZySrkPyxVvmzlOyAZ4dju+EmWrUQehIuMh4opxEjtU2qEagxgKODkYFW8WRwREPKgt9AO
Tcq2sbsNMJtc6hYsasjBThrb4NUq3d4ZUWHirDZGZxSqIwd8vI6Ds9AB6AnfnopqWj8kHY9ZyQsD
8m29xAQtdYRpeAsO8JYoK+Hyfs+6XYc9BSAS0rm4RueNXitIk/rjxPQ/X1V6mQDU/WqVuG9OdOLd
tKOV7nV/VwLRaeuTNcyJZjXgbbE+iXk4bK48PYh+fG3XjCfI6RMQOhBmpUhgqTvZ3Vhk22Ck2oow
qumbpNOLcAT857Xzm40uxlSm1NERmAIKGeFZNZi7SS2XU/P4r17k5V+TMYDa+UC1aiOWPX8L+PsK
Hh8QtrsdwwDZ3TM/zbnK6uDYcGa+x/xdlTu53dSWu8s1uhn/5GlAHcvmelUJzxQOTuo3sZ/p7Oe1
4hbraka/kt8g94KJ65fe68JKBaQghy489mK+tbn0H0Bzw1zJdkRuc98UqVXQPfYwLCpFPLP8akBL
n8SI0+nt4+8xeRwJdlFpCUHu9YTXf1Jmy0pKUz0qExg2krfZwlVvIhrvj7f+b8zWhDzRbqXfBvAJ
GVrRRjBqDMHGd6eP2zhdA7d8p1DuIUlTPYLfkOfUu69AUHe2Qr2Y8yFSJ1SGWtvf5G6lewtNpk/f
Wnv4YI2f7IC/7eOOgKvv4zQb4Dd5IWMdRp3msmKmvk63/R3GuTo+8oeWvu+2MU8s3jwFwrlSyJbE
DKbRKqFxp/U8cBCPdmiILqFLlDscTEJE05obSGh45sNvGYhQV8j+/LcXH0kYAXOPjy4/Bf0biEqB
DFSBYze2qRhoeeMLBDoWV01BLL+qR5h8vXVfvSJCU34TLfozkjtvozf5vWeU3nrzEHCsyhCKTMRN
T/3PW4nwKPuZcbnzwRoSIQe3E9nkO7MFWy8+B4urHcgbHx9a5ooQs7/Nu5nUOu+xlUR6iil3Stou
nA11lmWWlB/apvF7Ukjr68ps5OB/ZGmDc3IWgLuYSJlUs3MmXDyOh+6S2Yjb6JKlQ0EN02FObp32
SY4z2S7a5xOUQPsFbtuGhYDauYzbhzXx6KKrTbl4alGxjZbdT5vE2umUNr37gkgTJ60fZh0rM2Bx
SPIRQrifbuwg8Bm6+bzcg9fi2rwszvN5oDTx6bhzD7p7AWUsfh0pZJnxzy1mMp2NXhIFShZpxWaV
cpOiSb+mPx9ymvBEdlhVXVtvotnNfHvQIZeIvfGkmC3Uru4F6MEvn3rQP3z1qjjqiFxgfI7Kp9L7
oPQdyjpOJA2pDS9Hab1uLVrycg/uX4w3Z+3r8G/WFE1gnOY+6atdfhwbCLUwfX27/hylW8VqtZiO
HQeniI7X6ysSGaMLQNvOT+Oxmpq5c7E2ikXgxg7O2kAj/EJLLzPQXQwWqqklzGSSXmTny/xeouVv
gE7XmI5oS9yFtt3+t2Ov/vbW9Per0NVXEBCuDEr90JP0xUajjrqXVZhGOafFf2FPC2PMAvrrievR
Xjqtg3r0C57lnthra5qmvaIjr4SBXHafsofJT8ECuffeOO3SHCqR1gNBlMoC885PdWo63IAe/KD+
taaQ/OypGV7meo2ukJm6vptMUy01SXaghWbdizHRIIEdNasDjmgDGkwPsor9MxS4okI3Z5MlyWTF
S7unrwbes/F+YcqB9qUKTLvwAZWIfLE4vpxAZ4ZXzT42P+wUNH9JSAM2qckF2A6vGyowHdF+xcID
diyDytbo3cauyWkxSOW2oTU1xtt3C+vjk23Iyo79QrUmtTN2C65Ckwev6mltgbyk3Nd4W0eCVwYa
bE0hzR2wOEqrbRDY58IfVfnBCpj1pRMfhjIAk1H2wqYMKCDaz6it3RBc5JRubicUt1UV7M+jNLgL
Qs1Z0+B2rN9hQNUIfNQzU6MPZcUHKccaTfwBOPC6S7BxouGiu090nUJyLrFuRtH+0WXpwG39fk8z
HsuAiGA08CFwAl9lkGF2Psthgwt9fuIy12NurSyA+oxfJf8jigoP84dubu1CUn2Rt+6BkUuWsGGD
m6/NegyaHGttElCUquLaEno1VvxmHr3qOv21eqa7QoSs1P866sks/uatJY8rXk2/zHTvnpL+bD8t
kEhyg7IWIegc0o1UM76p5aa1pHRI0U2v4Sf8ULxWDiqURPxyi67vJV8F9smkk84hNEXejPTCTSWw
kvcYrPSrwvhVcLipFuuKn9QwxeJrGKiusqOdZlNQ3MUGc+qFkE+t8/s1woIuiqLI9EhAZKSSexbP
yO/YnsCZwcrfJj1tgwq/B9FC4zxEezVyweNhUHAm8cAecM/ito9jnwp32Cw8K/Q8/ADk7+Q23wP0
6iNMnotvo64zXedgUzB/+v78JrJ0QEnJY0OKzKnItLaPyFbv/+v67Q0jtq37wSdX0hjmstQJheA8
2UOKfPX4QRUOw95H6MkA9E9VjFHu106jvE0YUvGhm2BKs81XGx7b+j/1eAhEydE/5xngzpXfayPa
HZDEo9lGJPNAAYORSzGQ+ncdEetKP5duNquQgjDMdLpGZvzSmBa+snp/V/NYTLzvquPpCRLnapJw
hdB66VQmpd8eHnOkcZwJ+fvwQ3YRiAZckxW43rbVaYC2ZGn/vhJtIfzJyvG7noJXpmgaCARTNPVn
DVX5Zp0ApM/rm9dzoaRoSawYxCFGdnjWujle87O3d7FQBscUwcu5d0U7MW9r/1D7m5CIhcpM/oSU
gjq1Jmg7cUQaZfDx6TptyHx9sy4rwTO5ZSKZINE/qc5m17GRr9Q8FsFgaCI6BYBGrs8+9ShyKCvZ
hNMgJP1iV4UBrxkxO07u3ExOTwzttTVPHFpfFwxOjDxaepkEvxiDl+ncT1f3q6bMwZ65YXCawd2K
me4SEhAtcx8AE3pl/IevMHDBq7tKAavF5UB8qxqveo2QXAfKUvusLRY6zl1WmqeNcKbqSwi0tC9e
QCBkzYqmMJV6MHxhCNxtAFd4l+cdl6CSA8r4mW4tgWBM689EITETPDEYaord/6kWU7sclFp9M1hF
ALPQJcUmfd3yEysjnggmx/5m6te/u7tggZ2rKrv/eThl2IctgSDi15E/t2j6ihrsEfOKVobCq8wV
Y7EvykZiH8s/DyN4XE7WJmHnFBGYgAHjBFM5ZX2RpJwPkUmjeOlRzmxcRJwy1h6XJHGwTaP3KoEr
N0c2qRGDCzRL8i7BuWGJAZnxZ8kP6UwCCFghhjy56flSXhKp/xlb1Jl8B8cirS/ydvjCKjBDlWwh
qhijAeHZH4isxWV3a3YawS+R3FUhahkn78V8icQWbB+hGOJ9uJAqWN4p3Os4cXRkAtIOq9UqkIVB
5QSIUL3ggtRD2hsqr01tUMv2JJAQx2lZb7KZZLEfFWhXuSZE7jdrOSxNPxvy0VSZL5ptENr1zKef
UNo7ZjcgqO99a8cICGSEizWglkX+uw84zJ0VKyvgFQ6s7fqoJ8+IhiFsfpyNme922Ib8lssRahet
O2wLubQ80rqsXNvdDioxD0+Ar/YqoI17WVw2hOVOPpGqAPz86HRiEIasohs4dSIm+ugtdzXZ5J1j
+Jq+lc+JHvEDrcXflVH2gGFlPM+IKHaya8P2Tr7Sqc3xUGDr6lwQQdVS2UxRTUYA5TPJ2MqKShBZ
FnSAMAZR+4xI6JQp9s/NePj6mpBHKVwOnL3LB+3Ogo7d9OTS8lmEMSIbCToX1InVetp5sBvdht4w
gckp+PmLD7qNB1MZrKC6/QVSCUAtNhlUxisayh6Rm9/eYPVk14/+ZfLl+AMm5NPIQ9q0x+97JSCz
XRIOyze9A6pFHiPpzXqtdCm64Q1S7JvnhHzcV9qJjefNedekgadDO4d1PXO1FMWJ8CFQ62HQcmFw
pzC83x5kLgr/BUI7Ct45N/PNn0poYh2aNEze70y6gp+xnB5cEq7lWo9z0fBe3uvONPYazS9niqnR
HnjP4ovJ91OPIfKc2xJm7yxFlRWMfT9+5sh4GwNdZ+DPTP2xvUbgcNHNmcHzDcZNNWp07hrW7gPy
rl87ccUfHt2rdPvPYzznuBR+UcXl6cI+l0bOdvoNeDQWGW1V6rjFPiquF4fPM9rbhP6wvGtistbB
ViYWnqnIfiDdC3Rqs3oRRCyeWVy8wWEIUjUDu8UnuIj4Bj5cxgZXadQL7C6q/evdkbrTNToG67H5
rFYFLEAKLujhTWbFwL8HaNJ+7cN28EMRW63eVrEYyrr5NyfQfvRVJn9ph0KQWAnmqNBgNj0AUtj0
yUHNS12N4fDtKhkbYm0nia9IuSKxNIn6na40FVMMGauI8P00JpEj0rSTeDVgL3sBXtgZdzO9RM4D
aU4lL8lT8ouqGlAYpyYWDhxjKYyfobKyHtmNYtBnMUeqZvH1yRAVaRSZ5XXI9K7jbzMX4RgjHJGU
a4zeR/Zf6S8xIzBSNOGLcVq6h8E33psrHDHyVkCi/Rap8THtisxv0a9B5JIZbUVcRXSLx+LzPg4b
lWsXTGAV5Zot/c4FG24pQQQaBTfGTmTo8fhGEyQLCgpZR1Qkwip5QDD5M7DX2qiXkBR3J5Y+cagh
sLiXpX0wlhM6xFjvcwmuD+mGKbeLtuI5OWdQzPAj+tkgdzMSHgTK7zj0vCgeV3wh7ymv3FGjC6MY
qQyz8UWD1dvGR/MmFF2kUAkHe4Q8EJwQ40oeuvy3aIShJszbK1I9XefQHLv4GNzGxotucSvyjJcQ
GHX39gQSCJjt9KnkKSLVERAOFKzCXaQgnWMu11tA8EdVST+VirgTp+uHzNwC+xPdynxAruutcZWF
AO7BBW01tBuCss6ofsiwKzONCSM0R7MUPm3In+KkRezjxmT9huadVn/GtrWLLDrMTRKrB4AfoRYO
lclSveQ3U2JfcXsnuT9nWb1FiTuQYY/YLwlzdJE1T1QlSe0rm8SLQbTG89lcLzHFptOzt6+CE8MT
NwYWfxsh9lUDBT512/Rg5bcMsADjjRLRJKmgRPqsG3hwOl2o0YMYny2Y5fy13JMZidFsWis0dic0
KDxvATYmQrheM5RxfCwr2WOmzqsyun3JnCJGRaqp/EwFBxlugzwRnKVtQ6aav5FVpODjZiMbWs95
w9pEFxBJyZezs+gCfhgjab2Z/myLB3MO/dLxc2u5aT662JjtBcISUjmglKko4mby1emSenHlgctl
ZO120NP2Gb8uNyP1a3DwmjSioPiMhI3y0JdB9V7j3uVKoQCl/RzngZB8yKwt+yYtUlEpRCHDmxgW
0sTgQZ54OH9iLnHtYbiekKyYutX09MtVTOA9U/lt70XyVNLzS4Sys9+rKwhRj1kyPLI+Kj1Px4vk
k3Z1i1+wQ7D01l/Kq92kO5HGn/lMJcSHtyXNHVDfO01hF3cPSCOsRZ8C4hjmBclQWtOiHC1OdOmo
2hlsPqfARssdp/Y6q2NBSecot/+vm2LqMGWLqcrb0ujY+7dowTKigwcsfXR/MDzpsg7Q0ZkAnYdP
sf+KOJ9rgdPtxJ+aN/8agnjlvATnR/SQbvI1ZRmbNtgOj9lS2Y33XkcGU0BenwkqHy3sIDgE+Abx
5ukUDBWNuGdKtFLCcld8q0ySNb9y2fn718DFwg20xCnGkCBSQwgo+CeUZ8Hd5hXhnMr8GoS5BfiA
CzhJwvuxtetAosTwsla5Rcj4513+buCdBJFzZgde5n8v/5SdfSxp42dwqeoJqxWIrZNgS1du12Zy
9sLr/FX/ygcJr1JuCbGAPCDQL03iwZMd7w1ZOv3GgAqPHj4LVB7NtCF8pNxnOAB6rYl1OdCKoK5J
5g2xRNxmIqrhGCH3Q/fLNj5FvK7E1bQp1sfESeoHCh+QcI9jNG234OL7enrvW4lyqcllBE/2yPNA
pdKL4onH49L95z748tPCd/8HVzfUkf7uylnbygXNSBu5bZ1+7Lk/EmF1ve1+zInwz4EVYwFESpag
4jWP1btGrzPRxrEhEFZazJRUtQCa5Lu49pPLj+ZKVjAG/ZLr2cNGwUEZxjpVPAfO24HaAHTt+7g1
j+yYwMR+/cSeNx8RjVhuAw6vLNilQtLlbJEnPUyXRyWbEMoZ9yZjvkYMxhePvOKrFytbz9amHyPC
TIXpZzMgsiuoKRmAJoM58/zSdinHnisFv8sgDqFYGf9nb2lhTvmm846aL+APtKbl+myGjtfJCQ0N
aKxzRmgk+OWZ5yAWOdGnJN6qsZS8vZqpU9AmiPSlY+x0kTSShOeATFvoiDi063a0INrHcDWfQvtZ
zHa+N3gWmuyDiFL0C2vN+bTDvjbBPZSL/UwQnpLaWg3lIZhNWtE5+SmcYWPlCdnVHnzDDzVdQ56C
Vw4T0ZvVkbMNmXAHy8/okW/68PnXkiUU6Z8Z6FS4b0oDN2Jjymm18JEH2mWM+LyzVb8HRm/F7JaX
XcYTtkdHC2DaFuMzEHv5DOl+EDBbKO1fPhLH8k4JFWnv963d7u7kKACzkF65zHkIndYMH+04kKJE
t8Y57n30e9PYhGblxe787tc7otAdlh9zVB5eqcULQXKQ+1ZSgYt0+MxPnuzVY6JJ3eAEBfUY/CZ2
IOH+g+QR/6hR7FHnU1XlnwgW/3LxOg+ZkMsatxuGzUWNg8v8F2z+t+j3H8pV2nF6B8srEJE6jZey
5u7PqrK3ahZlSgUVzjGyr+IH3NcrmxZN4aYw+2BYTQ6/Lyn+am54a7xxgUo4dVkm5Z76nxSEiSoG
Bt1Na98BopB/TdhnoXCw/xbrdGts5d/GvsnbiDnlL0fQQjx8CIRUrQZiyDLyU5dkuZ4ajGDThLfi
uKlbpWEYNve56UFobf7VdbV71cYpa6ll3yfa72VqZNhCLqJ7XM6G4bhJtz90YpkcgF810NtJM17X
YSDKjZSBcpVHh7Y0DTXw4BloNbZWTWwTwclFR3hErRan81L5eTk+3tLNum95b6cOkP5A+LK0Sql2
S0Y2G3w6PQtg2TZuRtkMJonPyA1XkQoiRdvQB/8DyEDyFckRBPs9hDl3iKp1jnDwET8G8ydWKu60
KwECtTZ+KXc0xGGH9DTiJVIhZBzXLRFLI9cQlIz8LujU8+LEliy7By1W8ir3AsIkLM8WclvhVIP7
mwgwKTK9sTdCdqr6M3R60FdvMmU6v1UAwGHVNX869ezzdbIMg63vMjIczGNe718Qddt1NtHiL8Ok
PjjTcHM0Pm1WX076d83n3kweJuH9BU36EJ4a9zqly0R1pRCsEV0+HUKNzNWDNUNHOrIE3/ED6OC5
IsJY+FCenEUy0LBEJkjXxSILvhfVXi/jrw2zGbAamKoy6hnZgXAlYKyHw9U29cuA6AoXugILIvUP
16wGcCU0uF7hCIptw0uJ6vENaftLWfjH1sNILHhDGDsXG839h50VcD/V4dQXVqCUoxq7MS0RRH+n
sf8DCh4g+XtJe9uJkfhoYN4zfRE6kLtIHQhR4I/IZUiV7WGFE6uzBC8lbsiO3KqmIWCt4a48BW+H
FwFfN5BxhqfANktaaGKlJSBvXZ4zyK/k6Cf27Sdhxn+3UKde+Xnw+yMpXYQQe8mJ2OAZi8BNFLd5
1n+CV54M4sphtQgjcrG1EFZd9Q6MxukqgfVWi4kn8mthwEelwkS5JmqicjRR2swnDFs2SJlMJgE5
7g8WMZ1RwdJKUfVC6TZbi3sA1p9mVGCIpaLxY3rU5B7p++kIekPrRL/Pml11dKsQylnsY3/qsVH5
yEK957oxUSw20GXAgKCQg4sqs8Drlvtr3zLNT9cyiUvTSwq7Pp+r50qnY7xeq5lPoqqnfczX+osR
NLktEuNnYuPXrt47VycdOWbEYtTlyTwVRt6xillfjGF3FRR7M+4/Q12VH97EfZ7vu4X88Qx/PeB4
D3lrhiSUKwsfiQbWhuh0vxPRGwy+QztyR8fpHZkbcm6+jVwd+7M7jsWULajmGTQW7bbIh4efpwgM
bSZhQPWk57MkwsmlS8SFpq+KwdOyK7nkovK0LqeGognmr0Duj4vN3MQID4xp4vRhS3IEEn9P4CKw
QLKEABAGrrU0iYNALru+afKg/nHJ4lClQcRyabXWkUYuaJnvKhRxNVzindPBPeZnqnQxlgAyj3sP
If+4aLjdWf44oVPV4B72YJ3CtrKgdP/Bdm8NTsJ15y12/beleCtMxbS0EDyBlGi2UulcWs6FUyfj
HxNNY0LkjMvtdshju0jK3MUyWAMxjCLziKfEgWWzVjM/VdSeFZ9bcWTEJKeNRwc6NKzwy5+3C7l2
hOA8tET2I+rIZ3yMx8kI8nzVqv3BYyS7CpwDQkU7b33J35cs9iVTBs3lwl5p+Oc1BUKyuL1pLLba
IM3jsUxQ7Dn6BDsCsdI8ulxqAUX2d+pW3UN19e8/Mb6YOD89EKvpKTtk5IzSJWQFuh0leB3xhOkH
YGvJC/cpkt0lB1OMZnVCmRlv08fqjVgiwLbQ2OHmnao8xO/uU/OyEFk5lSMOrrm3+SFfcLpvJ9Tg
0vYziAw1d0xgMNC197hQ6KsxXPoz5X20x9ANje70Xzu5VpWVtzzVS/RcWiwpVKmYSWql4xkVoe3C
QjsiND3Q2VUUqiSyNMCA3lvevU7ZBo9d19w8wbnNn3IGNd8Ox0Ryx8+kaJP3zR/fc/g9Lq/+wYSP
oPxrgdtDTfaRZj12T8XgEFtglKE+sCAIbMIHPfHZjAxif0BwJneOLypndQ+9kMt2EoxPWFtO8NoP
B2/epjnwTI3TNDXRPcBbCBI8wNAhtbUtjfxfjozTJTyFtzuAb2frrzVkGkQKdMJ5Jl46rFpGZ0qg
h0qhAZ68lbr7r9nKWHXTpTFP7Vdz3tej3cYBCnsOjGplrq5kF+W/lQFVcHGPyZHbqPHruhBS5MWD
SBESaIe4r3P6UOBq7ADeNUq0UhVWy34vbSrxLcpoxAPmv0ne9jvVt9iCSteq3B89ZUeRSOcXoTeF
nsufmE9j2Sl05fJ/ck5pqFDDi9a8/8JWsX81EXU/VHX0lieAQfBXFn5fwcqYlspaVz062iotl+qt
xiI1rLTimb/EQUWy8bo2S8FlprqKOLu0oI9jjazmD45YE6m12wWweGLW8pj8ib5eom2LCAtgcQaE
pNdoSNz8IwqKENVS5gK8VhN1iW4cQQAlzL6ldJ3bmCRpGMWdXYfJNhXX1FPzDGXCrmuxOTyDREfF
sX/GtuBBBioEBTwkB1gWyjZLiLHrp8+aD+8dVlsY2rKE2V3M7aOEYrkIIsTHdEA49IgT9DpRzmvP
E2fpkhq4/0fd7aAKWQHFy2m5cYPWUJCcy9nMjw53Ez1oLBfxT20/e+2yt0JKlD/wt+249IfgpnYq
2P/vz0SenvlEXH6gBsN6ssrZpEstW3GSaEJKf3a4Vg2sK+Wp+F8acS0eaKT+UkqsLv5CFhhSnrAT
wyRG7H+01onANgyRhCdcS95YQCFygzDGzpHkE4BpLN1VluJSf8lHS98XkPDgDK4jW+WDVadOWQ1p
sEnX4xY515hPgovy0dyjFzc1nAXD+q/bxhnnlHU/dMso7VQ0idzijuRFrsKtEqFrcsxGBoFPksbt
YDSZ0/rNkr1OUiRz5Frjxi+TL8dUPJ291LoLG6VMC3ibp1wEnK0X1XID12HEC7tzD7cesWYKpty1
T370STkqnPS0QkU++RRzODsMhbsX7XLDbRb87PqkHgExRhHngmUFwZrrZpk3BtN9tTXU/q/OMghP
YfkERb/Fq26QqB8NDf+wrdKRSAyuhi0+MqqgvV8xYnvBB96ntVXRMExSMnv5neNdH1j0TIEvreG2
BCfduYwjmFuQEp4EG9V+WMB10PfJmQadVKhUPZlFbil35HL+CLJh6/wzSdw9SIVulyGFdrklqd34
pvxww3W8wYVSYq38iFxgk3y8i6ukSJcksFFcV6C0uEjfKn4dcQN9EC3k9W3Or6T60j7DL8S/aVS/
m7BYkEMP6eq9n/uMksIUmQQXS7UloQIM/C4ONO8JTKzeqJj5g8oj60u36IK7D1qMxNrB7Gfj3vMf
WS4qcUxe6kaU9mx5Uy2Eq7Z/nVtca/Iy10OqIpylTvlCAUeYgDXKkY7PYrf2iFxgVAIP0xyttzLS
L7ZkTeHC4bede2IB56jeHUiNDxHtHl7rwJGLnYg4Zs74uxlMNiqDdIjs5EX5ROjIw17r+dRSB2hc
9EbgILn12OoOOwFnaq8X5pktyjXNbp9Ew8MaffsxB92INYQGYj8XSlgvajkqwfW7SgSgT5yGE7le
2Xf97ThVMMRzmj4rWQnw3wkq4amJiy4ilbOgL9qGW7HdF6vQVE2DlVqMU0l9JLkxpKeNcj967Va7
e79qgE2nlJphjbc21fpMENHE6gVdxh6lzkvohAL+yJxqSwtu0Z2AqopojhZWRlBpDX3fcEpDG1sM
6HLjqzrikMDlpae6zMU5h/nkXgstPM45dfKjDJCgybrq9iDHW9QbMAAPbiDpZiYdsVPz2rjeJDSL
lH4FgYhU3WzG6SEym1wtPv755A0FaD+UoK8+eiiNb+k0Znopis2A6oi0PQAd7G7dtiUVAeKuCglT
2kfT9dMtrYFqTZUBc6ZMJu6AN2pKekTzsVtz5MjIfHDgmM3iAYgO5Vfvecjs6fTnNQ642Fr5Yqs9
cU/mKm/MlHoQ6xKoKreYXaJORTzDinlj8Wry001pgALycBbfJ2enKBJAbZdYaFWwpnSKPDuI+u3z
r1RgXGsoMWff3jgQH6pni60+jZdl1wLaQTT+pGlYkWI4arAaL+9gb+sNS3Xun65mN30fxgPs5i8T
5ymIZ8WHbjI82sNSJgjYDiIuTfFLfWVduP/p6hcJYFsOx088BBcR3WWhNPKVPjs0RyCyhTG3/h9O
svy4aHTHJfS+P+RMz6PPiKXEEu3BeZXPv6yttSUR7BJaNOCip9b4VII4A0toizNBx2EALNf30UbF
fSRXS8DVveNEs66Q+jj/wZ6H6yqh8hrH9s7+3Wk1PU0KVeAZRX56rLEJcw1AVkqoLfmBYTitJ/f+
EgJnSUFIY3YcKIoz2CRXy+36rqiv8TIX/EngFg5UraoEYuOQcnePPjXOJMG69fj088Ll1QfoT0Gv
vgh8nSA1i29XUqsEdWRAvo9SLhx0+kzC2eE5IE8mJFRxH0kf1fXz8g2Oi1HRoQhbdx2Il92NrdpO
yYFwstMVmTxU2cSiZ9SHcQiYMbR1wHdqZcUb80PCtbJc0GoSLAyQCCts5uFhsmF8HlGnaf7tImEl
DNlAOQYI5aS2y6iqBaCi6FFi8/Xjn0sFb3micFALZHVE/rWD9dBpcTMCjK8tUYO/+8S55o4MxMNc
VUJJsOs7LCh3Rha5Dd7zxPatGou4q8fYTo87sJDHXZ9G4lJEl9uj++n2EjL9GGrKLXT9XCrqQW4+
6YMF97xw3aNLEwjU6rnHeXW7p+ERBuw0+5GUAOH54BF2jYyXqJf/fpIRPHNEv10NUsBq9IcHiSWI
cTgdqoJXN3c1zGuQh/2RDMF3zRibrDXBcUa3BJ0DEuHgrkxuI0uuOQRtRjBK7IPvSYMfy67wfKpP
MjXLKtAoJGWVVU6ySwJdkfVjfC5Ud/lYqWfeNlh4xR1Pi1057+IHEx4iUvattF5/I9//CH3YLzon
64CkVsxI3ludmEIgRtzB6Tsz5F84+mMkrHYGN75F5hnEbTwmsXQk32YtD9iOJUeUNoT61pUzNrCE
QZPzO18ptnlZWNGdm/QdLFcQpeFIgTcD+Rtdaz2urGTgaDz2mzHhgXYPmrLi6mvJR5N6qMUvr97q
Lzlun9uOnvQuR5KuDNQ+N6JXEDUSw6bAqBmDlD12NlAYZVv6opFTZWPSU2XH/rIhMEr0CWyqW1ND
vzXumk4c76ZSzBT2txZlG35QbW5vKgeS9TXEq7+5wHqpmWJo5UsZFFOddy1eiE36bZT7F17hm7Sp
ODH9fFlyA+spA0EFEFJRNuAhB1PXjVDfTrdYEkUqs6im99SzxFrpOk+99mniw9SXVLrw1BygTQWN
02AzRHiDICb5Fnjaq7lpOpMQ/d3Pn2PvjzMsR3y888N+8tek/fvwQWTttQkF7wgI38uh0vO2N84N
lqR0sQt9i/h7BReNUPzQz66/BX4uV9J3osxrSJbqAwYMf37eL80syxFk3Hk0VaGyk1rtbjyQTOuS
ssdFy7hSI11dN1sB1MVp+Wkob8bMNWh+Sw59Q2ON0jxNBs5sS6bp7zkO0aCiSVQs4HInlhs8LI06
H9vJSy44dKvrO9zMhHLLMz3TIaADjOKeVgaiGkaJ8SVOerelcnRfEoHyZAgzeIKKaVV/+GOoiw7p
P8ukJ3GDflJg+gsdhXl6c92N97Q4LRQoVdDxzy6hHt89/cIfXROwWMY0GN/cWZDJa1AeMKLlkScQ
vykp/CaveXoIdDBWDJUD6+0HdQfk9A4DhvrSqV7v25o6oGtb9z3SYsey9jf+KEBrxKBspN0w7Bnp
yut/Afst/qvbHe19syvdFtrynbJqW1UrVI9pxHkkYgHoKlLxvnrSUpzi8vkO7YCwkEJgHVZ+u888
B++9aOLTPf6iJ68GjF4rFnVRbLFIIGt43vmN3zOW6PeoQmT+7hbDtoUoM7TBxlMm2o2O3DSdT12t
taWtLMM/mc6boQOVbIJq+C7GJL3gaVFt9UzxTGr6V+nEOMXwY1uxmB7hX/1SPncDKOIZQHAylsRs
pH8GZDWxeh8MABlARQhAddg5px4OwUDuN/Ttm5CN2HynH08FeDDpjOUmi/Rt6pwrn41KyFyvUoOU
rVgZNbu2BC+SBrge9o5EloEw6s5U37nk61dtDmsV/JPcBanixAGkpYu0N8K1/bSpn1SoZFJRE1Ku
VO0EUKL4at4vjF0ldvYG3+XteQld12MUDo5BJNRt75jxHZKEBS3leoooNb2TRDVbcKOLoIvy+Nls
I7K7/QFy3/3Q97bEWp5yXzCjf/kOQ/vzT0tIWFSSWBragSmfN8akG6YGCNjOecMpifKdaByYPKpJ
buJLTYjTa+9oNnC06zVh7stYPQrXX4/6nADJJh9gDPVPzD5gwJaEFOf4XdzKVfRlyLr5/o34bRBz
kjlqXd4yod+GGFTnIjKEpAZ/n/kBVChSVCBxjbNXukFre82MmOz+VZn2/LmYrBK4Lr2j+OkbhiLf
QUR9uy8+k+UPlPAfUj8nn+8/MuRc38bRRj4hW8Uw5yPn/z6eyts84WyDOkMQaoszgkZ46Oxyzlt4
Cu8zPv3mkx/dzLBJcz/Y9QkMwHRmq4Igghrkc/T3sNBvEtKqrxkEdo7jcQh3PH2YPApUbMs4djoN
BhE5lseDvtAQ1VxKqAnv+Z6/CyEvbvALcV3GrAKkvBAXfD5CBg9mSkayw7urKVZtlEYhLBtKTzIZ
bJ1XpbrsjZ1HjHv9JWohUfOsrMRKXvW19susTULQl+Szeyqz+SVlIHDaYj+P19Q0GJs6W2nfVfT7
HpSgOeCuibwchS+lkjUw5gU/lMcyXPFdBnwGBez0vKMxIlxHB0FxoIDMr22uop9QwNU9Fn6K+ehP
YoJj1u+OV2xo5WvW9sGDVDJ/I/OqUUxaq19l9Ea0cdBjtjRQrygAjNRGFmWEbnImy72R6rVRuqI3
/xeSmQH0TqABEvHESA1dNsFmrghb0susS8hPK3wkuLyoI8SvFZMN7FqhvRs+njidDjFmh6WK7U3Z
wEb8Dg10S8U9d+5vxvmQPfI36GWq4C1lkaZwvabzwESbLFbajMKlCFXYphNinNSGhFkpO+nim7j+
fHWIcHBZlLGtfe8/fjIKeT8pAKZ9MpqXR+8FXWSInWVaiqJKVaXoLVGyRIIQddxsxRgK4tssLvOp
v1+TnRQT7zPNFx8cljrCT6ykUEM0Y3Pr0uA0QAZ/lHsZ/TwvKdUuY3302hT7tLkJFLfk1dpr0uDr
hnkRXyGqUeu7Z7GzDurFcCvOHtqslvoohhVo1NCe+L1hfkeXM6yZeePZn0iN0/sdmQEE1DpQf2yO
cvm/SV6WLqGB/iRcNvV8OZO/+KpIUAFP3O026Ut50Mw0mNct9xhcYv9LdrWIqIgS0MqGSB2E4ntw
etg/ErCHbeiH8lHJn+zN5BVAsGsGVrgtm0xtmF4GYOfGVOP/21ETwdZJvRPo7Bl0UiSG5uEN6Yvy
qyw2jK3A7jRZT5mvu2mi58chE2/w3pDEwbbfL8Bi/ZFcXdX5I9Re/1h9UnOyjdBnImQkBSro7CfO
uj/FKqpix4jNEvLTi2sf5sLdubHGAT6SQ/xNdxOjmlCPDW6YmTHHyGKkIIWl5Sn5DVoG3x6JmgKW
UUqq+Eb1oll0IdBIZkdGnkso+AgfMuTMDhHK8YYcJbPnFz6O6SRD5jgdHwE929o2paS8srOBDqjq
uHvtf3duSQGo3hNXeO9BAh5Xh5dugsN0US2Uoed967rj1XFT6vHV/4c7tj16mFdCswHdsTG4OxIq
K0ob+xikkPZspEUei+dIkLzLPiVC0Osz+8FDSBBpj9c9L43Ck/dONLmS4uJHcrTzkS8qdnmv9Zt/
aYYmnLxGOjqyL7+S9oN71BUylPwBKhPKceFGulu7Kg4f9q0uMl1tNbb2O3LSI3i9TtO1wnCzQttH
SIXUbd4diGM2at+9i0yEGE1JUhluTr3VXa+eSnrU2AGdiUu/uZcVhblhhp8922W2N1SMCKOf1+I+
Ok5CyFi6ZC6r84y2U9qQwjyj2fLM+EckAitFqKy06DTpHzm3fPpNzAFz3M1SeZCErMzImQewqvXT
TKZZ5lMiy13A4DwHE8dPTB26L1r1N+xVqr7RqKJEWC8AuvcZoZfZUbwsAX95GTvKeAXLANkUowrt
GDScW73zHjqYXfajdBrs3hnUzyEsg+lzkUfpAwTtFuX7bJEdkNze+P04o0TJa3yrDa22sajJFwQf
HRBIxX46j8cOghtL2P2eM/OCf8yfv3BeVRyGc3Y1hsfXyFrAjTjpajc6tBIwCOg8VarPQ0/W3eVk
Q5m9lRyCZVHf7zIcazXlnlMYJHsLUSJmFed2xieVDbwEzId6rFBp8vfRS7Lttp3WuvQBOWWEGgFM
terwNerNLwvVtAuA+Lb4foknI7cq+IxgdfESXYZZQvqhrtpVcLp/JxxgEVQdHWh4MJwK4O281M6y
kM/QS2C7jHDAjNPC3g8KVxMh5WPZDalvbFs18N0Jj++h3Bbn+VEEGlGUNvIfHHrHfAL0zwnHR2u9
sn/bnTwoYAGy5kyxqg2EojFcKl+WXIJ2JgfSzP4neGoE13qoVNzdrrNA9uBxUZr9Z70if/8djtxI
AZRU+eY1HL4f2vY3fxXf01uESsR0/iwyd16WBgfU7aF2AUfanNBa2bjByMUHHCxrDatvVgWS+Ytu
GbLufeNtcdGbJabDpTJiKyYYeO1Zc3Mk/ZCqgXE2UfzhjcSP+YCQz/XR2/GBWd7bL6Zpg8/GV+HT
sawMY9wS9NRN1C5XJx9JTm2p3kZOb0mFAr3DFY9ecGpseuqcSygtyFkXQ40/UDpBFnRrbEGwjeil
cI16Z/p46PxUGruLFPh1K5/QU5TamQnUzOo79veYT3TweGpva6kJiM7M6Dte3pdiTUbNjPoRqFaD
sC8aVjopd9aUGlNKW/SXoL2tpjIeofEkuw6VX2kKV5JdFpQFmkMRZN39N6qAUo7BfCgIA6AP2KKz
AcHXGLQSPpE+L4CnaB27zKpqFwIBPmMrnNodML1ZkcjKj7gvJKBBCf3lguv4SoF4ziQLC+6TSaU8
9SCzvhFWmQFt3E1kCRI/1Plr5QdlqxPnwck1RedpveNVQK8k4HhvUOcspmsOROdSMmIvFMEiHl/m
0v5eu7xOmmVSGKdLFyysMrKPE4Ygez9KZjCM+FYCJGCE92f71iOW+qgZs0ZedN8De6xNbT07MSeI
J4k3HmDaqPR9OFdBzSJHXajVl0qkqN2mCHrWc1Kffkm3iUaPSJT2AiAlG3EjsCmRIreGPhYYfjqC
pbQWfA6v8a0FiUrxfeQ+bZEx5KuAPRpT97XuLkQWATpo4IKicID8Y3ID10q87wp7M/Y0HYVV1HdI
eUm8dQcngvk/rtFT9xws3xtqKiHc1gB2HhhQ7yYQM0YzEmIlQDyrRsecr8SeUFHmr0QdqWlU06Ff
oVvsO3D9CtM+PQHyoAJFOT9sLcGqkyeTPwShad20p6Hd9DIlqVrudBjpJWxs+PhcJ5um0BUQpgrd
JkGreg79UEIGiIZg//MfyG+zHYSro1mPTZY5fQgvwTgG3fhOch+DTqUK3QEq4ruJJNyumTnB/+MR
I5KZVeAFNjCKMKoyqtmCr9SRgbPaDts6WsWLcWblqMTrxxVvsqWSSM4T2er63Q4rA4O6KU0ZETXd
EC/aR7jB6Mhd3AK+L6vIS1rqbNCu1DjSi+SCZ3w42SPdwe/E1xTCgwwQVPpYF+ndw42K3ayBKP4i
vNta/mplKcPuCH3nzC/1zXa2uxInh68B9XBy7xkwR0vO9RMXtV0caHwEpq/yudIcwbnJC9QatLPU
R6scXGTtKrvZ1BNPdKgdljE9B6/nNV2IxEfuh1tAtqJpDyk2rqAupviD0OKq+oQDG6qykxaeUmoK
BaB6LKNIL67mGotFK3U1ryWHa0YkUimtwLU322iNV7PYf1p0LZam/S8Q5O6DgUvS9+O1sVbUAedG
3Vhr+T3eVFFi9GXFnZbnRkxwc4dfDYTtMdvS03i26f6zlSoLvJwKigd3NHjRTDIX1sdEhF+imBcy
+VqaF6ebaoFCn4cUF6qmnAU6UW8j+fO1Jiw0SvfJ6emQXh+x6Rb0ys6f6d259SR/A6wrgGAYo3IW
OEMY7MNdQwNy3itpNdHUhEKLJQXd7O4BqlwzRwIVYMAW5R9jy0W4jXsAjGyTOyybYptUifThefq9
oRCi55blX70dDt0WxPetuqz++JXqSsshCqnsL6jukRX6NbTvXdXiwr8IvfuAC+BukLpm5iQ0m0tD
2KLS3JuKDehFjujUY6sKkhjdhVNL81gIJeonaipQQOip1cJqWhPmhtRCsp4qj0lHXN8wY4SAy7pP
bMIhjik1ILFIk/3H1y2ng+Q73/i50SG654ggFJDmXg7TBjNsC1cUXGmaDIqkPoQfYjM3ViUduJeN
Cm77bRRDxz4j6jBQIQtlyYH7BWlzUHCYf7vzIlOPlnyzO3wQ8zJ4DuWC+HBBCHjNzNaz+cGcdLSg
S9df7O2yCsD3kXRoTWlOpFx2oD3WIF10k5VH5ST4lrKLYoxRAOlIdds4Kt+JK0BVx+nyCueHgSz3
50cliUZMQXddPvLnSu2SOs10Q6osaMK8wn+hKcDGoi5p7UvodiH6SiL4DiFq004rPB16jmiuGXsQ
xeCneoXHPC9K3ZuqOg73ylkJgg3ZvM0DHIQ8dzaAHabTyMKi1dcul6IAB25PuL+lVIUcHo7OhOqm
euMnKOMxEl5ZBHwVNTKgnhkIpZfdBUBdhLxNy2ZCIoWzfA8GGTL9phOHMDjbrvvcpVV9tRLuh165
PPKS4wi0OevlllvAB686WQAA395pJov6zZPoTPUD97QdYOkYbuI3J23vRgm6GhzVu+awjExf/bdG
RmPb4N2V5coVqmUk5V9iTopwbxwZ8FxLzF6qJ67DFRaH4XQfknT9GIyBa+QNgG3zbHgt5oLvqdsa
707Z065pZW50Kfw3anNTZUiUZW+W0VANhozjzWqSU2FTm4h4Pb6JPmkzewtYyPDSV7byGx4lCSna
14X2vzz40jI3v8+uDDFS1T7L3X16N4j3A/dhaEXuYLP9n4n53VO4FVq/PMgZwxPNR0pIswkSbbNO
F88KuVC6bNk6XNC6XcXXrOIqOeeLPQVaTy9OnaGLivIfgWIpk1v89ElbuzSdfkpi7Y44QnZO1af0
Ie6Aljxkb1JRQ35ViwWYuq362D+57k3hYWpxOnEN/138i2rh1FjtU8pw3UiMpNglUtHi86bSg36n
UYAyi/xlX2BDrGvvjFfmLopGiCx0NohY7XLBKjdkg1P8nhnCxyOjWjY1pFyjbbyMjYSSgoVzN8qq
fqGgLksUGqmIbiAUxcdc484ZJmu6mte2FMz7jBt7k2GSSC8iBGH2lg5pQeNmxtF3e7LWytiJbD60
d1vBOE4SHMjxt0MPnmCPlXr2qA7pDeyuI8qIqiVJtQZjFeSisiR97mJ/AEaq5r4Pv5XN6dQ5hxLS
mgQ7sFkQpYpnZX9buaYjcVXyRG0gSgxKHAqogT6bv/tmvBWmOBw/ox8GF8O2UCl/E+zglVP3GaUb
EzNKeSY/FbQT1L6oUtBslJayYFjLa8WoSBWzpiVEBTfxbagCZC1LFbqigP3XE+ohkN2hphyCgY9n
ICfdts1jU1llLIah2Rb+JB/1T4nJKfezaRsyTXnxLwNr036WUkeoTBI5jUyz9Hmd4dZXVsOaIw7E
BW6Xjfpy9LXQ5Xpz/MDHAyPe+c+G3mR7E0Uknnrnw226rYUePhx3Te8gUrDzoFc45AGOtQfOlHpF
YTN2fJyfAzF0sjLq++4GHP5aWdxfaptppeToKfcAsdEtJZAtjS6mW3QuvJv/+Ta8Usr7M1JbOxHc
cCSbg/cNvtZ5zN4ua9iWYhBqEE+bj7KgkuBi8UQpJ2jSPZU0dUPu6ZQRpWgK9bqTFkU4UIQHRqvJ
elrr5zSKywvb64+kHpaX7gTzTE5LJLkQ0VhF25p/1ne3ggOBadoCBVQK5BTxRehCZN0nQoAFEAqu
A8No+gpFnaucrxWpJvOgKB2ctXIsz/7OLyzw1rZNsPr1Cxti8mOcX4U4Ovp+5AfQkH8p7tgiuW7u
PnjEhKXa5JYnWKkpurqStustRZ+35dixxz8TekbgiwCxUKKhZo1GCDBrurxNcn0xEVqSJTfyWMZy
tgziKUCxyEJQSYZlfLBdh7+P9NaOFCaaJXGzzbKNTKDjvUwjqZ0rtMA0tTdLcXlMX/0cuXvgP7h4
EC/DVnb5wxogFmqEeWpWZm2/Bk3MwX3Q9lrbkgLYHh7yQDU8ChsLdYcsKEMgAEB7YIV/yqYcnajt
/ayLZMzPtp+lfRt0ZhxUXCTBdS51e+zbD08Zumf+dFrLBgGF59FZiXV+8ogG1+01Cv1BQFCCUxbQ
cFu+RW+RSwozVIZTS7OE980B33ltk53EFgkUXa8cDmsP6dKRwcKjzljaDrCuPU2lbnKkQt+ggbWc
cD0d66P7s4EmB6N4TSEsqkODlpYZ+hazEjatDXSPuWvrSt11HA1L43SKsEzmXUqZHbMht0NwQ5v3
rJQidvG5ZWfnl6GeheH1oLIGmeXh3yRdbg5jYLyiGOaQuf9OcA/ex2jTNgR1/TFf16ju6Q7hhMPy
Mm31P2uGaBOkLH/00KtIgiu0bjKyYljVfv9KM6hW3EHHN7L5UYodZ8CUsEnOt3TXREDshXsZdQsj
1LQW0Z/EvLTKz08/rV9u+ORoNJnq0Kxv0gOfpRQEj5cxPR+UWipHGqohatK5BjaZvDOcY/ngn2AI
b9miaqGkVGXRfJ80udo/Lwbf2+c8cItnUtIRdofn/VJukmE+Xemodk8yyCAFy3FdLwqmkMZ3oVn5
ctF4udnPm0VEMsDHiTWcDgydflGuuAjny8rLhEJFGSh32PZpjSepbRYH2oay/s+sIHfImEa3VfJS
oAH9DHxZ2eD6SC8LzocPap1llFIbBMJTphQoOmsR2zVYIOzLoMsZxuP6UDXbDjNvpPWqSS5dEzz5
vl0GNb0bSZEghA7wuB/8XFO0OULHu0kG3wwYAFzCfI5ri8EBdMWt/cBGKW96/9QCxKfpk/ta08kU
tcnVlZBPQlb7AJRS4iiB3we0FxCPbCPeZ73/LjU5QQbzPFw5836O0ibI9GUwVdtHo0F93qc+wb51
YPQMenzhr7Xuiq/Ob66bXIq+yoOHOypbwg42zrtXOyfgHWcuSNslf4hneoxUg5JDVKVs03R/Ycyg
5z0YDLfz6B1ZBaSa7Kwd4P2R6vn0Nl7/82765GYDu1LH66ncb6Q27YCnzUlBxtLuc4utBkw5cU/T
tOvLw6Ef+9tl4s4T8oqrXwgPxA80UlvG4OAxd1wqutvmYtAkQFwZWJWfgaWIQv74rMAbdbxtLchd
4EJ4NRcX9ivVJY2AvHC9r7IwoL8QdDehdU1NEvUsNgtWQqEtMwHy6AdBOF9LLqSsTjlLfVHlwIUe
UFOLPiFG4x//WZGG9K3pJZKfDuyJs8AKZO9T6qRzhfSWykI1xphSnUM19WvdgV/Cb1HfRA8kT0ZF
9xpyrqaOVNzUtTU497JfQj5VnPy04QBOJsafwZb82xpgt0rb8GOIxrI6AbSv/x4BKOrRl9y7O5/Q
ni7ntTLBbnPz+ZjQzidvlfc3pKwgV/nBZLfqKNok48GA2/Jctfwx/Adi8Hrz92d93ERVDCEL+/Ay
pF4G+6pDVGe4N0gVw2zyzybUKBDNi79tMAtc0GUrlU8fECBNC9Qc93GDtN1qJTCiSWyc2tz4lT4U
6m85BbGa6z5uIHVx9mworWbpX+05WmcNmvfhcEUCUn0Z6RvuDAOaetTi96Pb+73Eai/RU0ETL1sH
H/GaRq0BfY2fY4EHpxiov2ReEan1o+BpSQSrW3odrBmYaE2GmfpRC/T/onFRhYn6sddbmbZo2p4w
+DCOFPioWN1ut2XWGd8BZwPri91lfVOmCrY85AmvQ8nUAnMHkiS1q/FNEUyE7uqL7Amhlyzpbezo
Qfh3RZqWOlruf36Vs8qyCEzRS9RkpAGwVCXVFyjVWK7jmWNbYVj7Ps9TdVXHU6auZ3RHh/p6debx
kr3fhinqppMkbqcVdqHrj/KMxORYWW5N0fQ+bPmi0HvdDsrMehC73Yty9rkgQ/yDFPM2MDVIlHYx
dIOhELGVgWgBbrpiq9NyKiXkaW5rxQhQG1GYQL/BmjL+F5ofM6OFh2/47rmsnVf2mSCULu//teb6
vXcB840c+uwYfuBMy+lFFNycEt+dasgg6CV3Pbu6KiW3fnD7B/uVTqRfcxLX243AZk1tO+tf1d0E
873TgnCHDxnI0bUFz/1JYN8DsreDFITSnzWyXwzrx1ldDmwjViNp5GrwXk7Nw1YhdHLyawy4Ab5O
56oaqurTAzfgegkih9WuHq5H/WoqjoeBhuCAB+7JijG38l5G9lJ0/zmR8iyUoCiP1GiRVxuhQGjY
9SyXR0YErltrdxFQsbWN4hByyUR4JIesdKO2ilUy1tJlXdB25g1qqI5VnpaI1NDGHuXTm3Y1WDQa
gTrURRRhY54ExVyqtespYPpFJjQww6wQc8nBcPvI83RKq+rEBwzLNEG15BBfwGnBWb3wJsHaT0Ui
dRNrqGA1pE5K9uhuW8eLdeWARNJ7mpyf7uLHlE3KmE3NtHhhMA4PStc6o+iuuEgj6r+9Xw+0+ugF
fc4LYJgdi8QUX0PT8y7zvw/Rl9M6Yxw1g612vbviq9r72rhtttvYzSwYhPXX0VgfHvGX8zUql6pC
pwzWaewm+oMnGCB3IPmmZ9MbcB6DHbndvWKOvLgCTEbUG5Qs0C0N3W/HnWMrVxNxECBiXJzARK8C
wMOAITojtsVyqbXNeN97EYWuBY6S1PH3caHlu+XYKXIQbP+So5q1PhuScjxYtkNB4Fy6XHQbkxcF
mMezFvaJixagOYOrm/P68sCvUeXlsraZR73ssCzXTjQmCwu/eQVlgqPdvfWqv9AxTSSQ9QBo67nJ
wY7yN6T0IgwJRTPISKL1iviILzMscohpU7IzdGcTEiHrAtMU+gHd/EE9Vv7XmlJKqx5afd+EZRsU
iu8hX9WbfSNTEKouY3Zk//h9Bl7jkwV3OFqwR4cVBqQrsANIx5KVvGD7fSUKomTB/47XAuDjdK0w
xeEojsbUbX/dde4VlZGL4qU1M/1POG7UwK7ho8rUXmi24e74/xMon5JQsNACv0e+3QdMrUzrXbdw
133a0AtMq1pIJFG7D2dGeTNRKQ9h/7OZhwmTDLWpwysN3fOMlgAtO0If5tGpCnFWC0mxJ9dyFLtB
bndGdPC9BDvPIFbQecfAAFCK9mT+9e1+JLAWDXhYyqk6rbMfKlCaZIpY94w95MER9RAilUqdAFWb
Ghnhb6J26vmYz32ykwuO+d/dhwKw4MtBx7uKiOxHos6aC5Wz4AmeyqHxc82qnZu5HRal1SRJ0NLK
xur797ROG2mggp7B8nd33uRYaABOQh4eiUE16J4g5VqH5jD7fqvdfaca+I+Xy/pqOsiVb5KLnkMH
xTjk+imyGnyz9TD/7bP/EjI5K3grURkwKTbTMThaGZ44z77eaMBbY0qLAySai0Et7Aoa2MUdNOSx
VGxQHxyjKxjoGrxf490DoiHUg3W8dNxNodyFjh99oZOIvFZLMllTpszzh/pXywt3P1AQAVR/aQPg
+ssIkQXpjyYENM8jcN9pqPKPNJPjYbGkHvijmskTd36tfRHeAff91c7B6tX3LQ+MuPCVNEcopMy6
llX10dz3WPnHsbTkhi6phYtkW7WVtnIK/DiHj5pNyRWojGGrgjKfhPuCZtg2w7GlPjsWol4i7mxx
H5PpAxUzPEXANXPCYesUdjFPB/a/gCEBZzf3VeXz/oTvBDhvfD0QWhHsjZ7z6YWKnB2SMAUZ2HxY
gn7M/yCP+VAxrFFPxOvykyWuL93A7mIKszFbCCJp3mHkXs5BFa87BkuPjdmPKo+ieLD9iWfYF6uh
2ndROf6IVVYVLWEvEDouLjy1HYFH9iX6V96l2dH+t65lPVQOVf0+DkqwNMe7/zKpWpWkHjoisliU
L1KcBDxGfd39mQQr08INBX3JS/torSK3YjXakgxp/5SPpVVEUjSSikMYFyoQjM+zIkrnNRvP1zDs
TBVuLRc144q8Sb2NmPqt2+goYZ80xElFy1Rn8l0h4ysBbn8v5ft2+IJj40Z0guDSUEAXqdh+fdoY
H5O1gFWjDmOunV/GZSzl4Sq0XyIB5Nv3uuSiUFK+uX9/IwSNfNqMM3LrLjRBtONuK7w1xo7omPel
/SM5mLGbiNIuXe+IToLReD1HAjBkQfhOkRaxZEBjtxgRCWqz4mG1i1uhNlryy04nbzhBEMPn8woN
yknuAvt/e4zQ9R5zeALzqRv4YEy+GfdGD9pEa5xspK5jcA1VbL0iLpg6i1kEDIE2GTr37+hCmHAN
BuDhROLePGFP4LglEsqWVIo7Q2NO9rnJMSH0xXOUGJSIPoUhpRCOshlnLaIIgAxoSAbE0uYRAM8L
RYvepccg5cW9DYcryvKJrnVF+ui6uje6KngPJVQWzmuZ47fpDQK+K0Vv4QneIvWU1osVEfEEp+DV
vftZYlIbX33CzhgzQ/jRZKP/UzEGNJcuIfC8WS1XKqnTgg61NAOXMYfxelDSLsyfMC2+vRoUzHKl
rqYz735SC8Mrp9SqHti4Y/I7gleRxooKiCLd5XKgoiMTMDfRTRNiQp5UcXuZ0qOIiFNPuKzUMSv6
psk9l46AMFMWRInJExNEWHjpRL2GVuvDPl4BVy45wMsDmh9r1NOCC57+SbGCcaWvvqMZXk65Q4EC
y+4cxzR1z0YeGosBFi5wAGqVDsGB9zMLHTdWoOcVG4GRpJJJ5iSvA7FCg/aGRLyXklkr3nup66Xd
0S5Ub+enBMr7ubQhivDosRNNOHbd6aP578Bz1EgMb3t9Dlhtg9SgDzZsVGMelAuzoy4/wytQGkjw
FlJSxHWL+O+aLTDcOTbiSRTaO8He7lfVkbBdkZJjnPupKeFz8qI3i049BpkI8NNR7eTXOn3ytpfb
EkStlvGEXnGqBRJafMLN5tgcqytyYKCACVRZVQkIuGrdNQw/Bz7KGOxDWvlaaBboyEGVnz25UuIL
3zUZxiBU1dJFHm4oeBOMlZy0zaeyJ0nHREXhhxbck6Z3pjp6BP/RouU4nYkGh/VazyfR7cumfzY6
kmy0NwJjLa/Pn4QxSO9ZVI9POGmUAjEjOsmffuCLKYPqGK8Xc4P0Dx+nDPnAJABRI4v5IN7cFijs
fNO8wmX5KXToFRzQdEC6E4dCQ9jUczIb/S1PvuzejpsFGL5NXLiCYF7fQslthwD5erA5B9UHTktA
Ro4XOKVpH2XfwzOwofRHyztAbjOyXn6S6JhxhvQgnNhlEe3oFxEPUrlhyJbKy3Nfclk1yi2hY1AA
er5ckOkkQ5dKmJDrbF8u3+sfCNyWtNsbrUtxJoUoplf8Dw+oHPY6toXpAhlT+If1ltpdtlVjqQsL
cqNA8Q6FZwXuU7R0/LcbZ5jMRLrlaJYnS55EQty1gXvXjTpYVFfxMVteGDbZUugwzkCoRcBUTTpy
2sNpwi/j0VEXI5eqv9NI6ZVr1p1I8/8THrJmIkWvyytgSAG4Pki/OrbsnWrN5sKynYng++HWXWpM
vFfD9nY/JCJzyySpRDuN9B5SPoGnn8BRJCkQeK5rI+dZQtuyqq3QW57T0tQxsJQxYZs3aEhe5cis
oNY8agbkHOZdO6RwOlNpcu1prrDqbtJwV/v/vJiZUXISuW0+MR7pkpKOj2gQVe8mkh2IRmxV113G
y9GXNsvMAbsZUv+jrYRbSI6C0rptGwd+e1OvZ0SV2WN19gTpSN5FlwmMHrcAromMPzZz5IRtJ1od
a+1uFeyBjErw+TKlbuvPlAdw1NUAdUBodWi7DWU5kWh+vuaBGipTaFYP4KSpS3XJ1vsEPIvDQvSI
dl6C9lZFpQG45nvy53sh14X80wVBPur70CzdGcSz8YYyIjPDsgCjx68nqpLxwEnU6HNboCaNwz4v
2FNF6oI6o6/F123IUqJxunPZzJjyvn6Sa3M+xP0gdOKVHp4jp20uiVZtDgGjeHPm5gx/XlRTC8Ge
LYCqE0mYHTTG4Z2m6aI7L0fVLHgbUeNKdgxxqRB8Anew63hnsNUC84qcAYgFYl4VZnggt2mooj5m
cEhe+SWcHRrjsrprnWWqtFma45LMfi1JA+tZNPosqf09aZi7p9AK4gnFLXd8VJ18WXetoCMA5MoS
z3DFaBt9aXejuRvJt2oPHaexTk8H047pxykN33D1n1Zqh8GsFJldtnd2cEvaY+OVrLexrFdrM+H0
pBC1Qif+cZ60lxmU/W4W9FFc1rKobpy0XGenl2qDiX29sBI6aGSA6Qnrr0Y8yvoC/2hri2hYfiq/
3B918/Vo65H1JV+wDZmmv8Fbi0kgG39pO1yzYTtCxap3PkZCGwgTaOPstkfbEkGNCDyPbJD3lulA
MF5aHrOSu8ff/urHO6sOU6nyRD22SbtNp0xQqjLN3nhygGAx0pPn9iipmOdVx4isiYjhLi28cUxz
h2Ub4WrmooSVXiN6CdaVUsB7xXSE/AtDTYOVuo0ysPZ5QfjVP6mkPUwmlg3+UzwC8rzXc8WLmjuU
67+vASyl2RRnlX95WkjAfsNOxOyKeGEDa3MgVS+9SZgC77NrcGM5xI/ZqI5uHB4CkVMZdu9VbPDa
+ggBE0F013/EmOWqkL4nY5DaGB/dl9dP+iQIpGLfqpKlnT6qBlY/vdc1eecUq8p2uIzNReLde6cR
MlhY+Dw9z6PSgoQDQhXMaO0A5co0r3ftm5zd2VlP1CPJvB/gRSMm8b6Khc26lUem7lwau8fUJLvo
LkC5qeoqdRjWsx+TULxVdf3x4zZ831gWz/GFg9h3jt/XZRiWmjIucCoac4dwVDA8V6pqNbKBYIgx
83xPmo2+1Ws34J/gqlFZjYkaXaty9x4z3iAAwGfRMlXs2bN3SOJiLQ7/akMyKftLgU7TO9BgoVX7
5E4hEoHsFyQc2gkRQnOHpppvn1ib9RR9Z1YDMalT4PwqcUuFQAaAtpWQkRER0tK99kl5IYiUveOM
Gy+4TX8r4+W4xU8RCiwk8+Pw7YrX2/gO1Q9eutsY7IsSUM8GE9IRv+twf1P2rjPGzRCrOW7mU9Lm
n7yIh3KBp/rxqT3SiZTgJA4rmy7KvDwxnCSXXgrKMbO6N/CK8sZdtavKAgJTiSKPXoyx1gt2I8vp
t60tm/A45BKtfqa2OUqv5O5b0a1DmbuM4+3CpeOyYfwB7zpoFEDxWM91vydQFODanmGZQKw5hvl5
ibGBB21U0y0nkMTajZaLsMUFZYpRyr98rMblVGnHc6ZXwJxc9UK7IS6/Y4RVJXlaqYg6f+kivMDa
OpNjwSZeEqwqplenurbEp2CgMwd9LYtUoG6Ad1frXdNQt/6ydCvD5fz9Bv9b2FD2OeL+caKfoxJg
WCi/QtpW7JtXP0ENFvzrfeqI0xi6lMTodG9dCNMiGYwhrAihaZYtx2KwPz+aRyYHJ9koWNfhmzLG
c7L0+416pTxdea/bKy9XnWhVA40l1YqklpGUfiOZgi9ze6MOawXgnsZ9eJ3vPQqR6fuWFBnixeND
WnkgKMq7/4ErHsd78XNWPQ3l5FdFRtNnLO0dKaNk7BbAvRXutgbPXzp4M2TD4oeFPyAdxRFTL0m8
Dculcyx0hDwpCZgaHYtq4GH++ZOc4jZe34OXOSNKiUCTyS4wJ3TAFZgaVd7H2IG7F5vL5JraQORS
AOj+v5eO/zrepuZ1g+FWjIKDLLcKLUTH7qR4B0zjsx1LH9Gry68XqZSPxQlzBlTC+ZTYl7zjh14g
UApT/i99Gox2zqcr4/2aX4ssk84b9bcZG5hqfXkqOSKQAU7zTURPzmg++DzLwzjWe8lNaOwiv2Ah
ptfL7ICtBSOo40BUULqAg1TvKh2+zp9ImbVGM9ds+XEhSvgJe5NzJMh9PzOKep+UR/FidM4hBSqz
+T6RwO/SvgXVSEZpsSuqQ5IPRia1RHLi5Gqa2ikNlJKgcaek8ZhQg0gNF9Y3dHMiYOjJVOwfmyWJ
s6FrI5e3Prl1m5he7yRH2qGGYLCWfJpF8j+KkvwUNMZZPK88klgJvM++bu373uNn1P73QbTjUbXC
RMeSIUBcsueCPLh7xwYTeWAae1vXJR5gkWhk4hTNyPDySKP15wUEPT8Sc7HAFxAQgtcVtMsjzDmy
mEF7F87a4dA5j1igHPdrmUe1TiJhrb6Cun7UvRT0IGBTqZB31JBep73ICdBKkNRxzeEq33BgP2Pr
M36mZk57y4tIZ2qlYd/DMHWhV7ETC/oHbCh50W9xDEGJPWVkn+UYSWxTu14uhjbvtrktkqKJIS+Y
9YAwmSHayUWKOtcUaWxYPP9zamwLmYqa+TkHoeYJxqpbLUhLuWmDDquYvAHBwnHCbVHHAaUGLu/4
qAsNBjrHZlHVd7fGwKR51udgDMB3JGSupIGWvlvtYqQYiTT8GlB0zWaabAtQ8asnA2SyPUfa0bGi
yUVViVUPZ6sGPwrg3EVHB2HFm+a1nCzMkabaGSjiHwjgmljrevaeI9HAbotyzc06ywg3rb4CiwqK
s7COs5w5tdbFVVVxGr0ghPEoBHXsRNlpVUmC/pwduPE/zQPMx88OkM+QjKJr+z1C94T6tm7KC+je
cT9dPl2COVNaIdW9GJZQqqn29QNCkIU1evB9SQ+0shNoZZIPrre6HCZhyPFVTVpiK3xVVMLHkXN3
i5sYh6cqXLhtisI4qBTPA54KjNAspaPZIs2E/2oN/6Wm2IJR3Lk49hBg7a+AyvRnhmUk35K4Ojf6
TUtXzZmI4I30ihbONRc7h82IWQ1INurM0E2BbCeoFin6EYYcW4VMM1aqo2Q6fEoIT4SIhFX6G+vW
gj0qs5la/Z3QL61XsInWZac6X3YWoNzZR7K0aPpWwgamtRdyUIK3KE7CLmHsknskD4EsgxQOPDgf
BJMhk95M/guB3wdr4JikLltyu8whQsuDYRnlLEA2lPkaMTc7NhzS5dB1S3QqC9MBGr+zdJbYOl7w
klpDw15PX8LlbPMkXoei/gNKttGb+qeTNMVcf0JK3Kxmx4Bh2uaVCwGKZmqOD7rWpzFKFcfPEYpQ
pczpwWBADLJFA03lDFGnn4Q6Q/hXkh0qxcGtfWRxcShByFvnJ4F51KwGe5hE27xNGylRlYPWRpTX
EnV7ABQx1AClwaRsvgI+GmFhV4v08uMf2hQWhOk39ugvL/KU0neaSS5DITHdBtaJku5aOkqr0/xw
vlTnmzq1AQA2gd0QOWKNADCZDxorjHDQ94wNaPlRJhTkgz8oNYtkhWq2vans13TuFJOaeG+UpPdo
7Xc5Y0gT6Hq8skfnLR2yQCY2gB4f62sFRNTQxdGPA/cL+h20nmHmPg6Kl2fRTS9kOWTgwJAZVRJJ
Y5zdx5bWmkJukLAXdg4UrQeaEBe3KE1hrTktsO13Tve6UIlYWS0QYAya7XtUBvMm5nozgx3wmpmO
OSwuiefCd3DXMKtQ1URiuyJfzRRqpRzI6LbjiNco1Ku7rDE5/fdx+4Jm0oj4TPPYz/6NDj5/i4Gr
6fO/Eaxcbq4fr6oBjThNuVYu1+5R+U4xBCxPmy7hNPFgo1KEGejVF0kn4iQnN/2RCyvOyGqgx10m
CR4frqln5Q+bVm+gaEnXaAXS6Id1X58OKiFu6HK8FwXrLShvG2x8tVHn7ui5rsTxyyA+zPkKO42z
RstHCyGW4WzHiFzPCvyBafZPhE5XJKVyNtSS1E7jsIptHL9S9UO4He9Qi0iqRUbP+PgePJQKVZSZ
x0Afctu+h2TB/OzUAoeFSWVVZeIrUyfjUGo+ukJYg56Zd7/BYznkexbR9uz22qvIOQ8WeagsBVme
XMn7wNumVaoA91x6ViGqVqdrdvrzpKCh/191WBuEt/tpYhR9a2NW6L0Nzf/l6xR01rEhf1z1OhpK
FVXr3GoC1cBo+0xbSXaLHE4F3J/94y0W+A1aJtzc+g0lj6700gJVX9VYsBxU48wm1F+8TR/c64Kx
DjFvBHUFgbDRrDeT7U1idHpwul41plGX3kA4WVJbXziSveMDe/qukhR+AM7fVU44dvVQ7vW/YJgM
nyizPAKgzWmVv2+3qCkXWO4Tgkp4Sij1nEZPgccqGy2ztaM5Ph/9DhfsyYBROvYWflAnL+3A4wM8
8/Ykeb4rpOusy4DY61K3aPpfaFtKx/L9Z/YeH8FgOEafaD7mJzdYiybdpthqPC9bbLzEjGkNyFt/
3/nK2B2Vdot8LXG/FYsXQqTicYeAi1q+VC5WCxQb+1DbwIiEWXsV3V2PAB4ln9B1NNFzHJKGyyS2
by6tPJAOX3Cunx2z17r+r1TPPU3nSFBKHi596Rgx+VJnf3v4S7NDgn+K+IYq2bs5JDMiGAEKPnKG
ajPY//7iyH5u1GhNyF83az9rB1GAe8Cv73J3uNrYgWBsG4GlgXf2E+VIN1/VQQ/xaohhaakr7tgK
hIkJ/X2rI7RXSfGpoHMGcPiGCYqHeE3W37XrO5AWr1FmGsQlqXKYD9O/btIsnouEYL6cys6FaORp
uMUHWZb5R+sB4u852fiPNSt4IbKfDreoILeME/eV7mjf4xDydh01/Cy8svGENCJAt51mUjTOK6Y0
VPRtg2HJWG/SrSR/qHeQkqhz2zWOzKmqoE3hj0DOHNNQQkk/f43vI3/qkGPolmo75fB2Hjdnd015
3EBtLld2WzRfJjS4/cYZ92X2lmasroAMK7tIUQ7AF32GjiPE4HQpWXUlgy56XH0Qh29r3b18+V36
MaRWriZ4ywttlcrpQjUJeQNuy5CBftSWVtDFra8Ds923WJc6C0726yZUnSTcxFXCm7yysat/rpDC
r+O44Oc4UeeoaibLLUYP3vd9xdXcLie0gKrcU8DYRiPml0y6U/wRVLYCjtf3tKh7m28cFmVo2Soi
Ze+WQ1sRZqRwdiXtqmerq2egHrkPWZnZjgGPgTq06mXIkp6xhWtMc6e+QM2jliFiNI+ysKMM2DKj
xwIPl99N05439YoQ3cgdpQo2CS0Fa74PcnPdq8hU0IGtD35EW/GFzLpE3NC0YXIDWWMMH4CwtLCT
1gTrUizmzIkuQtS0ZCoLuNiOrIEjB8yDhpeTae3jHnmyHVgPYxuEaQOvB1puLKubQodJQwHD9p/c
kS58vUep6tGsQCZUX1xQo3pstiNWdAuqt1o4KyeTy27VJysnPtsgZnf0i7UqVUcYXWHcekYluOvJ
yOlhrC3HdyV9ipfd355kcAOrJ+fq3+l7zwLYuBOL8NZ9rs8EwbtQcxBjo4O/rPmMwyP0spPZqeBh
ItOaaKKRxoAEWKkWhIaadoSvgBMappaKEjyTLnoEv2I8c6/2Gl2DxBDmK5pxbbLoP/m7W6DDoYiO
VDTaSHU9SHtytJcE4hj6W5uqJlb1koTBY+L3cMsNNfQW/2IGdNFyX4YX5I8PKaCVS5ZsSCwbudTL
3pPJg6bAUKR05wr7uaQyZjMZieS4j26sI9FtdmTkJUQOnR2KoC4SqAZOgb9I+fK8S+IImtbtpeUl
bwXwxHxlO75ikUnGF/utEYwaFx9UZr8ib8VHBWcdRYQto9+UXUoBllIvUoLYxfoDRZSpWR/KXfqh
+Q3aNeSoEz65vSkNR/b5HeLurVe9QcmrKU7XaIRR4FIsDFhQOoGZmeEBUNbjz6SsA+TZrIOEuV6+
Xb8ADjGomJOGpbaOpt8Q+zfTqicdvNw31edsz1ZiYfxrbnn+4Sv6byV0JSuQ8JeKRSFy10o/DrMx
/231VlWovTLHUTnXsMZoyeZkKr16t2fMQcVXqBsqsFZDkVbe+Veg8Tzw/9iAN/PGZLguE55Y0z0n
iBkWadwKgheqipS4esYG8Dn8aL2jy4WXGQplk7XpNftdQXd9MQmjQ3+dojBMVGsTsL6DyFIhIZdy
ZsH4uqRH5atWmMSSvsNrrhB+4rR7ZAPY03jP/SNTNNqUPF12bby7jOl/KNf0YTe/nVIRY8ZK4zJU
+GDO6JhIRjH09sNdSDYhuhnawZDxwnuO/rifd/YhRl5AWdKNN8lwUmsaExWdwbwRJGvfg+/k8tPh
/wRSTrBGUMcpWL8PLhf5mbaXe1DC1rm2avAR+v3aGrbe9EPzJZwMUGko+E0YL3fxEbpqxiretMFG
qZ3RqnIeWBzUE7bSpQWgHOnN+cUHsqK+IZmemeIHDivJRbi2AChFQcezcRoTGmjtgrubSOLQAqk9
tSmYvb4e3RiBq2SUtT/qwlQYfKM9zO1AmbWrjHAnDtqorFZWv3fUk5LXzLi8X09W6rJRb4T5jp2t
xCEg7yANvdGS/eSsyn9bHM92WkvlwaJO/XI8janimFPn4mDcZHIfIuYuDrlY59Mo7M87SmwVJTMF
u1BoggAXIsRyV2B1a5L/jbbLW60ycmewH7PXjXFGbYFdi4d80cZzVQe/3ZqIrYJ/u4tE3EEeeX6D
9b6z7Rmr/D/wMLUfJZpWaoj3fEPeYzw3AG5kt6IVFKnxxF7LE3MgG1YjYxVAV0lY9DnwfEduti6c
GXedtMbuvcJtgWPJTx8XAXeO5/LogvYIY2e/hXkebM164IKS2NtQebFYUb7htt/L8xsmmt/Z84L/
MI+4ThGzNspjCO9aixKJ6ccYJ7jXyp61o7uk3iRvsQM1AAU/EKxpDSNKks8m5e8bn3xotggyXOdv
rNYa9z6mVeEPOVs5RBVFTxIlqWFe99UuO9VhqSCL8ugJiHsGvN0Zu2E+8rm1AijfED28T3A8F77D
hap9/c2ZZRnakxWknoLv3bdkMK5KyU7aqdM+awgnWxI9e4lC89ldb+J5EnRv8F1AePcqW4mbmy5t
6WZKLZmgR8nscP7a4jsZqxlLKL2FtNSat53sioXzdSMz5jUUkMCB6wauoaLqHh0CDKqSpZcmFNUc
hVW5oO7BxyQO7P6Oc3vA+tezeG83DtmetXKgLpSoLc61waLyCwqcNtlVln3P7lnD/05DC0p33Eip
GLJxUZ7LVC20Id18KnVrxZb+dDjbBzdm4aia+uCIVhg/DuRhXENqZlg5I/CQeDwinXQd7EWN6Kcg
65r/D5in6bVb1lxmoC97PjGhUkGpeNtgvfaZH/bO9zKcF8joUeg9F8dPgY4guVfOHNrbn8kP7ghS
GU6LA3oGoaQTEfGbjhFYfmkRCV5MXXvrJnoG3oIU5fxLWqcQJS1iuMqf7wzrnVcwWSH4WHvc9aak
zAXGWHjsYRSX3voKUMJgdYXVLipT/EkoMQtqc7PBBbJIzzmki6qYQKJ9wUs6MeKrnAg1ZMXlX+sM
rvehOQOT7CVar629PHc5NmS7bjrB2N0/GHk1DmeqxzOZDWb2dFgPmplTW7P8/DwSY5eg7F7A2x5L
9PtUtwT/eCZg0da6+0bSSuxro8BxqSYTRgOfCyQ1+NnBjaaddFAIaUeBB6g5wTVpva8WY0Yuw+ee
8B2Jb35405zoNF60qfl3HPwDbNDP43RjvE18/PHImyRnTSSx7crm9D8oHNW4fJ0bMTMzx6ShqyKI
/I4xKkdBgpgIX4DVS7ykGNX9pzxc/xPsNT0iCzE68bkpToUQFPvY1B94LDl9xqnKrXHfFqBFCXY9
yJYJqhfaKL1rr0gc+2agi8nFMjfbwYw/HkB8/EjIba5azsRWwjTb2AMlDoDzpFxG9MzCKqtIneWS
0Qtm48wMqaL31gkEkZCmO/Wo1rHAA/6Q5IhbIC8I23itZj07ArON4cifDzWbWe2mhxPWhLP26aIW
gIK3L53nfGKiDUKvp6lzwEwfPPBhu3Zk2EC0bG7z4pZxVe+KkvofksbBoRECPnXuYsRMxafcRuKh
D4BYylw2gINV/62vOUxjyciGy88Y/TbJBemPVPE3KvKODfZGFrmM/ujMYxPduMN2oFOAEJhvfmdQ
cm1ARC1P3oBZyMnKBUd7rZNitHan0fwMqpmPQA0adH6idzSsf8a+9iv1ObrInRo2fUxxe6G/si1z
Pz/F/tK1DkfIsg8tx+tWuliN0qPx8T749hV1/OkjwqNA/iz/voap22JeeQoYws1ygC9OEVKzepma
8NbkI/Yo2Uc1J+FxsEznrhbqG+OZlcRprIjH6DpC3HpWNVE4sP/eKwMgodU+XJThRzX2RcmlRtWY
WSA9UHoQ1x3n+5r1bPA0fnUpU5HUXI0jlzOAOFn3eTqSfXz/KDUP8te4xjK0ZuRGFxMlcOM1u7cR
IEAgMJuZia4K7mzdWugP5gQfNf1FTiu9e54+SNaVdnOb04AFV5j3TfLlk9TLnq4DeOQSm5fSt8D1
w+K0FoPbe3pNAn/i/ufFiKWHcvIIQDTuP9QkKJtR/p9L0x38nrzU/wlN14snh+1OhBfSbDUWy9ha
aslf8osOs2whAct2qhadu9pMXg5/wrEB8RYtjKKdGK2xLKHm5GtfPTHNAC81041nPmVYb61Qo6Rb
Ae9U/qwrk1tsrYElxRuS3SBxkG85VHKCojG23Txd5pLL00LrQ8tMcWX3Ehd7MOPXQemQf4jtfNiS
8LdGk0vbReU7dPg+XyAoDddwbJtwaz7T8eI96JNfnaQA/QiHKppAxRu5XEAl81TTsGLihcqajggo
NdLdziASp26Isv++PkZD9TkWxC30I37SM+578soSAT50wwkBAv9ps91XJTnGeY1wdHKzB3hax4Cw
u21scguPAG0xexujnoRgJozAVuJJ2TBRq8mepPgecC+vbQRWZ03Ien6915iVY/b6hwWTgvmsffP2
ye2ym8eEQrBov+8LzpImwZA3vpIXIhimor0+RyEmGod6wswhSr++poKyepax+eWQTIlJT5jrKuYD
KnjCjYi30bFRi4bhAYX9L/VW6MMrTWnRU/xZXfVNldhPCECDKF384rXqflWzHqVaiNVq26FzPm44
PwtafZ1EQPT+n0iACx3Heqi1oUNEeoZ3tlXC7NDYuYkDBilOIauOoF8v+okxoHl8rpDpgiajH2nW
k2HSOQ7d9s0Q6G9mTgKmSTRDRxV9dz/dhJQ4clpAJYZpqlDE6u6EsuHqtLriG9gPMxlWPIoGAFZO
jr6apanOmkaMh3jTbvbSbWTe2KvMv05BxnynI0T5VRga9OXCL0XsRUvEBJK+WoC1T8gyrIrZEX5L
miR+ImesBZAaoTlwIG/z8/ai3VbSwBlBAOLgj3x2B83jDdOxE/vy23k4BHcMy+nUJilAy+xniDoI
7NNoL5tW5NK2MWp39SAyHO9ImD25IIUpcF+f2xwya7GcuiAYjrIzu2uLebsueH3WzQb930syjG8M
+Zo7XZh4X1KfC2gjTGtM1d6Y67vkiO2H82YNF8nS4uyUGSSF+vE+N3jSp+wSu3ZIYYFsanjnEQZO
0z1+tiKf23yKX/R7qqsI0bHT1CUiWTHCwvKasOXhBMrlmGBit6cABKXfQ2OagCp9B1QCWKCMy5eC
sMM/dWKR+YZ2gVhbKTud+uXeC6bq92lH/vxZYqAG5iwLvED7P98Ywaabx9KWC4Q8ex22pgD/seCR
D0HB+QJmaZoTu1gQ7LBXFCQvBpFQNJXg1H0raTl9p5CpbRf5YxwY0ZLKdgIEQqzhuRCPj5RvhlNp
3R1QqKOh5hK9OqRMmsk7vXPjijsJbtmnVZ9tQ81Wb7wgPuy8+ChzlS4OlKEQLk98PpHFR02JmDby
AyiDQY1MNUw+jBgKhLnBRVr/VNBRmiF+75fe8tcB1MrXTHhKxGEdDLbb/se1DtwvSZu7zrLpIgHK
O3nSur6w3XcNTxQDkdufPfHRys1ehvXuqEUUk777wb3xmFFyXNGBXCPzAB4uGjs+eH9Y550yEDTd
E0d+K6HiSxFPt14WskyNaAzs6mF6SObi4okyRu21Fcl67wpyHGv2cFDZrxe2s2w2UH9aPW5ZwVTm
EVAwGT/xkkLx5tBbt3q22hHp5F4a2kXaCU6x6/PW6mPX5Nh/0j0XVGbHzj03yS29vs828JEwh4FS
mK+yXOs03mVJWNfdAbJcjCxHp0rlFhRKhPmvQngVPacFWEj7y/z3xK3bo4aw+urowRPRlcyEChs6
8ssXZ0OyqmvdvOxCqe4pCDabeRaGwNmv/40MiSBhzRLHlqFiAi2sSZdnz0ImRBvici3DaI4CIjGQ
L7Van1D6hX6dhB9unFJvlzP9TblKh71DccFhbGDTlO5noVLjXZrDSLabQqT/oMDTyV2uYGTbyvgR
WQR2gtx5FB2JgRJYPUkse/0V+Qs35EgohDmPdhBcoHyhymujYK373DT9kmLBxOWHjYt28kXgfm1A
Rp+5e3v8AMbUbYGZnnsU6j17R72cI0k/WYYxpIA5kyLmgfccyud/DITMrAAzXgFaP3uv+I5nmWjY
08Plr8VCGv3TQ4o0gEV65JDovw9jLMoYPGZWiNuvmIxlkiq1hE26t9YGCf3fxRZUMU6dvRqOsMQo
dHDcsY/K7CLBu74HT3FVny0yNPiV4H4C9BT5BsGnC060I0YscINJiPrxfpojwSy2/6FhxqE4x8Ix
wV9J0A7xOfrWbbRhGv0YpvEbEe0b5GDBDKbGro9mmu34jdL7TAfTxBKWa306N4UwJ8I67UntYoVp
6tChGOtMnhUb97MEVLwfAVtyoV88ZHS6Axev9NGzrc+PLF2Qr+i6IfzdbxuXrUnYJP4quX71Hs4l
E/4R26dZ5C6UUiARDcjnp4ruqO+auWOJls62LVSS2FkR1SBGxCq0XDEhx+5HE7IvOwWXJ2KA5ur0
5uReYEYgDSPivhcNohY/ZP30v6CUHC9Vu6sX1raDB25rxud7eEPzMO/7rJTwDb8yIlyFWCQvcm1z
yblhCjh5KaWGOiEhEyeqjTdEPQKUEszRrCqvrvgq0QaHNj0dDgRjMc61/l6hFb0N9zEf6dn5iK0I
bUaEC/H3HpyG2Yam16+QzeXfh2HAtj56VGRrn8qxCverLfqCHRcl8pl+23QEjBNYYW63wH7rTPlD
cE7rpbD+5o6MHJCoEGuzh8DwMqbaucYHXyAExsRXTfVb4WfRwcstXivU6Eh8PukTJspSqAqPTPeN
HO02yCaco6T8PGRP7qyGlIFxvK+AlvUpG19yarfbQgY2+tViYovM0spWMsNPtt/SFEcA/sHEJhx2
/Tds0XT+vQWRKfLq4TJLs4GOGEIACuKsgzU0vDViW928Oyb000ug1QQlndUjg0L0Ln81gpXl7UZW
9xwQ9bL3s8Bp0UbYuBOjGwlTEOcqdYsYYmCjbAnWs2DrN+sJTaxVRmmHbhHW5atSQIaYLD/G2FOG
dcqNEbY3dlcVWiUF57IdFwV5HUlIUZhmPB/yf6P481v+TUZOmmQKUorTVFREyDz4f2t4TbRMOvbg
eKjg35MkDMabrVnJA/CUZvsUIVmq1CnRUpN+479yX2yyxtitM/Qa/aHx5Nf/3iT2aiUppxPmVJDu
Lz8kSErY5G+C8PlpSaU6WESmXMzdBdcv6jcMn2o50yEPeoonGNlS3MML+9LtqZwghhTDZuMUL8Pt
Z1Iml0QbiV2q3CVECbKqCRCNSN80vQgCDUVQNx69rVbU5E5W0Ai1v30YBPsQnJFxb548Tdh9Mo8g
nZsduMUZitPcCTSNEHOmmsHgJBSRFBdjl21K7RNr3Sb34QgE6hh+pPuJkhxKBwPIjXseVDmv08qu
OzsLwSJ1yElgXE8YjV4UY8zuB2V1Gk+X+s5Ioowc2saHxiJzWWYTZ587Bw8ai7N5FRp/HG2FKU0K
l54QyR3cmR52+JorG7r2cBUmYeinrcY+t6jDtPGqvi8dlvRiTFf6f4R69BXzix7xgb+uvqytmQo0
nj/RzaJOjNPVs35R9/mrXvHPhKh8gZrDnR+OMtflUNQLnGDKNtPfVrZt1gNDCI6qRUTg1Y869INS
Rn3KfI30zUbPhHY+7/i9wO+VTEM5VYi7iLzbaJrbmEu9V8LR7QuZE+Q5COdtjwmOaA5pxUNR+bPC
VGZvgRDMS6Keh1FJIn/4y6gxAClKj22Ni7/IbioD96d/xuLLE0bhGs9GAo5LX3j+i/1e9RxJHxIg
sXq9GcJfd9Njuu+fNNvUnyDZvXHyEnBfFj7Krh2IQKnGlaQr13QTM5EiZcthHZ+6SksqmBGaWOrV
kh1MWfzRSrwqTHiwSX19O8CKdw6+uLMO4klDwSoRd8T/dT81kiO1F38RcJl2Sqe+GxbcjlUKtak0
msc0azUKuuhGcGRm0ipzgHDNT8XUZ/jWEWCQUS/tTxJkMGd27IUgpZfXN5LzfM87R+ayZ3N/f/5y
m5X/0aDsgz+fm2N02IVFBeA7NNkCr04UWPTDO9iVbxcJXcc7mdLwBnBDQBHV32SVNAUnMSqgi0jG
21d1YblAnGhKEiccS+knOlNVdquZTAASskjPQ/uzHHXu2yOysltby7cfPtLSAve9QWskaqwzY8EZ
KOegif08kbKqJYQ5ntTZFbtZI4bwpc1xUtGv9gfOEVGnZDaAbpAa6+UKRa7YrR4Jd7RLdx5e1nS4
SdFot2RSe9fGodWBIdUSl9jJlCZh9jVS2Eb6QlrqP/g7rOX9FE8tkdlp3+5Ul4eZkCsdIbqEaJqR
R26llhdxA5C8vKQgsWjYM7d3WdbMGw0OfGimgW3nNaVNJ7Bg0bwN43myRXhrYKUoT8bmYJL9Ejbe
4v4qQl4QgxLlCs7wq9zy3H3zYb+OKaHBonLUhAe6+aSs7J2iifEdU0O98o7rBJ+lKIi2d9VlTbGw
iw5iUv/jQY2GM2TIPLY6Ew6veBkLhb8rKzljay34L4+Om+O8nhp5wxXu+ilspXqE708IIVS+Yoj3
SPeI3uslFW9EJj2YixjOw+5rQ/9eUZC1nj5EzKQ+DNhbjbian8HhA59qK8OQyFGZovZyUmicHsPM
nLtUkfqVbNj0va4lIM4t637zjWLGE66Xl4IycmcP0wj6RK7bJ3MvklWqeo4KjIxJS+LE8/1IDHDk
tKMW7Mnyhov3oeR+N+qsz/81U36bqJ3TTg33xhDqZLyOCw13hy6ozu7HZAeDrIHeYVFdnID/mmyp
YhO9y3clGTbVPkowQ+t5SVsVH9okbOkClR8Op9tozCTSbyJXbRQiKbNFIAxdjD7gBjkU5tFQBVmZ
6TCqA5cV+nzR5s7LJmIzQGB93KqlW3lR+Y8nDcOrWsMHC1hyElkOvU+G3Wdx8d6ossE17U2ECszZ
5TY5ZwD+v3Iz3B6qDC/kmSpUYEiEtVx0H2DDlGT2AZH/Y1GpeKvFHNgsO8mLiJSEpbQ6yIO8VMxA
G2BYOx6AT5K75e8fX7oabBJiuDR7TO8kGGn3BtLmVsGiMQsHZNnF+wBqHNVkjvV6onOcArSZCq5x
PhAmYj3SvQRx3BG4Bjmvf7L7U6sc9TOCgyHop5pT/D15iphQzCNq6RPEYMD/ww0qZA9V9Estf8iy
VE3PJZujVPAaASWW+ghhbx89hBOZgTRVAMJxaPDJaGl3hy2fYNDRG4UYnenhaWMBdm7KS+Hfeg7e
Vx02lS5Ymk6/knDZSdgHrquhzWp288vQfqpZlvyBl8qcjlF/9u10PL9N8TYevBDqWnxuI4KIzQqU
EfFFKGeS83Yo1vMBp4ochmhtdyc/wnq2CV+O7P2Ouw8vyXEGo/h9rHyAhV5fwdKx4pVxx20H6n++
JycbAUx6JGusJUf276MStvebRBVhsPkqy+C7rrDsrAwGQX0+70PEjM+QwZRjSunGYqPxtReseFGT
ekmjLog99LNauvC99PyYsL1Om/6SOF9Bgt/8hU634rBvOhrkswD2jpsWi88nVjQ7Wu2czU2uqZuO
0fTcGZc2dPEwRMrN7Y6LT5GIEXCpkIf8I/bhuOXu0QiOt9/hmYu4Zoy9BJs2TP1Rng31xdYwLd2O
ck9O6xCiWlEjO8S3hsGwxpa/OKROHCxFjf09r7BwzM1u5+K3jC8gBNHNs+/BRYSX8n3Ic7FfspJT
DSz1zRo9XcBGeyIsM1GhTXBFEN9N0QSKAiQoUoQiDVL5+3k68QJhytJ6c/wXuOrdVuoc3yO89eef
6Ym11+1OW/43tRGUoOuY2Jbgy8RyyaX+/AjkhMee4O52pwfScn5tL2s+vCgiZNdD/xfUBpmu8QOT
3gw1lUEGTQWeNIo86VN98lreYtT35ImHxQUwK4D8pEkb/Nx5QXAfQ7Wa/SAovtqGubayyLZWxjv+
iQi/K5oRDsCMsXG5gpuQkpbu4CvKgoVMXuHfGKBVEZ70NaVh8Rm5DGhZYSTQp3mXPfPgLL0nigmp
ocqO6ElLXAGekQX5RH75Sn+aJ9ikr87gW+xWzwLa/iNlSRsLZrJUYBgkIdmJfv0DBxZ00bcO8mds
AhNefoch2X9RzQJ0yevIMZw+3r2ssIqe+YUo3WRsWDzbZu1i+upEn/y2/j9nNwsWzXSekzrt5ACO
oVZ5h9gzlo4CQzpIPpVR60X9tBeRmi32+/Z1CepVz1H7+z80upHDmXILFmt3JTgtafGAiRQZZQA3
esa5wsA5Ca20sMxxdRiLK/7x0Xh8geZXmLgH2NAfcL4BcWbPuvmMlCZPLu5iedn9oLtGCN5QJ9lk
cBPDiY6yJDJp2cRyY+jtgT0tSVAk5iI1g9cWhdYbwkfW8iZuyEGUpRfC410rw0fo3IX1VF5+k0e3
4bjD7FUkI1TWUE9lTBkNd2xNRPxLxSx6Q0aR5VBVXrikktodWIQ/gTRt9F7/j+okLRPtZjRResCm
ZR7LrfejXXv8o/h0cVfKJjxiMcELvXMb/6kqaaDRZOO62rN8DgWSpufwNAS+RWBz0LDkE0LkVtHv
UFjgZIMng9wW0nX9/YBUlvA/yy0AwDFYRF2YzyI39GYoWRaN+kC2ovCjMMZcLI2YXa4Pz1z8HQdc
kjYPZ6JFTeg7WQOYRUcKC35wDaWV+FeQ/JyJkyUbfUabrFKzcZUAEc5aMDGkOXf3cc6wu/QeWBY9
NTjWS638Es2qaM/pdUaSeALK9A2VmryZLRtRHVj0xLPyW6DZCgc4TY83lbT6V9LYUFMoHnheWbiF
uOymuQoOqMHxNAWY4rEMF47Ab62sV1nljP00o9ygXhlMRiP8fnOKgtYbFqkI8LWZz+7+HA3vKVgP
QSpzhWDnN09pZ7UUOZNqveVRfG5KLZs2e7fBb+s6eWo1vW/nCB1N/Wlgdjd6qkgBIcgWERO4ah8T
gDJgyQEaIF4DSWYAqMiD5ddiI742t8gNEu3WG/mLU3s958e8+BlIBF6mY/pVTDODgQ9+JhShvfwd
6l8VLzmD3JPCUz3Qm/U+ldTR7HQaAVFgDhhNBF+ZrUs6Agdwz0vISoBQt6+vGlTKJb/IyNTn3hoh
qRFAIPE/o2eRFeROh3xJY3NZoqkjPPNvBPTqQbh6W1mIId+l3X0Ly2lYmlcldSekdjlq+A4D2+IB
xv707NRqJL2cPj8U4iAox/cEke5rOgmEbeXMdcez2QFVsfsFGqvHIJf8DJRsqBXKlojegRy4R7Dc
h1pM7CPidEnB/+swYNE26ooOA6OaCvXjdtawTRQgcqxpCvdC2Aik9PBrEHtYu4TwE+h8d4atLDun
jApSHEfOK6L4Bxg+WO400MRBM8lRCEByOsRczBI/FciEvjqe5ekTBvAhxU1nuNu2fpj3/U4Q1xaR
YiK18dsQaPVtT2sgkG5Wxb3pqPFEaN5iy89TjW1BZup00oTLV7gqdDm5C3XMJ75+zmJzbr6jJIqB
Z5tEA7Rcjbs6Wtb46nHdUH/98LcvboIdS3VDMl1v6MB+sFtGxCCX7EfMD8jo7KmMdx7GRZK2CREX
ehKXFcU+X9i0U360VOW9jbSMMOIjHgA6cCtu5rgB6AcbkLZt758ROVYlMAhFdWJe6WstCzyfGCJN
mVlpaK+sCWTW09YA17vhloXd9IewWVsNvKdFCuETNzqDrmW6yAM0GsJev5yawSk/7gMr1shcF/JM
SWJzUIXgLRBPLRIcBzPycq2oiotkYcfXQqtblQmkiJCHQDoKYwaUcA6ZM7yADgMr8n7RUDEI6Uzk
YMRnJdN5IIn4jOonL3veWL5F7HRPOA51lSwe0mhkxrsl8i95AbqlRqpbJH1FOaVSjY5DyBEYzql7
5wHY3eXQrhJ6SGmh5wgkd/sCyClnjtpkCt1X8xrg9bIWIllP1eEPqm5Kky2hN68FSg5/gLYxBYss
sUHYhDSSujAmzkqJwJHAuTELB4Rsm33ftV3CU1xLq8ZidykuoKtJybYeD9o7iVX2I4tgpRjSbpwc
Oaj3vt+Vz0rfARdLICNbFmA55Jj/HPxW04AvqTOPFi5/8sh1b+sFP2qNM9MrxXj9wqnAeeWeIIwX
Ckmb9+1OUioq/DhyPXaK7UBvbN7j9ZZbyub7WX/rDZsX5KSRKfK9U2g8VAKF+B8F9DhjfnspUPKt
n1blJERvH7dxeNhFSTybFA7ZGGQ0DkC5a4+86G3ArtrYMuqH3gYRnFT7iEFtfv9zq+r92q/x0njW
TMymS2/Apy5NZtB1o8g2oQDKSxPKk19N9jMfEtnga8wwxTbBr/NCrQ+pGv+jAN40KlQp88HJ3k59
U5lLl5VAqL2Q1moQ6a02toRyqiEh1bukFW+Hv2o7+PfVXTqUABFBCM04jTbbRcUtXmW0TYJYzYc9
gGwwwafjrJkYQeu+iteSO+Np5Wf2va3hgOI6PufOa9Ne7oZrnctmzOrMcikbdfQvzo6IPa0oNmJP
F24GqXr/ON1UxYstduQFuwmrdwx2doQ2o7bmQRfYJknJ19aCDEPqLGRGj4cASGbLNHfFOij/KTwS
4ojM5qdSFa7GB3C3dUNyfn0k30w3KBJ+b/FidrAKawLv+QbaCizDTcIoRLa1PFh9x0dHvOEuhQVe
FsugViZkiMoL7dElEJDBlRVOauGdzIiZESDuM5vzbpJxcI6Sxh7fICF5VsQKbDrgYX9QQz5bMh2W
xIl9QgE9jRlS19+BtS7dFVuDU5NUGyFsYnfo8/8GMNRjovQodoSe+TFLmdowuWG58k0dMXidk49F
wr4I53vndMpA09J40mDToMojXBDjDJXv25Un6YRbNeljHcZaNT6BeDeNmAfn3iqsDWrekkb3bHFf
zFKSxWw42zfxC3Fy4XYhBpQaNs5DDbKKGlK9UhMV9IO7SPHaJdY/LlXre6wYX1xK3ihHCJh9reax
L7N8iOPX/vPWHFCBZhun8c+X997Qi82WgA1HNYL/RkqsuTwj9O1jvWdgfqzL252QAMPzCwjTroR/
UCF7rXSeENB7m4xNVRa7l4DR1efDoEyGDyqbLW2F0tj1qsDFNd465wumxeQyoTjS/N2XWZP4d3Sh
CfJ8vLDP9iKr8aSa6BM7AM9w2vsYb7xT2UkwuqdwhoehY98XSvEhDJ2nD6QONoed0PoM4mIqrdpZ
+FI0iN0FPamx7ATJRs0aVSxGA/3KfnrlMQdlDFI3lo1RaRpYvRcxhfk8sDEgJFLrFAVlETf9NnYb
EFUq1j8o2sD7lBGtJX8SwsFGLaEtZQggql4hqGe9zESXmMZqzMeqlXcBXV8QiGL8p6HoJCKMcQkq
ESkRGMpwZ8aZKNj5TtGveq0VV72SVK15AGfJOKMsBtKG8nD5quIXcBvP9WQS0gRHMir2jw27Ca/D
HzPMdU1cpUHai6URSC5F/Yy9M1kl3DTl0PZP8E+nFp7bFWdhxFGXR1DcCaes8xpxbA/u1TgQIc7W
RiQ+cI6WkHxxudNDwVYDs2kOeyN6pIVF8KkH6Gs4tiB8d0Ot+T1KHQHsKCDQ0E0gHhTZDMuziy/g
9A3liqAaZ9TCyQ79fWiEJjCr5WcoozijaSNnqDjPnYmvzf0bwbUX9cXQr0lYWNgo1WmipHZdrcW5
5yWSAG4hkGG/xrowljIjT/l7d7fr5/6ZzAk1zjlpTYpiGfyyGTl2Afdt4U5PNncpvI2OEQI5b/zd
6wLS/lfKB1Wi27qqCeDyofYSgvCgoHI1517OI7bu15dFoO9sJizvMuCOSeJrgwxPaG4tt1g3SPAo
MDLDX3EbHfJJT782IZ3G9QGvcPWBxd/Gd2PRaa9hogqg1S26Vq+SWlrpgLU7zBRw8oP8CHd/bcL5
XMFFmJfkpHHf+PJrxChCfa0qAcorBod5L7TIo+t/Vm9w0grC81/nuhO5qEHbO9ssufTxljhPd1nI
aRdwhQKlpxZBZEXVxhwSaUnG+w0MCDiCTaWvtSA3KgxCxXJIcJL1M5ExLJ8cfIdK5benC+OY2Ljh
PP9F5PaulTzyKD1ekaArFLXMSrvhptadZYMuYetKVsUM4yfcZOhwB5dCEvyIv7uFuQm4TVr071LW
Mu7ZxS4ktMssPT9RcyDoSEfN6EFsoxEga914XVk5dDvCZve2sP1F4RHvW20A9I2OPm6T9CvQNIEa
3oqYni8bpRiIyKe+GyFZUFTFdWZStJLyPsvAS2ILte1LBNKE3iiRZLBFFoumKopDTf6fGP8S4EJH
/fWzaH3L0TM6dpU36y0KOoQ1AHLSJHUV9bZCLDOnvD4XnPyaUraogq6C7cgikpIr6Mzie/q6x0Gx
PsPfgoK5tdRfmCTQTKbSW0eImKtgNN7bDX1XIrJLC0A3nFY0art9L7pqRBWuE74F8e7AOWTNh2U6
3S4lUPNVlEBa+4kDtm7Fa//poS6Te4s/VGvgoSmUwwQzIIycZR1efZaQ9ryP3Hhr9UEMKwqqpxB3
oXqZdyLdhlDfVkI9mrIHxSgWIQ5flTUDw63iOiExICHzQDxpLc0s3tqkJViVYMY5DZc931MuNsGE
Alif2vTi9mbHfdWsxC1O4Q0r4yhIroTtW5yUkmyNSRRMZI1BVUT33oHYiosTORckzpdWs/tg8+te
8UmDapfUU/eGylrDBPToPCeXNBorbwzVC+8zdgZyxuBZp/nyH2P64FsDv3w1NncJNhLjsWD+OVIv
nrI+aBjvCnv9okqUKKCdpoupifPXXMqFWR6BOVj4V5yTuESibEG0+SWRlmMcKnGVECItkEORNw5B
Ryf0kM2PBAFLOE12a1pMeiHZit3wyl4J9zR9xrp8/TjJLcY6vlZ6Vxw7yY8H8zdg49sMca27Xhss
12AtHOiJ6YqyPh9Yvp36TU3szW87vtJLBQB7oyh1qBAiz6WpJDRz6JKxbqP6MAgk1F7aBo/BKe9z
w8c3l/oEgyNPKcE8fPA2W3H6A6npFaKc1PQNlHIqhE9jkYijNEM8e8RkCVqSEQsqlnWbR7M/HqCT
8b4mQ/9Y6BL4SBZGlmcWQyKwsRGe4ZDTBjlZvCLdNEkQMQKxTzv8VYd04TkLLvUsJ7ab24gBAj4n
3M+0k45PwSqPmnzdJ0T1pwXHsOnE47oErTJwZ1iPHLtdE8DsAvUGT8U5aYZXitwNd4YkwIskX7SV
H0dqpwkBT5/IKBR1Abl9Cv0LYYaTHZ2I1/4E78mgfe2u7zzLXE/Hisc+RWlT0PV0jvdf7XYMV19o
nFLCTO8Ij/QA6Gf6w46axCNBlE9nqsa6ZqzkCMGVs4W7WJgmXZI1iWpeQ78JEjChKW+N/yTb8jAx
yD6gs4nUlfzv89ulLOaz2cFttvQMbeCp9Chk2x95bnY380E6WI8OydRkimt8mhyPVc+8C169e9wC
NBIQ1Gk1AVedhSFuDCoeQ+2hhLZc42rpG2T1hgZ9F+M4mwjGntssfCK3H0wcVD+chuVW3WCTfSdI
FXtxgBlSct39R5+7YU9OHwM9QpJw9yEablNcF247qZ9zc0huBw8s5MaPqYYo6aLYEYylda0BUn+e
V/rnKez9R2XYxozH+uRE1O7BomasnM3cneHOuMn4Zpnk/hsqIMGH90nFwW0NgT2vkDinGjBfT2Uu
CNAAGybf5lUEE57rpdpJa/etha2f0w/FQRrt9tDwJAsmdo9CoIKTBDJXQ624HOWk8S1BVKgrhfaR
rpGkXCmgAIVDhUScSPvmxNjFwvlQ0sgsBeCVGoDpKgCubsM+3czWG5oJ64lnOKy79AW8lwVuAtUQ
iPE26+MLzJmGEASliAc/raSK8Ho/fEMCMofEhlHrkbtqfvRhQipAR77r8IVndg3V5fqDWDZ4O+QP
dmq8LNMwECa8UpG2ZQ4sKGTNfpP61PfY7ObiZ9Vq52Hqi5pNa47DONY5RTipO5oOkAU4dNlpNpHv
I2jEtJAuLKH1al7ckHy2T/4QBxkH1tKaN8UFRH0HxIpSRV3F8rBcZArtiFuwCzji8Vq9aAuMF3kW
9dJi/AuxFNP/P5CeqD757I2dcmekdkWAQCTCUvddtg3JsJhvgqa22lhMSWACib5bgZ5skBFEFk/n
JOIglRFQeNlOLoa13HV+3RPPZb0M1NZewWmeW2Ub+3LTdydCF8FfoGFKI7tpS6ATez/aaP9P1SJ/
rbSxCF9UeHvgM16qboFSWSD2aTE8Zn6lT1hKYAZ3RnKUY3GHAJWwnP3cbyTN/tKQ7hIZyN7Z2Vgd
WxQlX2pYp33XpRpMKOv4EBG1tB5lgadB99XKdypSgilEFmrY+7Wqyhoxc9qQYR53MDs5YiydRKIt
8PgyDCTs5GKosTWu8wpUbsizqw9LrUSNrxEfXlivBCyIV7JjrwV+icYZnm8mTjNBtTSSKSopT7fC
v+Tye2k0tP1O39cpirMiL/+AyPaRgGawAfuGwIWfkmAgI3ZPLrfcodTtB45CIZwsTvw+G74dtuCF
D0kazHM+q0EI4NCS8Gd4fS9WNYKNfLJavRY78H8tF/2OOg05wZiFN9L2ecEChHaG9mSn7EDsuFt/
MEZFqTj99DRnxLDD0kDHq62pprkB+cHglJcaeK/PKeyWS5EY0mcuw8fPpETCvk5cEd8cY8vnRxQX
9yt+2NSqWiB0HM5Ep0pkb4chwAlcyXu2auZsOdr0O+gIM120EScoMHPoJfoU7tpkOa1+ZbYM7wbz
5Ev3V+NUAXtYCAaReMSchmoYazxF13nDCl4G0nztmoRCTSXKCgPg8UH8kU6QBmMTqkLxJVrYD4FZ
w1NoDlzh4hWtRH/S2k6QuF1bSmuOdiL9zQ5XqjxzB05wb5k95VmihlNK7G88J/+qwsdjT/ge+yaY
J9fpf74Y7UnAv99iKDa7QG8MaW/q4lBPf4ficRTuTRf+piPPj+R1xKeeZcjLEpzvDgwlWHtxtXN/
SJdWO90ju8Zu9BFpJ4ri81AzCkZvTaLBDbszyP89g9PB9e/XK13qfrwosSHnc8zBBZaahesfuRp/
2lsawM46gyYLi9Ur2mOnw0MxKOPlgc1rmzy9dTYo9/z6PAvFTyW1ArZ7hgPP6uHaafkvGBFtjx4u
OQIO1sbKH7TmL2QFmWsTl2D0eEUT0c4F4I5uy7d2PTa+ikbl0gMcPJ/F9iehHI2sJdE3eTWXC8tt
SrZCUdufnNN14QGZDZK9UtGLgxIpVz4vCqclX5tjSP6RHcUSc7Wsx2DrXaeDCKJfeXBc7WFLaD6k
h7Ork11UsTtJSXElKB3FFmYzpJ6Y+D+OAbl0asj1eXwinD+7NdU2BIxKUEGQOGoqrpzzQU0thGqF
84nZbmzPy1l7X/ffTXppPiAYotkgIEcb5m3+DNBecx3vw7x23pAPvL2t85N/fj+REOGS6HtulVB+
qIPjJAQcohumx+YodX4vyjBD6vl7A+U5C3ysxfi9CZ2yBc8xHNIUvtUXHDnPkL4G44wXaLr2SiRd
3v4omauoEndjUueSslhNcF+VBJfKa6OpYH3sUGtcglwPZvsJt2RtBRQuNrLzpALIHdzJjinPxq+D
e3hZ9tG59aoreI948ApOuGaW+QhIDLrzSEmmrtJ7hT2mB2Sv/H0avmXQLiKBIf1vpWQp/Nujh8mS
4/hhbCgEhLPku86sJb8qH9gmYFmMLqFcp9TBuB+5/oYuNdWOoKSbEbkkwmH5yedwKZ0ttYcc5eZr
BnmotTenx7hCI55LSB0yLSOn9N7CAGi7gSOizSRd1LCpjIroRyGtbIKpQrAsEDGoKQCvstXrfGbq
IsX0w6ilyH3LSHX/avrhCTktvcBItYvyUaa3zw4XLxQSLYG10Ztt8wh0RK6khDxhiVtQTlLSPesG
abpd+W+SK7/VaSReB7CyxX6aBu2YVb6QmbfITOlL2dCDIi9QxOc0gW8ExQ0Ao5SheD2ZCnI5KLx1
bplY41UZ+vwd6SEqsaDpMkYjczHMeeHXiVhor3Wfp2/Zo3FUDUHO0mc0uzoyvWAbhDZm0kHu1zs1
5lHdQGvMmEUGb3cf0CCaSfUc6LFIjH9qpC5vIWbLTKvSqs5gzmgF2ulU9HbrKN9QN4ISxy4fVgwl
v0IE6lagrXLERJBEOhFUWAB4Tg1nnSCsBE/aoOVE7iVwO3dfQqmaLxIZeRNMt1eatiXU/mbVysGH
R/gxw01V8WuHqNGNfo+H3MM8mfXJe/+Ke5TemWBlOmYKjrITfJfcawv5VbKvuvlvPjclotDvBO0f
yJT+mQjU4phbdV8ddnfjqu8gTGjSaaZDVxhEBsnbWCVWUK/vladX8YdCcAKkyAC+YqhhOUx3Oues
pnz3yC56rYe4D79NNh08/pkS2hXgYU9thSDSkzpeqP5KB4Si3U3UjHhqtI3Xz66ureW94XhoFW3h
p0mHaKSUIO3gtM8czmhSL70Mb6FR2SYPXwY0tNp4ErfyXkZjd1HROfNG/8xnNzhVKXC6e/pLJvDY
qL26UmobxejMIw8F0XVx/v+jrl1Bc8SegSrQXQr+RzfpUMtTpQPDB1Hm2tC57UqJFTF61OxNRn1H
o48SRIQyWTWBb3vV4h1So5aPv/2Euxm7mHTIsoQRx+zT8fienG/WeTIm05NoeT8SZ2YLNmc8D77q
cGiTUfN2hYZfxDUW++niilLU9AoIdoTJwbzVCnYkrFR1qyCPspTVvmxAwrnjclOfdpeb32EX4hii
6lscWs8x6BV5g4CIGNDQCd2yDSdE9s3ArQuFWrKwVddTB80X/2go+uNWESBZoe4qWhZSJm81NtOX
ZKcEq2GJ9e2xBqfcr+SvG9crg0jNAvPPlxFeZ3w3ugpI9SHnIiKaUhKqADPKb8vZ1U4V4f6vzCUm
8aV9Cbx0sN4D+FRxk5qzwuaUvd+kUEPeLy1Qo5EpldXibTBCaEZV6g0B1QMVDhwOrQTYOy9el2YQ
Ju7V9ySHOzxSE6Aa1WJf4kAg9nChuEK0PB6tGzQUc05y+qT82RrvP8/eECd3EWJGe/B4Fb4pywrg
moEQ3iMNvcmXbXs6qrHqhGk4nDHzw2NaJJM6Dz5/uhQqQo4petfx3rGqyt3bEIijdl6qh7ssraTb
+BWu2fvwPuO/5/JL9WwodAmnOxTPA93IFSAM3SHWcFAzB0yO3UdqRYHOp0qPLgZOqdOgvx133580
mC66g2HdPDZG8/w+PHQe4LVH5ZdDkG1X0xuvaxuwDtc3ZK1I7BmVyUvzsjwFY6IVmg1Q63Ki8rnj
TPSS4lZ8v9XFF8JX80zBPYMmpekjzVLhs88idd1/PPysNDLkRz4C9cIn5yNyO+jSsp0gTtl51Cr/
Je0AC4eYZXRTs+DJp/7pggv4Ca+LCBBero09la2Fe3gFBWGZfvwYu6J1dlxD5UAYXJQX7V/zKKPw
guJzNaf52KitNXGUFaMR4y6wL1Vyl/1xdp1nteUJP/PCm3xJ3OOYQK3sUPdttehR6zb3Ly7aFqpc
n/zFHnYDPVHwjYbP758whAsZQBnuyDPtUpAcpCgTZM4vFmU6rbVhZ2aMFvMfz2bz7aFEjUmctVmA
0ByoCQE+XscMk1TbTaxn/xN4cXWxcCSHpLhlcRHMO9ZFVGRalqlKEq7GjakErWzdiAlldKjnhm5h
zsenQ5GnauP4/ZYUF7h9VMnCTxVRTotJMsjREornkBhkd33gHihbuh4z17PvEep0Pp3K8P7F6vz8
F3Hhd/eMf+OEReoETbuaKpZBb5SN9ur1QrxZPpmOjldqfm7floiVTCb+cJH/jfhZB4Bi8lcx/eKY
7OrwC02K9/Z5YVOV6vGfhJoEQ1NMYUwvIYXf7SRNO7rErkXfsPsIvGuSIUbvXGkgdBpZloC3gccn
9EQJa7Oyjk1i9V8G8LEMf56MUnOHZIOahj3fEKtqbDd32DAK32tQyhN9LUQzquyT6RVhI7pol3HQ
Gvs898RcpM/uX2bau52l+7aRplMMeZ98kaq8C0dnuk2stilccp0ntOom2g8s7BTWtSBoHooM02Tm
HiZ6KFaAc3ozEcn7v7M0kr/24cpoqH3Rp3CaJ9zpTBXbUx4+VjqZ4W0Sz6MP/HJJdLmX8by4NSuh
uZJ0uGWu7c6/Ke/1tQKx5aPu2mlNOWaBhnn/g1HJxOfc2CZosuXQamc4fPHuUQfxdDYG/KJ0EvVi
0sn7jAddp+O4X/cuqD+EY+WKbaulCx8CFolD91xpTp9jVT0DTZD80Mb0wxlrV61QeZrTz5iYIWv3
Bcbo7pl5xM+H8uMzaTFNKO2B/lg8JSt6EXObdlVRDZcMQnpu/83dsrsGgry5n6bDc0rVSQLu4y1Y
EzQ43XVkkrxYtJhhJ9lKRqxWC4rNE13dyXd/21ke0T5/n4BsQuc/buRGJvvgbl+TR8IsQ2XYs03c
cqOxMnERhusgcZhUx4g6/25B6D/bRZx2viig2NFRamEnLZ7/+aTcUYf2ucknLHxh5o8ej3o+tkJU
YFuPoCUPBb5bfU+F2LU0wbCHZpQux+IeanuzE2QIpj7bXJ9b5dwAAq79hx9YA0hiSsmbwDnXnV0j
CvSqtgNA/Tu1gkF7o28ZUsmqjgWBiL82kHNiX8s4L0wdNY6mqmWljILN93eSr8ohrmthYlgtdKnZ
X98ixXL/ZjW57Y7B/aDhQQbDxYsVSynMEQm97qFn0dCeuQqbctLfXA+bBZsZRrD5BKKBboQ9zKy7
l9fOxov4m7oJ4Eqiu3605LbYZyoYSAIz2uSDXZBww7VABnNAcVaYG9p4bw25oA5oKZ3KRhg8NB70
1HfUcDXL74O1o2E+XOblJQd7GItgnRkbVG4tP/8rWGgaAvRcITkJm7KQut7z09zPtpV5mSmozbel
YIADaIbaTXbzFpUEsmqD3DgM0e5IXaXYArTNPnrl5Rkof3/FhCG/kk+K80sajoS9/KCr/pcidKdS
t3NhVJNxyzauw8/rgZ6TZ+yxhVWqToRxCcWCbJ5d/FZBwt0srSlAiSV/Eb/3nY0KuAmWSQJHc/1b
rspxe47aodgFR/8cMtOrHuYTNH2vqLpkDxiNmHL2G+ZXCAaD7lAoW9mvyk5msVCOEbFuNVj8dQPR
My7Eq5Hv3WWsErnunKXx3uoiB5MHsp1cB2PKhZ1LUhBvu1aX+VLmdcY9V95NYVzzR/kMX1akO7Xc
RLuc9ZbwmFqhfpytIrbBUYzrZh4xqrdQK4url68f8IHv0V2zFWU4kb1lzzmiKkXMoJrkqpaVUoRK
PH5lAOYin2pjomTcIuXZnsGMNGT232bYsqiTjCWbLmkzx4+UJ/3d8R0023E+ToQEFJjT5LFALPEA
pL/4/VGkMQugCU6CyE6tY8pE4345M2+r3s7C5pUXXnFSY8mjZsmuRntXVjrnvJr6/Alpo8KENMmF
KDX5BtYDEnQ2zxjRWIimk7tOx4PoAMEy78Qs4oJ4ZxPplk1A0bSTc4FoRMRjUC74gd3SFUZg6ZqC
Vj1VgUQyucLWpiN/10Ikf4dSN8TuYOEOxZ4j0dRMJOdhMVl/PLqETKYPsNoFJjPBQqCFiPlKiIbI
F8F6yfqUgmRQEe5I7HQLnDgmcYdSn5yKJlOgcp7FABJarvNOe5ZtmY2IPzxYn27nm3x/1qFDHYdZ
w2m1a1S49eQz4885EJyMnLEAQb/xz0FMvJxvV6bAthNrdXIIJC80ZhCS3IP75agQSzJLWmK+eWnu
Ng9w8pRPJD3jPMLejpVfV7Pf6rQhcLDGl8LQwCM/fDRKA15SCi9awcYF2pnSAtU+09bXhUmI8pIp
t4N7JkVLetfronQLekiVB/fR+y2fJDmhzItgU+l6JI5iAP2uOjnUpW4qBvOuKJMYSI/eIpm3ZXN1
TlAr4OOw0kDxzDFczSwzaARzVK73ZHUzfY7uRtOpDe8OmWeHsxG6RVyrAqS/eSs87jbrlA0ict/P
i/ctNChZj7mDBJlMmtESyh3Oig6IovrMFpZ72mb39rznhivXy6aC/TTvtSFwHsx4DWKd802jPMjs
DDiOsKpECUDc8Sw8efbTh1VPA+Vu1qlGxyMDj+DcUTtl+8pknrKsXcV18u+chIO6vJMWxo8jYOpv
0LCsfpDYbZ7aqME/Er92+hvZ88kHESzc0rCmaW4x5lJ/gAbqBw3KDQmQvy2kr4PH9N27H3HT9CW0
IR8QsggpjeSx9Xt7YMlC1C0jUQVVhmcaS1VfxzxOeMCIvN7jA3A7sGYXxGIwt/6/mXTk3zE+kOr+
uyNwwfdiwKy2CAHbvUH3Www4r/RuePk6ChgixH+hMEOOvTMTcZBRXPFiwOC5alQLv4Foz2cNrD97
5b0SOSgjvgShTaXde+h+JaXaC3fZozXdD99hZyzDn+Xg09JD0HtY/o0yLtZUWI5xasB9mdpSti1X
WY2os/4eoVpxgy8sl1f8g0NzFLMFjWdWIUMGPvdtVCG5wfGU4GfAS9YHscaBv5oRs7lxzfhMbLl4
3YfZ0wZ8BE9hVhqGxI5zEnGM5UF2l81MRl66R4XsPkBJZjq6wFhMsjSTXKxgSwoQ5xMfDT6iE5fM
SXWZxmeCK6YvkZfR24lSC4feEs87wykfwyQcrN5QEx9QogSUHgJEeN8S2Sn3eyZLqrKLhVFJxnsJ
nESZaEwWM3jhepB7nSJ7wRKpfgZFoeqdJCx4Dxhu9b95XZyMNMbFanF44XYWrUFIiMxLhdTB0OPm
xuD4bhJmg2hQqT/HGLPZ2rmcZ2reZ2Blvyq0diQbKNh2uTwPTru9vwnJuzSwRh1cAu11GNp5ppeO
zPh6NQjDTTejLPVAu5RjS6roVq9zinORwQ1gd6gCbBpsk+76B6JaXwV+qKcqVPlIvW2DuzoGNZC+
HK9GUSllxrRFv35inwRuAF6iajXySZGZZvYn7QKYeEegPThkrUKJCDXS8PJ7VYZjg8nzqweoC2OX
epwOrFgIRedggXCSjumkbVN2jZ505jag8WdalfNBb1ayfPynwGq+YRTKALL+TaMT1F11UhdhDcoI
Tv2dFwsiV2sZICPhYLWUkJSnNeQh7b4KR6dhfDPnaQI3TIem422yb6q21tGamUNYVG7Y9Lqw4tIa
9AccgocYKSg1dBrLdqMyeTZnE1TeOBWP/N+87o8otmZd7UH2M1+CWG+kX4dorxETxkhPE4vDCMNF
6cIQYwX1TXLmH721DLaxlyC6HneHJ9ut3IAzgAIHe4FA9E3/JVbninHHPF9hjpHOC3pM9kkJ4eFH
mSHxmUdeR8B0Rnvo+1LxUcgmVJxxO2+fkaZOOp8w89UoecmeitWyjWqico/9n0MqE2XNVB4PwJKW
6XbGUUEBpq6W6XD7XsnKgYMayF0JN/S6NDozh57zD8/LSEnV5FsJ1BhEiaSmgibeleRuq4cnH5EX
DsERaEiM254ei3uimGXepklpWpr7po+Dxs6mV+Ef+GiFsd5KTkwxPFAJRP/7AOnEHDajcghTZjyI
nzkZcBjRh2lvZmuoHEP8D2r4e87QYkjeUWiStn4EGLSnKAXD+StNIQz7rL72akgHPaEhOaAu2yLN
pu70CfGyyYdvSsoUPytPGBTc1HfMTTGG9TQ6ZVxzXK3KUActT4DimzoZqBVej9TpPuyN2MEEQ4JM
kB/z0H83DOgzpfKlZbM0voKA/0S+Q9XjYWvwhuIc3D1iN7KiNQ+WNLNndv9fwPAWl+DEdbh17bSz
4QYFxEqIML1K23M1yp1utvGfMwxH0CdOQGVFupUu8Ali/Hc+r2H9yGYrIF78xa1AlGiOU0LamzRx
iCwcBvz6ElseRd/4KrOmp9SccsddxODmz8WOQVAHYdJEs6msm+G2y3Iigs2ZQ9iHdK7t1WACb4ma
eYrt5IJ57d4P7KoDFSqDbkdz36IYLC1FhcdzjA0QMZuzQwRHi3Cjp4EcPVI67kGdYNDDeWOhg8n2
VOKUKkw31XCjM7ygkUcL2gGSqtxOJL09e6LA4QyVWAomHkVmxq+5IB6toHIDJHieLE005th/MtNo
HTMkW4ZnVCtsmORVQUjyLh368cw3IBL7Nqyg0rTSxge7o9HvJ1xdS6NR+JVQHWxbgBTe0dvTj77k
wY54coDCi/3rko1UGBkIaM9ULD4rlG09T4gclecTCwKMkG+29mC2dMVd/D6+pmCVhXNpJgx+Qevy
ou4JPAXPJR6ZRHUghw4ErOjOl1IXAtdQmQ1h6LWxQ2axQe61H13LSrXcQY+WEvWCLcQ17hTq50WL
md4BAQNIPBi6vqfPEacx0f0Bz8NcoblFf4ykgTHHgQYxst5+nHYjGYGGDPOCMC1SZUmiapTA9gfJ
Z3STbN/YhU7SImm+6zl0j1JoOT616LScrFM2zh3vNKTID1L9djjWkbeSCrBzNvUMUu+mvaBFiojY
/w7YYsQbJ3Wme1slZ5fqBPQme3I/wxwqu8lcYoLIrNX0DNn35rhQd6vMY+8sLIL//pjiYyGvBZjl
5frizqA+VfxXQIMwz+dyft/fFZtee5QjrLa+LitRAQpZLo4IXIMkGLM/tqN5C52NIGzcFO63tIJx
xLCrEFPaIHgFLVkYU6ooEb/UlubxIQMxJyLJHkvzLN8rPsRYVWJ5Wen5yEcI/IJjndOxUo7FdNVE
iPNuqDWuaISvf+x+zWoSWf6mNep/QEzU5Svfz92Y/yk+OXJ7Ysdi9u9LyIwLv8OEA5LVORImwpNi
R/N6z5UvobzOJbFkjS6E4nxAleWFTOEBi/veVHRuSZlDcwicPwg+vPqNAPpCcULdJ1vbho6CJSJ9
3rheypJPvbF4kVINJPfooOu1rQsvr8EQtlgy+CyNWFD48TXcR9RjWYmc5bpMQe0qGreqa0OayDG3
jQwDw7ShWrho6ujn9ucx6Al3p9xFDiKsBJfo/tHwz5eu/mL51UkX2qiRZ4PF2+JdFFNYVlfnhfua
5Ke4IG2K9NYKv4J6e1Nsekp+2hNlWB03H/r+x/rW8jx6KwZgHGIYYu3yY8A/cOyDQayy0/FLYYCw
vXqTaTUc00hPzH8zBfhk5Zk2A03aymHGdpvTzFNxsACvOnrdfa9L+etNEgnb5u6YDbNbECIjNix2
w0wYvhqltq/SVZ43gmAn1AeNytxVicLNiZb7G04R+v3Grl1TZX/bzghoXZODE8FVdWND/vJnoKkm
jTCeBlOn/S9k21pv9/Apc3aH2MZHAHPeKb5kMIPsYfupYAY4oIehjoAguQVoWpkN9lxv65I+JVx6
3fA/CuZA8IvciWf7Ad2GjHRZx7EaFy298m8EqDEt9jTVTx7QWeQ2I3goYOZmP6nxvueHmtBy1etD
+90XDUuHcOx+NTXu4HXlMSe/7g8Xgkqon+bnMeocHMUHNB64ekbCfoGLQh8alU2THt/eTdXTeJM2
Goount56fTXOQbbiSnVKrl0n9tG2vM+T3SPQbDKC0cwGogESPI7U0M1VRVMkhZtpxnY8XjmaVYpF
+Ii16++A10CDqMUFIpwH5XFu+gNRBLemsriv6SqX+OFzEzLbyRHvFvOjn6KO+SeTWN6/Ff5z6der
i9n8xIKC7lz5e9UNQxebQdFI2GT8BFWqiiuVThONLifynV0bvfOwKcjq1U1ePJiOYBhbV6toB0PA
+UdIHgq6W+BmrBDaIPFofnUxwgVue5eKZzkI+vrHpdpxSESu1MWLTwaNJhnKpYRZxDyhJ0HTsu4J
qOPlJRENmscINH3bfqfJ58ZSYW4PydE/4kpCVORELQtnKmTaa5n8vyasJ3teIwOd4N3tZL8Zz2b1
20Rydw1o3WjCkBhgJIOTolDR29VejzjI9+ceEEeMjPpOGnyN10Csqhn2kg/sMl/rHnWnrLdLEmAt
I2YzZJta7mRV4a2iq8ndVOEdtDVjIBV8SisPTbMzBVrrOJXD592o4ABL17JEOWEzt6V6tlYS9/96
SoylPBJsbrZuu1cizj7aezQIc/eH8n8H3eGRFeyBVjSTg6eKhDX+Gqs2qNPb958kp2OUPGr8pJ07
0C2H6/AZeGyNqZA4YTl503GCLNMhs6eK+kmv5vvehHY5YyWQ2OgY7OQu/FSrIEE9TLbZbOSb2ckX
227qNfp1fMuxnT5+pMczRkYtw/vqZH872VlK9hpWNJ2yRy/6FaCsIE/Tm4h5biwMD8tWZIto+JOK
YpjWV9y60sTM1bZHVGlEh2/CS1hkwtRIhLWFAq5yO2IO7gDrxPPRWiEMcVubhSgOxVhN+H1x/oTS
ERDFhiWbz9M+A6Cah9RLu75ken2b5/Zqd6gznxYuM5kBp9aVxcF6s8Icr5t6ab1z2eCvDhVw1IgG
i5uDKq+cs3D8f6jtCewa1Ocz1HQjyokP9gtlYnfBxfg/vGGZNuXIct6Md8sly4mrf0zeN6JZwgU5
blO7tPHpLqkEeZ1DRw0LykZ2qhVyl3ix8J30DtsK8wcrsXfqs5J4EQwgYnpAMV8LFK+NjnDgDNaS
EWbVpCc1kzMZBEFRiJ6WKC+DdtB2K0z9yPPCAab3rh2wC5R/P0pIEcHsgzMc/NsXVChXHFnwnbTX
vxS0JuYZdNH//ANDqvYhawpsCt843PmgnTqKYVmvbUKdcEtzV2B+t/LAPcAig/E067wu+c9rqvIE
Ck77JRqlNnEsWbarHR014lY2KLy3HxNEzbMdnJEQMB9UbibePNJL0DhYP1FEW/jGA44UsKyiJ7Bb
8S0wNO8HKyTsA2/fhUXJUc7BUnnndtbRG0CeL6BSc4lhy2jOoxQgHaHv8yB/dpZddYvm4yW9VuXi
9F2yxDnIkm9hqgKKXDZ9IabRZQ/h91lxsaIy5ufCnyn6N3W0+C/m1FonZEJo28/AKCrh4RJMCaws
ZChC3SXTcygUh5JeCqYGGV5j0w0VzC1D/yV2BD4PrwdD1NXK/wVRxikeEXCERO60obsM7B02DxAN
bEUIfWgzSHLFvOJdUZ1z/v8di40nXCAF1xhJQ18QoFMsS2BPHHeUFdZ3g95s+j0DlhsSyRmD+QBB
1CkoqK/8M3WubPhpWqSD6xdQjlxrGXVvTkUPFym9q49n4/IazeRQMYNGX+GjSoLBDT+wEdLJ/7zG
UOiwI/a8e81OPOisZ9bQmKQpja8w+J3Fr1fqxc0mJPmjTj7SxSaFqzN0RTeqojt0j/42SFnkgSex
vgw9X0qjl4MKukm3porXMrTJquL7iVIQvwGtHy+Odw5Yg47461iO/yCvi6DMjiOMXF3Hu2gxm5//
ayAYwvTZkwNJm1dtZLfoL1/Tttq50gxPM+Q5dR8CrDRq1WiDQOjSZ0D6rWiKYLAm11iKcG5hfOM+
uKIPXpfKTrIiVp+a48xZ0bNjFw+thDN3gXcSQhXggDI15b1hlDvgM7JcktaTUYAiL8L1b9BtVqZz
95PIz79rNDa90/UXhegtKqm21fbL0v1mlSFSzyErO9FqtE8mFa0EL5JgdhsMrjE13bcDCnxlf3+X
f6ui64A5De4GCxSkRmL+N6SLAIu78f9q7ug5erTTLjpW6Lm9pQUVklJ8DPhknCqSoZW+/uoJFECL
C1Dr7AwTwV2JW7Z5dsewqaUpDs8MN63TUpae9Pv7aqjG/I+nCV4mljMw4g1fhZeHD85zaZ6jl9aQ
Nde9HkdTq/47sZf7m7k3TR/hsBy252Vw42p86YENXoEOPKBFWA12IlLQZRWewO/xhbXYfbk4Sad8
2NHgX95rKGtvFA2bog948H6J1dNsp/MLfGghNSKFAtOu5MqIEwFbvSUZRwYjgz+oTRJ7MKWr+vpD
rO3o7TLRV+TjFMOZV+mycGWOkF3AB25pppTpw28+M80yx/WimiyWqpk0Pn8gnr9xvEQlEuMF6uMv
h1BZajHcMzVRVRDDaKAOXYvSU029c6Ed2tOLBgcVYTkgUNzfaIq+5HyAbqPnkAu9MewVkV1qCyVg
6xJzbaAz3j8p5XfK602So1y1B7r879QR3C/r6Eq5cWHF3tjpcKYw0sPI4GuNqMnvIhJgkD3tM+ec
KcldL7wikD87mk1s2LTnZDyOg4+6hvbxHiiT//WdHbTnGptIoKX8c1zwEQ23xJQJ4cWJOocd3PEw
xmEF7VLeKhePjtWfH52oaSPROo1GziUyWqGv49dnUI3HBDPgil3RwewWFbeZ3DOLPCO51IZWBAG0
VtQr63fe4JXPq8Y6ZVozUI26RaaIkmS0sweGxrq5rD1UKJrgQncBXobbv6/ynnTCWg93jjzrbllv
ImGbkjGfbXB5Lr6fmioXcUQe++ihgFLzl54D8XXGXw1SBQnctJKydzyQaRaZshMSbHETA3lNwRO7
oLiAfKti0OCVSVz6+3J6dFo87YmOvfvaR8Jdun2NxE9TmUvKaSyqEoRsyyBh9HfjkIzX0QSAi+/Y
CKOqxiRepJp6uGyui5b5EhFH2Gb3S6rj5WUyAoyMEo6n3pYolC52+iUII4Ix4KgMASVTLzbtIFNV
YsZDGqCPlLnreP482ishbfeJ13tUNJPInWes8yHcASeaDHDsrWCWcVgApEC51NQwFR7Lz039jSRN
bc/Notq6kWaaN6VEko24y6Zb1xXroi3jXwmSwC2QnS5DpiNJkzJP/9l9wkvXZrp6jSQtnilS/cq3
2a4jyXBl6LW8s4t34VhEF+2C/lldGoQaHgiUj1aQ6hxhDc/e2QhxzUAPqhDYj+u7MMGjUwLYk7X4
7VzIX8sgwbeU0BntAZJJE9UPXpeVtIhWr44l4S0CklkIod2ttEY/T7cTuPQk63J0NDSzhX7JqcTc
yHOGlm2Y8im8ZcUu9M+ecb96G+OhLNM69VqUIHqDIv7e9Nr1tKW6G6kQj5PIQw0Qt8Jl0U+TsVrW
5JtQ6VIlFUKxHSedTjlPXGVQpzv4z/IKdrTmXE821Coi3jEaNtFTKx6mjfYXUSO3JadyfXXlPy7r
dhAbCkUWB+PjY5kO6Ln4KihwZ3gv+FJJmrBLQAAkC3fxIiqBJfEsamnP03RN07HA38Yihd7Ywxwi
FY+HIIMFguUhy9ZuHpaWHHfQF6/FwHjbyb4BMWE//zTqZh/vhUKhqBaa7gA8kDgWcukJ+Sh7XY/w
xM3qkh4MesRHcFwBvcEHOHd47PoYT/e1q6LkQ3Cfk2GJ/AtQQw3s77x8ki1XLnOKl9S+hGW4s0Db
TJmMizLsPjQebOLnDqn0xpF6t2aMyOHhtTwao7vjUsf6NVRctxP6VFk996cgTNIpkNq7EZ3Wqvun
mW7CYtSNYjRj9wzfX8uMSoHNBk+HhZvC+R0T7MDq+AGC4HyltaCGhj78kkXNwh0dYsZHMPo4fPyI
z1Di+Tqw+/gd1ARj0vN/w5fmHgoKnLueq1jhH7276RfXhZUhezgYHdg0OT55pk29xUs/y7g0RSMh
W8pr0cUNo4paZ2UFA7aWVJPFfIHf6+tvrrtBR3e/ttWz8DIfXvzQlW0feJ5vo5ZKm4hiSTDmOuFM
f5FIrzm0E2EQqzNaE0KhkJOsBTxm0iQCJ9NiNFELMeN/xNC0X0XiamThIVHqAQidJ0FnUJgGjB05
H6TG24djNwdU7LpNW6pIIcrVtpi8Bx8FxxVpa6KQts0jMhSzD5YRRtHTJFkeDPb2g+sry3i+gOU9
ujGEanXYFkE9qUqsC1v2QCEKksMpIX8+V2wv1cIufaaMS0gegFd6psP7enSLzL9AWAhMGCFhQ5cO
G+YF6TxlqWJAqqpBEmoFGfgEVRzxxKeblQrdH9q82rLBXHyQsJTrFoWMa153kscLJbuGNgnFIIvd
U35HD19VjfSZoTxih/xnNvC7aLItLz0saFsFjjkeDwUFQd5KchcmX7HI5fFuj6TSQQC0pTudWDx7
D/wHg/LHhgpDPtvUe+lAkMxXuKz8XHa6nNxAut78sbQ6PCRgyDYalKLO34r33J/cLif8CXfGq/9w
w5tboETf0dB5c95ecov7Qu8gVl6YLhyJVZF/OFt8GQnni14K0GGgVgtKwVhVKtmJXyeOcPakFQPq
33rHhAD6c4CYaYDx5KqCjjlA1SSS62Rjp/8NyjFWKpdhO0KOxbWIN0a7HmVuglRQMk/7/+I1K0Nj
qrCpB01DGTLlXRCdAHrmfJiEca7F3RD8gp1A+mcgqi2XIz3Hlx+NSVfwbdM8++D7zQ1hZIfL97Kx
kqgnxC/PikyGj6q40ilsybKu/OLRJEHudzdIAKhSF9xjhRjK7OoL9w86t/g5uPw/R5Prevl6fsYp
8yWDL8SCDBLn+G78ZQgcc1YmJHogCPgcJuh92Wgp/uOjynuuI/cgPf4iFaS+kqsX64gj5HIzqvhw
fKAnmWYJJkUjXxHh3GHNTqMUTh6LKGtCbTccxoWzD/2x4kl3g5H7fsrTA3TamHZQy3wVJBh57UN1
LWVGuWLZ82xaAGYjaOyVvlSHZUm3nzLzS27fhoxnMjSTLsJN3Qb2duIl3mVQNcgB3TnE5G0nd8/d
ZAnAz8Ip7G5ED6ZR1VjHMOJ9IDhZ4wNUTjJk3fihWENNEaDGhqVP8SS24m8TbX1jgPsswqLtlABc
t4synQ79krqpKjucRwvFh+a6ZRp9cYUmGUgxMxZNN6mUTujM3H713Zrl5FVQk3ec7Q2ZoCf0yv0p
gOhF/BBrUE2xwmvbkfiq+scn1y0qss32PspWvPnWNLYuh4aCgsuyO4uY/EsjhiFVrQO0EGrqVwmi
CPCMIx4gRwXjfW2l9P7HypwqdzKczQBO6Cpve1Ok0GVatMALIwQtLujf1CSERep4RUstHCJWKQSJ
/asy6n/+u1DzxP+f4aw9psPCGHoDzZoz1JV5jBcyalxaUUdol67wkeqd2fALdqAxqrEQLgMmIE3k
RC1cmMJROczyU02YIQIHkLzM8gfAgL/EuEfaalNnWKHuEK3NdcFUdQ0J/Euli7KuAtcIlv8/Oau8
ubdmOxdQSDIfd1TApp2Zz+oqbfPXaU/qseXTlgQyNLrts/4DCOgJJtmZ1kIPNRPb34rdfLPCv+fY
ab+Wwf4lDIEg6uEJOLFaM8VEOi0QT27QqwEfHsVSbf3KoCLcmVElpXiJVWaAEx9is6q2ev09/jT9
cEpvaRtWu7VqVCabwCPz6uZh81nD3lxdR6r6AQnqDv9kbykF8QFE21t8qKRoj51CumeWTZxIrAwV
/JYjP7hLhAHMuF6v1l9MN4JRj4hkKZRD0nUKuiC65XY5Iqgan2gqJulZqOXmPvXbtYVuUoSPmlP7
zl2PYj2VK3++q9BxvDd6EDDF9PgOfabn7j3M+hxwjTejQJpyiC3Ja7OgolEqC/6tZ8gVdkbkQM63
IiCKduuOdIdaiFDB3vMI26PXyKy7C5b+GeHweCTJuYB/V2iinSeQr9xiH9YaKHrmTJgNowbDbVdZ
/vh08s2C9o4stZ/P2xbS7tQSWxRmDK7VAmMk/BfvYCbnKa262/vcAW84gVWzEGgQso3DFZfmeVOU
FkVIv95YyRyxIzgA6r6/PBluqL3PLPwvK6wNR6ix4EGzmOnihK1884XSzYQEYBq+ClU6jqhIXH/c
/cgW0zGcuz9c3A2Jwmivu/MH0/a2UTkDfSUltpQFCLGUF9aYr3LAdxi0rwwsiEOFzRVW/AL8pwa8
XrWKVETC2Lf2S/dZ7JLGdVuer0++Q/2KNbDwzGDMBTEODbC+45JkNWslCjjAyMZEOt0T9+Wi5Yhd
uTULHjnl/6ofZ2sBI5TwgK5ShthlND/Mwa2hWlYbsJ5EivssFrsxPgo4tMRJJUvrz+keqN8+AIJc
AwrGaxENEwAKQz6E1LSCbBLoDemimi6KGYWgkp4CFoVGtPswWMR6Q89ywxUvZc8dUD6jb6bV0FI2
cWEu2J4PuoS0Izb/moAtCWwdIhc1H+LHuVyE/WTO7KBESGVEqG2lyulm3Iiq9t8ymRXGAoCE+raF
OxCYbkC99aIJ/BA5LmR1wUSNLjagyUGVsv+PvicX7RTQJjbC3kY0ABNHiCm0pPiuGvDm6WJ7ikYQ
jRKvXhqFJIuBWCJBeVnN9qETyGCL2IRQWX0NZMATRPTew7CtnQRJWUPjcYRPjM3l5NTifJrwvw4D
sSlxUmWqHmC9ECuaUpv0g4Gn+cDDIIglZAZNbJXYCtau5xLCXTIRApURWZq4WgAyhQ8xX5hPhQbf
QG2RaNxGhOSmDmWHizguMtn3UCtT6M4mz953B0+WigkqtOd/Qz3TE5KYqiq+EIE19l+aTi+ftIGr
FPRyjgOwgAOkqmpkdkKf2rhTzfGnauMZAwmrV8VvqFziuVCacmIBZQzLt7rp7yF+pYr7Q8mOhb6g
/g++9BDnpdtqwqKQkgiHgbMaOTmfqIkDpfNGQuUSTPtwhCoynk6v9ImAsonvvzK4Z3pC1dh0CDB6
Y1WlrrISOmPgVUPJXRMOj8OM8EHZg1cfwvyxBaGtW1Z5amgosuLqF7q8B8fxG8wAt8O6IE9KDnV3
3X2TVk5BwlFpeXv7WX3UicwJHKVHadxGCXw/cNrgVrbNMrY2g+RhumuLi+86E29WGBcz9mSSQX86
EGI8vn8Ngk++SHLvBOZAFL5oa/t7/xj/jv61OL0wS7SC13bIl9Udoir34JGaoDa0HsErF4Zf0skg
qeau4ExUiti1LfKsMbzH1joSyfEYvOlhPOUOYiL6LUaJm8Pu/mCjL8joxs8VW1aBxxMIEvCz/eec
CWvxofg/WP1aIe9jr3hVivAKALuoNrqOMoX19QUuc/JvKyF2xfXUbC6SFMqrEMqhZSMZkHowNvtr
ErqFwl3hzHZ2dVHs6g6KCqHu/z4n/epLT/oJDjYMBW4+KBGevEdDKWVsfqT4h463FAXjFG2wet68
DgO1xGMX13JV1GcWqULvTPGbx5mnMiGc0/ngCTxHTnkNl29P6QihGsgEf41ETRZFlvOaFWyFBeXV
oI8pN9v2/0muPIi60ku9GkI4y2Hqqi4NamGwe2/4aUuBhRQOQM30Tz0z8D5x/tirSOc7aswQgZBT
6gyai1mwNWfvrOHZzxE/XabmIOYy3jbn1lrzO9MNTMOfWJusdWAVNvw9oUtmTHu8O3hhzzlpOgu/
wz+DzLgDu9pC+8/1VsWkAsiG5/e9/cknkaPkzl/I9uzaw/5wYbgH2KN/JL9MbFMIGn5pKVSJhnCu
JZXftfcLSnOVx4aauGVs0PWw2RE6usa3c8uLr63ShNzgZ83Mfcy2I6q8BRxiJoKnnHnpDLyMpip9
Hl0ss7B+CKumpICjbvt539Kj+mLnEhS/TdC1wAYDj4isjqvQ5iIw+EyNzb3CZ0O5Jw9ZqL5GZWGB
OcIruFEwnr3DK0S99rNrz4jNdx35ZvuWxqYyjdRAoD0/iFc5wWpSgTCPSq7jgQt3RzmJEe3ewRiY
pbdAKQlISU2KjMhHu/Y8XawKUU1pEWbZn+aKGLBtCqumcmKiIl2E3m1QiwwyaoWvLjSeJiW9S0YL
LtXhjFU8N+M/86j5DgW3YBIivGcia7Y7hl+v1eDVlCKrtUMemLa39skkWHAU56vZvzrCHqZNbsUn
7JUw296f1CbszAgMUkCVOoA370bM/hpEHmpzas+JVmkMkWgYQ+R63md/SevEpLmGB0+jX2pFNSR3
qXBti0PmNTXPPn+AmtOv9B0HBkK7qxm4KyWGAw8Jqky9Hv1OiuU2ks3uFw1/pVaOdaP28Sav2Gtu
jUMIguDhM4pt2FzGSIt3iFIktc41iU/rCKmrDL8GuwYos6LCY93GhBYmuCme+uh7wSKze13LPero
XJrDYryPRKiOy3vPhX3PMjhhxNIKf7JVRMTClUwhn1AIWHjtUcUnW1TXoTEmpbITb9yyLR4k2w0I
Q2PTARjvghybwXO0h8/T9Leycy8yJho+YBFx6ohJuVGGkmQDJA5w0HgQkzfE2pbz0Buv8lLI7f9s
+0kriyGx0QLoUIaH7sgebDBMCxQn0LsGudzcTCNZTheYkBuDeRWHizIidXbJC4ZBhzn4S7R2yvTw
W+qQGRlHNwBLcyaw/2jugLre8AhY3ICZNwFanrvsYQN2ViErSkX5E+E19T84UCr191TGmlXMdwV3
xrHY7kycRLZeGelZyqocjgFmSMkUiHqEHLqwqyJd7HOd6itUol5sivfM+GLWFnwLlFdRKTB7feMR
lhKf1bLbXrWgWT5O/uvf9d9KJhWifSCUS3irhQLquvrdxxw9qlT2AUv787ByXvbfuT9kabf2edB5
DvbI43ParNxFC2+h6PoSDjnz5zIY7jiivCd23tJvmoZfaH1U6OqBkvHVCu/EHRPgb9MFi1Cj1wY3
l6xwmL9ER58QJ9LtuKu+GsY0L32dBWZEk05dLfNPC+dIe45MVIs9Oi3OnmZu887L4WTXQsqlZIxp
/KfhsPh8dfybY3c30zd5vVm7ahgBdaWZg0xAlxJw1XcrmpnCZRaKQI4NTqUaAcS7YuJRcumSeyUu
KxfycBWJyXmoRsFBsFbthJQ1xvBpmFKOqZOijzbQRh5eV2kUIOfwrZ8BZkOpqAmgiQcdGFo69DXx
xE2zdSs0dTnDuaXZKfLWn+zD40idofIKD0WlhxCJP1SQKr51Hv1wBgTbJcJj1Gp60dIphOyZsQPZ
2Ct1916zbMVVTeDsUrIfp3ahvpOfqlYSP1wSykp7LGTotGE2a8V2Rpgac0TsC4Aws8HFgNbWZYbS
tNKvGtK8quv08egM6K+FlwhIEXLye7qU8LxFnkcR+Dej4HJkF4zkPhxoT1j5jqnkKJEHZ1k0OaXZ
1pAKGZbbMu26amCVrBDyby13tPzDR5dEyvejR0VLs+6bGsWHtGHG5onFzUNrZAQPEDoy4+6pTwf+
WFOwGXqWmkiYd12ufjM1Jh4Y85qhnsOrwiM+c4g8Su+ev3JDfR8QlAumEeJptUQfYsiYhCQLGFZy
9mWbU5baTk+v3/Sutwi0ltX+MneQaSVs4bdhPnLZsOR7lzuLR552BtUFpeGzD078W4PfsO4Y91qK
UoE9GPHu/o2XeoTZ17M8fAUuSUaAyEPFG5QH3SdCIUQqMhwIldzm60QYY/pQeTRGOfzbyRDbQ8fu
Wr0zVXaByE2nzPFqBVF/z7KVZ9ZmSfZkXhOMscKwcIdXJuOViOBe9SOT+GjGPvr0bTdWCsUH2JDq
w2qPgFa3t43U7Cm/GHWUu/mBMGKsICuReJnEr0dawh0ebiQzPAl5oxq9YisscC7Da7LtdhIRHan/
gqbVkSRorMZQTgQiU0G1qSlPmcRtzC0QmSoa0pbJEPw41KJOtuELk3zrz38DuqwZcFpuVTckQXGi
kqpNuOtlOWuH8JZz1jbhJlsLTcRATSIxQkXtqkn2IcKMcNUFKmpVecHvbZyXpAFJvpSjkKxI5BY3
Cqlnk77rH3K4630njQkvGIkdnEdZX/Lp6avuYr9HG3IZ/ZQne8zsNDMioJnRT2amqtYi+rHixN7K
sAcpxLjBrM9H6FT0kQeMX226mi3n3BXMwrNeasfdaphb8qABbuib9aPn2fP27gAmri8LiAMRn4mo
kq7suo0MwIzM/xs7W09qIOjgSqb5HagSAw6JKM2eKdaAG7FTz1uIkIBXkLmQzf8FpF0x43tNMwzD
qBThEh4gf7/wi9jmmZHDr7MxrrYCeE1xi7U9sVYzI++aVsDHCPNZlEShG8wKoaA1pqjXBesZ4Klt
scvgya4KOsqrs6QYJFffkm8Bg61sPGZVVuoWYV3VgFRC2Cu3gvhQNR1bFeE1L8rviUdN9cODAyFg
uPi7sCDX8pUs9rGYl/kq4wShAw81e/1ZxE9Ki/6+UxcARX6qSqYQXW8gV/JTmuy1l8btuciDF51g
JB1z67X1XinbEvtOL/9HRQEkRPGYRKt5Lj6Z7qKjICqNzVOnwpHGwR6+WEx9OUWqBT59AM7dt0QZ
1xUjqQvpatt+VxFuQ5AeuMgnjHntStdfo93fhuR4MsTrp0jH3aPb4mUnKfvIdp+z7+96p8ulkRxY
cDIUl8NEk8eZmVY86l0zQHcXFedkp7+HrdGaW+CyI+tv64rcf7zJcg8YvF2M9Rlmjbd6SK609J0l
c+myzfghLZkA8/+Jc6IvowE55jBqJDu6+JW4xTviUx9Z/HYxSCkEUiiInPAsX2fPKaeHFYGMGrcg
DUYx7h/5kCANBuo4MHwEbONaWPaNaXkGcy3bH+9isLYjAWLkGmR5GwWHBkJsfjhPFNBlpfewTrKN
92oipUzHt9p1tQVqlXoIkuGtmJSLvyXxMhmfZ+uyF8uP4tnZOJt+D8YvWoNP2JTYeTo+oIT5Gp4p
A2LJ8HhC0s9wt6Bcl81uQOgC465ZzejADOKtZtOKgKvCPNay/ZBIRG6oVv/rpqmAlvFvIyPMoMjm
vzfWZ3OzkPxpCnwBBBHfTSug/LeDsjPHnwmoBtWq+Njm72g46C/dVAisMn7rSVpEj13GWcc7Ftx+
yexlFWCQtOnwnIN00xy1CYSEK7olZtkfM47fdV76pzt+sofimPsyIsFYNQkfP1+AhIZW7ZWpk6QP
Somt4pS69mS1fv8RnEcqd4vg7K0J0fq4h/GXa3cQDj5JAUbR4JDvVtFkKbSNzKScaardc3Dj+oyF
A4wqitNtBnfVVHMUfQqbwDuElUzFMiXfsELRjiNEu+SCC57rhypjdt2XvV1Tbt+l6EBgl0tihs4M
c0e70wGrfmY4dtU2kiigmet6qfY4edBTaZS0T8dr6ii4Kr5bM+1WEdMhxg1metqm49+1aUsQYvCM
rHHkwu/AqU2ANWdsq8YpjDsIy20y66nE0fIHRw6GOWZcAVV9YFCVJEO+wkJdIyWk82IxeFspB9o+
mMEMczAIUObZhUdQG0xU+h6m2y1PpSOOjcuk1sF50KeJ9aFm7yUdKiUAvMcn3m4t7lPGX5ocLnMw
E7fUUv0gvS3/7h8ETKGL3Q+IEqZxi+oJE8DK7dk5noZcrBqO/qblPJ7o8IeuidO4O0gy6jeQ8Anc
2Md0Lhw69zQoyLobvfvu1laJmvUEJ0XaBGwtab9eocf1O9zMV8jMGWKpXrgbHf7VPBf6QVpb2lBT
rWqTOf6LobZtjjptFjVQJK07jgfN7WpSN+5ol0yODQFJeYKmOXGfm1DaCi3C+0Pmtr3XBUtpuj+e
3BqgUHfZBW61RAbty3cRvGQV9iigHN+g96WFBfwt8luZv3mgiefPotMPvSDiSwDF11i57uve2IsU
ID1jRPLm91v0UkCFQPYjUHkAX4qbanWATkU307WJUNor9nW6y9RGFBbfynFIUDKpUrdWv56AkS83
KkWoFsyLEx73esS/MP6siDElLOUlN726GJZEVymfsxb3kQOvL1o+9PR/qZkdWCeKaD0v6qROSgBy
e7DZfssGUGSowCOgDDvXnAJOEGhIKKV4W26C4HiR2w6DLtmC+kMbxMNI3B/ADAXdY2inB1TA3OOP
E2/zn5W1vA64YxdnazTrw5SgPgzMy2U1ImZVYlamLBvkaSJR+AdHcfYSzqWCWpW0nh/RicaaVmEK
lBoKYgT8RemVJPJ5tvns2OQUHU50RFEMEQpO2spWbsVUrtnZLynJg10k/Utl1TzfOymnu2pXibcG
uJzbgPlMsmfUdSrxuVnKEjW1D5QoReir1k07rASJ8cauKDqvsLdYYjC3l/qbFN74TSoo4PC4vxYv
RP6NPkEFx24PWfTPYvGvj8J4Bk+pLCm0wfdhlPCHudW8I3Q1Ccl5lb4S9Bfa9kxN1dZkix2mOx+e
cyNBgqo21CqZ56p4Hgnl3wcwC+b+AVzhkf1x6J7QM+ev42v8/56Ig3IqzMENXXuGuNLHgxvYAnUF
vR/2RzzKk5lkyCdiapJn0Qi9BULak8646OxGM6W7IMWff0X1pivSozIoesZEwZgPzaphJ0f4YrwI
CfL98AzrHKZ6mCv7FvfvgJmPGiKSLOMZj03dYqiWX8c3Yc7/xE8lmTyL8IzlG4P9GRCUYMSOttmE
yaZ4sozeyeqTKYnHQS1XE0W0l4qBj7Nqx1q8VFq/8O2w4ICFGTxZpZTD6aVQPFQaAbCYcN3arnmk
PBwactlqrI6LBpqNfN8jrbmtpKHQqd7rdIPJgi2Gb9TnhsbuiMePCqBoU6kX/CcwUksjXgRRuy1k
FGACWvCJ4vLMRiRQAD/nEOTlGBdcWwyR+SwflH6mJItLIFvuIYdu6u9NycbJOArfXplojy0JjsBX
rl6Cab8oEZPKy+mmK3kOEs3pEUnY5kNRx1reoMsiJWDUtoH+aCEUyusavOiqTpcCT49a171+UUyu
3JRszSKq6hu/fIL9oFceS6NdgMaHiXTufEJT5Fo9mUax6SY/jTHYl3Wk4t3CVuAnjW/PRScdrlUo
oemxzzOJ8TBBdI7oMw8DkU8KHx6+t2LhJYJt2D8wCYWOuwIl9vLd+8Nk+cDx1Ed1VEyDOiXQ5TwJ
kYvLuoI3i3vJzoZ3KRw8KJj9E66t2aW00cUgYltuobqPxsZQDUsNYdEG+YRVLo8RAuaGwlk52Uus
crAU8FX/ROK0sB4DPHMzmI4rzFMOqU4e/bmXfOSihVBZ4Himhebw5SoP1C8eI0iQ08lj6UlEYF5Q
KELu0JzgXDq3QxnNH9fIiyd6vP5NIRorzIY5PRySaB2POcQKJXLsvWbT1rRyU1d2882fjJRQpQep
RMrzzQwn70UPMjWV7Pyg4X53a07O0eE0yNBbYCJFw6TAEDsRVzTv3QVEXb3wriAqmGw45WJxtir1
c1WnhGHjUJSXaRXXW+2fvpY44oa8jcWz6Ptl96jrJFXN8qVuiM9AhPAxdT8nut1Zu5as4yd+RGfr
wdhBsQq276VUK4i4bwk1wjV+NLbc0QNGqgp2RS66vw/tLQXSloWM9App5QFzcRi/GJefezDLMfgT
LcVH+djTDS5Uud+zAHiWQ9QPQHAdJ0Lsxu0Zje1o3KdkcGZfEo9RrWckf5gN/xh++wK5L6qyhOwe
L9louYEdFhWh73tWI3u2SrYp5H5LLUtCa8U9z9xQcdwFEKEN3T/gRvzBAJDC5v6LsRqrSg6+YYlM
soEI+PKzNSBJn0WBm74ShURLDg7dGw2xaq8iUP/NVf3+GBH7BSxgr4jbw4m7L3haHLawJXQwtNNm
XMCw8zdhWNMiCehbmIR6NfcylkmN4fQWAiZQxmEgv9g+G9uhKedCTgOkonUsbaOpeHnze+A8H3w0
HwJd0PetUspMmSkgL5WWJLKSgOJZNv1QAHd4r931kT7o5yTU/Utoth9CF+5bPMPol8wq01+k3vjd
mPmhCIQng7YfphBe8g9kYdM9snTxoXK+wLl9HuPoExG4W1fc0Mm21SxlyrfCnVZOhcBagbu6B3iM
KEc6ura3Je7dHcW3qydU5iASRMNgcCpI4bGej6U87VCLc/FaKBkZ0raww70LydHPIbB+3KbYIb2t
BQaa25+VGNYFmD2GccjWjv/cqAANSQVgVcHI9RsWRe5nndEY8GC4Nce2ZwMn2j4YR4EW/8A4POHu
IjYISgY5kd4yTSixzU1u+VbSJbQ57L4Rzs3KQnrctfkfbLn1NP7g6jCS7j4yWvSHN+SZHZNGg+DX
WpItIZiEQmhX6s9ae34LwsM9mGdKwUeP7U/vTB23RMXwp/Ogk2ak20B1Ezk8OzpK8Mqdfc20xemC
y9zbdiHkkfrS/1eV5ctkIQOvsqNMSlP57DEcp8rrSs45Z1k2iiMCoxGmXPNSJf4vaqDXO/0QrFP2
BgYfVH2xBSeQnqamGi9BnEa3PVdppYrVxBz1btaW+uv8+90Ecuyn4cqUbxtMSpkEDJnAJylO+mCi
zVHWHfucvBrFssxE6n/vlXedbIW48J2v84FF1uDxRu79w2iqlpjiG89OMrMNLOaouNwcHVL/Hupv
WGYxyp0laomZvsK/WN+QBF1mWMDBZly+dCS2phuu8Xsw00YidePITBz4yK5KpZQclkm2/UjmRANs
NDdFFDdjN0pCT1aajXYzlYO9J9gapNge/rWl+f/XNbBiFe8oDv2WQRAwMbqGZbFIBttcz/P8Q8/3
+vn2rzWs9jeSaGSGAJ47Ff34l/gg6OU3EGfvH/DTzoYBDBYA0G1Zx+ipQzER0nd4qaOExvD/3Vi6
GB5mknWIPIx1REjT6H32VVjiCAuUVfVVEH2DBxBEM9ApS5lmGv8RtL2zEUx9T5anxGq0VVaKeHTo
HHEssALpRwyawXQEvUsVf3nIrnIKy/JplB3zhrwTLrSQgKpgR6BDYCHkkfkeVNribCT8dlfyrLzf
7etGunWpoVz9fz5nBX+HhW4K/8aaJP6OgrajJAUnOpOcD/a1QjB5gZnJzvMN1miv9UN/R62brinG
ez86PX2eNs/yrEEusjKgk51BFgB7GNTM9IeOOPGQsTSCz3ImGjS172y6cG4V20n0GNtHYcDYz/Ln
sBl12IUWytE4Ib/iYA0/3el8xvUDfgsWDiOceo8BP9pt4N4zpS1u07XdskLQqNu6WHakiDkWDGjW
jPPkNJuSTi45bCUaXmZ07ZMMYiO9yq41IyElHge3KYy08p5nkB1FPDOLbBYw5egk7E1BWQJYDGH7
6qCXCFX2zHX2mH+IKNIXp36ztLcXfa7M/D512mDtIZ/upoUCkgE1I19q0QhaFpcRNpMoI8vpkiR3
7fLsEIymn99G6zp1OeIpf+mGJPyeUMOmrjYcVKZbVDzqFhjyzdto/O18jci1D8+f6uwzNjjb+yT/
o1cWNVyG0fspq5kesc2CVj1xp4jIYLfGlvXiw3cmPjIuEkJytKx4lTqQvo+iHoXyO3JHJLHcnmt0
tH4cQYbWqgo+y7QtuZC+GGftIRmYLc+Z2mk61utpVc4o4uAd2gsq/UruKo+Io7jP/N7AlJBexV2M
CV6tdbzDhNbNK+SAHcA6oLuoi4wEqzeCj/XqRZ9snJj7hI5L30iIiUI8sdjKwg/8kpnpIhBK/L++
F1CKTpcO2mjL2MLSXiPbsjP3SsShjIsfqre/yxTzZG3G2jMY0KcIwdp4gpTRdnxws+gjxxlOnv2N
hVuFt6OAHf45QP4R03BUavAyjwmpK1DSfDh2+KvngtAjjLI4SMbn3Jk0t07kU8IA/RHTUQ4HPIDz
SYEfFhIuASTH7WjGJ48SLo4LZ9LdjDj5lw37hdoPls411w9JUq/v08RMjBYg1EhRw3UysjqPjd3j
4er5mgkYSC2fGFhB0MMF+jovL+JJi5MKER+aWSz8TKqh0FSxNEns4l9xJIYmfDDsTfFkPWieonBd
JAqTC0GCjlm4NhkEifRH/HuKbJb2rgSzL09qATljq/f1VvYYCmO0T1jruc5S3tPveiyTpbj3gJJe
68baA9Qr6ARFMhaFlYNnAj9nN2kVBR9iEQMeXkoKT19XboFEid5F66xfdDLLSEMgH+r0rxNptd0b
zp5xPJSN/bJibU9CwYLN6MmIlhY7ONHDW82TqILNG+lm2ARn5PIOWlS22Uv4ExChW6fyv3cJZ+Iv
9PU6Cre8qBCUF7uQZrzXZ1owTynU+oNiarDN26/+tCzFDkrbl7ZYtICdMzcH5WzEhVPEauP3z9YT
SvOpneo8gkcLGyqehXjFXXS1+yjC9HngY8YUV0f7+K+8gmt9+fs8kxisoUYNXoawqwD7cIOrDtcP
VYUbNywCDsIH/lyWThRrCI1Tb699hjHq4IU3KViwrq+ysQ2OpdCe1+MfRDDqBgugjBO0XXk2jgVe
Xc1kwPqqXCquPOiGLAfL2mJj/FeAFk6O1vkyy914zMNsl11pN15xl42FsnRiGU8A/ed3AE9weCdN
lF8nrg3UzbhBKqBKPMHiQmSh57V2Cv/NtdILcBLobx2THcRHJY02ic9U4kX9CUhh7bbrP+DImLSi
sBWyvQh33U8ubXNFgaN6aHweR6zyvhkKY0uXkwZ2xfS8K/fcJf6r/hZtEQuV1zuifQF2ZiYi6HgO
pHS16whiubYbTUcUlBqwD5VJRTIZn1kQHPEvlBjymwWQH8QIU0Fbz/bUZsea2NLQcmtX2YiZ8jci
f5nI9Dz6s9r2OkoJoSc+CpY4mmgWqHlkNEUnRP7GxoKTCreLJ6LLU9u7RN6gR3OFEQ/7ReSyMCEp
Q8QxPFVgCpw+4imzoA5Wq638fzCGLAhrZBP4+91vowM0zviNVqA/EzNeoTVGMSwTWkccPif4G9Ql
rsHKT9S1vt+rfFSWNDYBspTu3fb1v0G3KiQcMFXZ34Zz3/IKmPGJkemRd5jNh0CusocuI/fxF3LS
LDOr4ps47FzyGNaz8TQLK8Ar0UFg5kAs0q8fKPl4xdRgH9VpaTqCscEm3XUb4uqHimh/ALMA1bFt
jyKZPK01XxdZzX3h9Uo9ebUmU9+Q2/yx+aGWiBj+joxpuALr2IZ7GNprtUkUlEpDkrDsoubis4kS
QoWcYHo1PAd9Dmb9qHPxYGU2cm5EhrckSHlaoVnLAgVeKlH2BnJhjHDcWbeLa7k5LY5YVRQYQ/0C
jMuCVm+e6nn7yJAFLGNPc/RGMQV9nNhaYCyWk5UJSgWokJFIyATAtY6Ai+P+jGNaKZS0bKuTS+8v
iFprVoL9S+mfmDfb4yX7hA+WHXhOiUWAdOgNET0omR63C65LK5C9O4Fo9psA4VLfItqw48rftpNM
mL1cL2djQ+CPGY/r+AlX82hAzM6m9T3OeP42kgQrqL7D/tV734mT3N+f74FdcenbgdG0WOVOstnq
FwZP24Lphy6Xqh/4iMm7xseJKq56sbuz5yVBk5iRuLr+E3dzvghA7P34H0mWBHnWbWq03Gv2afbP
p4zGMVfTbkQcCDZhSK5AELQj1aYJeOvhz/T+6Bt8wgQdOQvgUU83HX6XuuHbIh/2s05iFfhC1pA1
5LGbdFtOjBxOPT9rHL9JagzrW/IJ2Sd/XDmCbyBAhJjh1BGZcNOi1B7BP5Rbou3r9mlQSEFu1PLG
PGfe+YkvrlkfWxwJP2gAxX+jryzjne8eqnXNQvs7iKc4H6grzU8DUn7vJaPCcSWxOsszJq7ok0ST
q4yiKrEaDNbj265jGvyoyWKsdLNolVxKSzGTVW6ssRqkCfY04WrKZVsuIWvgqHLJC6RsoxpPSlA5
Lt86N7aMTDI5G2003zuZBtbaes+4oMTxrdMg8kiR+IgbxTCIF+oqG6hHfQ74F58KwZal9UPuqO28
Wk0n+iofIbfei15irs9yoqfbk7b1eFsc0lpa09XVZm0ks2F1Edg7iob4sM27YZNFUCZzx+CM/52x
xQdmsql0AomKMFiRxC27tk4pMVaX5WhYTRp9cD6CH29LlLu8a8cw4a0bjst9jynJP5bc51v/mP0V
Ny9xMiVRhjNawaJ1c4OxAJWrdmKQP9haXKMBW63XG+uBwlnzoK9IIf6XjAvj5nZ7ff3+8IILbyg4
Rt2R+nUmifCU5nHTuMxOUzmVPLwY90vdi5L314i3beEayNmzTUJfiqVtSQHWiHR/YKJGeI3/431s
RTfiAIJ4t7owi8o83d0P7SeD7k3vfKHGwwBfODvgge1CV2HmgAoCw6AAf/chx0QhY3k25nJv9vnj
LUlOtUNcTHWQCwsTHV9eq7w5gm35UZHH8a95rRKBYffVgxmWYYPEDZIoi+06HS6yZ9wdpCkbATcE
Wx1BIB9ko85mO01eJYAPtLPemyhF5jnMxOXGLe+KxZ6jhkCd6GOw5VYQgDGtcg5uoS8UAGQX0Hmq
CakAh7+x8mN7iUMQ9y5qdqiuwtlCo8ylrhDxJkYzrL90KLVRqO+jp+NcWyjNdBbe1+yneCHBUOk6
iN/Tf8rBYx3cVLawZNP9qZxCU3WYl45U7/cqJ2CdXGaD3X7ppW/0TgI+Vlrn3SX2Hk2hQuZMx60L
f1gGI1qiT75JvFM+6D3+TTAsoaC4Gz4av00zY0tGcB6G8QCPTs7WZUv4ZOW4/GWJe0ITTFoveuLm
5GZ3g1gsfHZZVcOMx1IR3yADVdrPRDmp1OOs5pxJM8R+PLfzCbtmaLNhyKCiYRNO711683D5SRQZ
W9Lb3Yjq+959VS30VuOWDvhZpr6kfct8TBSW2+V3H84XkDog4D8qigLKBIta9QWf3Q5+fPNB5ZZY
/Z1n2dAmi5o4g9m/6ewUUc/GxPYnjhf5YeCm5Vr8lK7NOoNRJAhqT1Fafp3Sx6MRi1NxzWqm13At
iPJ/1GQM9bp3xRuB87FULmIP5s7W7AZsca7m0WCL0LvG8Npu1SJnoXazuaa+EvyvZlTTGYm0Zog2
qOhUjUhwIcwafw1mWrmEfZoYuaZUF6+Bs1OPDow918K6D6Plqukux7GM5DWoOkP2a4nwx4OtK5TO
S6K47uOth9zD6dASwJkMJwiY29U3sCMMW9+SvcrlVf5gCrTG0QMerR0Rzfl1q6vrHo5YxMnu1p92
tqTxEUmd62mJJDS6SBnmUaHeJMwM2yKqHGyxhKh9YvM104VsRW+oZj2TRKbcihGijWSgusIe7AW6
Z9PuMXfU1O9zHmCjhwYqLyYjGU1v7VOAV5XvAZlDBeNsAR5PEaLtwneRvDetPwcpnFyugWFeAvwc
PC6SQDQQYRW0Pgt4F2C1f8BL7Uk1508y/1OmRkzsIvOnhTBbfP38YL/ue9vZ+PuqYyDAuS9pBLan
WY0zUWvGkyLUPJorxThHBJ/M2LciMXyBJ97aM030U1vPz4oItCKE63Zo6xthy3BcE+kEslOcF3cR
ZQ1sabXCzy3hfSFqYhhgmu+69FQGD0ZpTAek2tf9ZCAWm2Dwc2bCPu9jMcDPbP3Nufez1/TgpBrm
EwzllJjWrTF5ARBCNDDfiXNe82nUnISFI/CpF6tQxcWQjdl8j1nnLm68dcnIPxmTosg22SM4mVPL
DOKIV6NX7Qmf1oRfd7X1B+lOB6FmrSEYZ828im/hExh/PX4dMzLf2EaNFaQ/JLGty87tmW2w2Ix9
ZHY346oXS7LXEf9jwQaPLFui7QIg74KOvn9UCb+CLgaelr36WarDHodsQb2w0vHaynuFj0IoUlNe
mYSffz5Vfw3Kxb0Sp79+ABYgUkx885MnTN2ZLSMyR1pNQQ3x1kDnsAkJkdhD3NLijcArYkKjSjhj
bmB6X3hzTbd4qg52d264PlLfd9/4PS2G6yi1kUz1aVdzmyz5ToPgOxyTAQ08ESMLNg7sTiBa+LeZ
3XQEeXhtcKj+M5UwcHw/N+7JMPlqTO9XsK5IaYC+OG5LRyYSpHOvUgS8ttpgE4Z8w4nCgpXSWFQ8
ZwV1K2UxGD9VBOUR0sGuxHXsL/8LZWY0nWE/J/x2zfHCV5P57zzCdmoWQjp3YENGyxkweyR802Fw
iEMv+SKP4z5hQT+TBLSPv11+vqlvBo8+1sesP5bbeiJHiETnhUofdGLx7lcuSQmetx0OQSlhNlSQ
954HYyWQZf5qErNFkQ5lRN6k4BevlJYQ5fZOvhGbkEQQIAuvDSn3Kb3cjqOr4IcxmWq9bBRJ4j+0
F3YkWSOFd6QGCx06E2RO7XNECddNSsJbsHOYquQw7J8i94mufQUwkP7eEVkGOnyLZZIoEmWkPNVT
VSvE4Wr2bRg7RhGJLnjGzXXX+k27NlVXA8F24jbFC19j6+rTUUNb7VPd5bcczk9sQbTCQ7PaqZtG
hODWl5qnq7X76on4mub9azGxCSDw1kDk0kK5FNJLZxqExamni0Wlyz0xUcAahzVrvZ3korVrSX3m
W56jErFL/u7bzm4S/70iD1TTSQJti9OULFo8gX/b5NCiutxuAonMev5/9A8krJkK/MDOomF3xfhw
wgXWiDGQkVrAN4FE9fVGJi7uphnbhnmelfVHGzj5HMUWZcxgE9kfyq+zlrj4G7wTqwmVBFM6Qrnt
vYSEZdBprV3QRxg+oH1xc2rec+u9NdSuZCJoZXcY239mbqNnnegK+4DAdSFpoZoL/u3aAxGOH6Ta
uhq+w9Sjpz0NBsMOCNafl+PhqNvo6XXFFP2wOIt4/62vDPoH8xnt64INSa5QEgICAL22PgzZFbYQ
KwueNnHx3oOy/Y+GtcYe0U87SDTcVRJGEu27M8uwjBw4ipz5SGma8TJYsuWOWVmid0cHpnK6sGPU
Yaq3JaEPTwvDLY2MBqG6k5VYgbD8nIwQO/ANAsqyl4lMblEuMqEh8htb/cvEEoVyiZ77gyfzM4Ww
s1353l8bKmgVijFlfRMQ6/bpuiatGwgyNO1bUtHlvGqc519ZnV1didOvFxiKTznnMGolYe6Kh9V9
pLvMi4cf4yz/GSspt2rdqUXaZDgCfwci6Q5pYfUrbsygxS8kdrlwcAXTEU22ilohU9HteUU6IZSS
jXuLF+PqXvXmW2fvljbe1EuUlK+14l5BhM1/m87DlLdyZvQCJQ8yT0c8lSLm1uK1t0iFy9ZyXT0p
1KCJRY8uMcHtoVWWbRzFZObF/rZr3jBRptSzY9zlfX4Ux6H/bGPvqKSTeWcMeS7QwJnJZumc4DQs
L7XmVGei2K6/DhxYrHz4vRqC/Ow8C5vD352OPGCI+f1eSe/X8H3FRWEQ+dtfLw7tT7B8v1YKbuwV
MlYArNMIaed78I9PwaHXBBxrUo4dTu7DR+F30/leMAuWsDI5CM8kl9H5qKZa5NF+jJLNwopG5lI4
H4UoZSGVpU9yAGFEsIaEf//Mk+iJiCXjfzm+zrEC3hfVXPhwvONeDy7iy1vhQm+/+zkbRMqqmPKy
EPljH/LMTBtZk1THXsAKfIQw04aLYmSAS/275ybjKH89gRLNxsN5FEfTKqyWFHNIX9b5PuZP/ek4
as6keGz8pCRniGxVUOpn9l6dlf/D2W3JvENUcxEJuVTPC0dzbVvnfXk1sz3W98De0xys56QRyESY
0JaIWdDsKXxmFoNlbChFHt3jvq1J+Y7GkjIFXD/ixD6iDLPt/8KTinb5BuFppHvZP32+Z5d6XXkZ
aVaHc9XYI9KK1ujV+jx8+JIt+5UTbef0SFgspU1LEs3I90CtIKBpVbAAyroSPzz+rOP5dT1Rc1HL
m3evDW160PVSypuJytfyzsNWkANdxjqdx2jiaC+Q7+AZvNESjydTHiI9SN0EG2R0sY3qc88v9NjU
2JgSo02fJcl1Z9tn83+j5DCI5VlOW0LmMDsXQCyw9+SV4+yjZr1Zyaod5L95RwWa1QK5crJNusBe
xq6IO8TyWlH+J/y50JdljsH/fAhMCP4Mn59E/Yymdfzrhl4FV61DQDXzNyRrr+XzrdQleS4N5+mF
4BchLjtikzcYfguFXN/8gtggrosaSWdEF0nDB1yiSkiNBjPVnSMCsOXban7SAiOZk0VerlVj9gJs
O8DF1/wkIo6z1y1TkFW57BcBjVeA34+8kdBiAu7nyN9g1bGIX5hMeFbalsCnya3P5i+IvJ4iPTRK
Ic+ZnWMLRA9mdjdjaxC531KTNDxWlIzq/woexortkaGYHhLtwJ+YfIGFGRgggNQpZD5N61kAng66
cdJtTO8qdnCeIFPpLngKTtkvoXljLZYNaSBLFHNHXDQ7na0CYYF0jXGoA+xX4s5+9i3dtzFgkuxC
2FljhULWDWn2gJj+5Y/vf1u950WyhNDqUftx9Dh1zmVZ5W5YbD+OghnAJO6DRZ/N8z9ZVmJXDtcG
A1/k7yorGgQI3fiHLFwbMR6kikxY/XBuJQxDvzrrSgyxtUnc3kPKDy2Kf7dKhKYI84ewiu4Utndr
14F2L/iQ6dJpBUz82bc75ecvURGfAXVfdFUizZD0pUYY8DnuTWleTKdzexoo8Tbwn0516MQdEpr+
M1QAT/kh36Xfcz7LAF80cVtv+dJt5LSufikyKgicXRj2ZQrygvHxkG5TIcLrsEB5O+HTKivstuwE
l/6Rjhlo3N71V7DeaMBwiJl0j9SC5AN3IemPfQ7XOM+H8VUdOXfEMMqsxgNo+aVgZlE6amPiSc4B
U/0ZWFAK649G3ARRIjBvCdETFdsYXY7KrHwc8gUsXsQAcyX6ZgnBQJnMCg3iRpkCwgbABURI6S7W
JRNIjLVb1g9pern78szn024Hi+J5RuSslFZdM5cC0qX8CIk9LOYHh/MLSWISP0P7TI3z0/TEh0BO
iDHtN3uigkWWWVEnctSRXr1RYbdvtN60LMtYIrhygN99rr40BN/MKeZHx1LNDjWdT1wzkhfBob8K
cjf+eDZqhQqTVOm2Bn0ngQ3ijFdszl9meLC/Y5385QRujTd++hZIsErLfgA3G7VI5IaQyb79BxT1
o9h2hJoi5WXMYi0Q/BL2BjA2+VSPhpv4stttmrv3OMZ1+wdWy7pH/TH1l/wqE3fa+ncKjBYenUPU
/BbfZ2fmWIW2gNbfh3YUB9wcuECx7Eq/PqWI+34evZM9+yVl11TKcaIYB/kOY/r0GsEwPcQVd8+8
23QfxWLYF45UkLwY/p6CVqK2HoOlu6rQgsSmSSHMqzpNwKaO6g2GlBZU3EnGPoCKMHD40fTUcY9+
iv8uSw+4aPDUYQnLpIZWVF3DDGJjfHumzPPga2CXaXsEbxBW2k6xOuxgnPLd1XeT4sl6tkES28lW
mnSMzbVBtT9HagTdyWq9EI+L8fdtCfzYGQUgz9grsM/d9qAj0p54gbALfG5k7y7DWOkwfk4bq9NB
03OIPzgzsWI/dwrCqi6kRu3LgKK75usW56v748uWKfy80THRJ/RlAJMA8tyUSb3e3khZM80e+kG9
F87gobzcZkKsFPbYzZDhZ2Eiz/UFDAijXvg3AhbS/+kIG6IhpbhxTsGb+eLVg8zfnGuoQcsQwoEF
cGH9Mcvji8FXx3lJF9aDYbTOk8wvDPkyndMRjWLUXg4gOypwcMt/oaG3mg28WiKjVX6HI4XIHD3x
spG+Kqgn8bu/g1eU3ATQdlr3hHdZWk7ijYkeSgAzm7PVvlVSAhaR8vcEqc7BZtAvx5AbauvCCWbm
QcPKKfAqHWU+AukjySRaVyU3kXN3fKIvkfJ1zf53y0cQfQvuslT/V6HgX+y8O487RHbrIrftCUaM
hvnEeiLseBhbjxuphoXlaOYhYaGqXDnCfhxudDO1gJ6utZCD33iJqF+Y1NDdHClQM5WUKmOAOVNA
2y71BP7TQU9dhEjn5mz+qI5JUdazS9KAcb16aLVszQfYm0/PNA3HLiR5lai/V8x0qwoOvYGj2mbc
BeW1ZoFEXOnT9PEeniDYALxC0BkBtnB32VcPjAlKJvKfP1Y66LYpy+HrPArejXdVCa6kgoaU/Xnh
NffOaZxqy5hwidLJEZDoFzhLlcXR2pUWcR7Zca9X0eGCDntcH5LGaQTWT6P6oOv9JqbYL/Z9cav8
qOekJp4Af1/nLyPQmPhBlbbVR9ITKBwFWMzHz/ydmv99DPF5tghyCeG/X+1kpV14vdbUWVOurc9t
N1FuQh/o1aM7LaMVpxLOhFhlnF5tQqRvs8upeRFrP23/PvF93Lr+YUwjgGCpoRWlVGghuw0zTl30
3ufbJVZJoSyk2tYTfTqCHB3BLCV3MmW6cRpctGgZmJ0LfFpjrRNASL8cuKM5mk+q6NFAi2eMogv8
LDmJ1gnaCCa8oANzljjNAwHOF99sNRKC/9CVxurWRKonUn0ocYLCMdUSOfBzj8EEiDknhsKMbq3X
CSQfbBoBYcYatOzpjtWz4K9KDj4Su00VSLq6xBMbkzK4tZ4OpzqKq27woHXAhgiJEvibfHBIDUS/
/m7PidXD6he987Vd/KPF4B0DkmzvMOGZewt83a1tR0nULoSsD9FLb8WUH6K2ZWlXRE1P5eK2fZNo
2RbZZLx5jZ5cYSBuDCgP2SIiEVsqxfa6Ri+3YLZEHVRSS7PRgLreoNHO42L8l6zEJhq/bwwahNTi
d+VzX9BTwT3lLcKer/wxK2iUWxiLLGzxS763dA3V4kAQcXNMiwp0BbCuhsCN6QjnzvplqRHk6q2a
EX5v9gRYUSp87lnyZyqQ8jBF5pUk6moKoGs7RsO1Kqegdzz5jfFDr89SpRcAOtd2yWVBJfBwhGvZ
GCin23OBsH8X+/1CQb90O/1dKP39w5HPNZu81HGBkKLirkDxFoJesnV1FXLOzZp2HvAWZMcu+d6g
5OTp3ixNUOc5wj95tu+1lsHyL598l1ux8dm1pc7Ndb42+wl1pX5oaW/UFttJ77Syq6pKWFIe0X5t
iZtRDN6EcwOLI8JYDKvB0YFQVuPzbuDigi+11dLepZwPDgZEnGqYr5Uij2QuQ/YEn0+G3P2UUwtm
MU9D+m+DVSHJhqKUWOnCY4IRoYGHiTfKLShIPT5JC0csYuFOPxllQsaBSGR0nuvkePNB1/6ukyQy
yEyhZl7hrht8m5Trtion9n//9Aad9Vk3c+XvxA8edPMJAyL5I5tYEiXwHkmO+6WouDkpflcsrmCT
rhIu+fKPKVReTyCi0tV2jsiW+OmizypaFGEZaCW322EoAVBznp84VW2vqHKmYHVfhrB16uINXIC5
8wy/0d/NwDE0aHEiMXhXX2G0s4f9yLti8+GAS/YpEICkfZ5y8rCDhq8BmtVndVmPuK9f66+v4tbl
yYlJj7eR0/srKpBNWSQzC/qPu1aq7UgqhzqFnn+NphVIhcEdTJh9Y6OQvJSQyR7jnPEpbs3OWrA5
MDA6nTivC8sxCfbbeBUQzQ+IwAkmUZpfOwGN5bzNFGmPaVAjuDs4Px11BEc74GMuBdblpOmRK/e+
ixcx/TI+gpQNuFK7uxeFJfJgJUsUvO4gXFJQ1Sc3vbS5GRK3TNUenDGS8EwHB2sBAkPH4fRQDDob
KpvqEX/SrPocGFt5ZKRm0qvxZ7PB3Q56XG5t1Bsl4+Prrz/FJideztEiAUOe9+TI8I5n2JBX1BU/
467fJxxVt5LBgetQe5ySREmih5I+eHAnNNG2HPWSfBIIPmpHizZPqkXJvII/Y+HkAfBBbt4VApvE
rWOs4wycwgE8k5g8yTwWuB/CRhHEy2gJ9zZqrNYg/oSRcsuWY7JMt6GjtepKEEibR239IF8IxPm5
mEVZBKRiyVeZB/TGr+oYwWV951RUacwyF9ApbfDRQBIlVrJIry34u8cCgTmyNlorAicmvaB/wV1m
mP3q4pfOF2NcIZc5nxXH+AGKKThSxLMxdFkFKsCqjJc+xpO2uYrCiKXtUaWCd19SzbBOk7DZRc5W
qQkmIS3KsokLBwtCSnj4o2GctEe63V+jQWOpGZkk9R9M342tRwbYWWTStYXRNlyE6JhSVFuTlj02
PATg58Ldc5pzi3o43gROjsW43YNX2+r7GKr4G0cFZyILEnpNLstkZ9fJeASHd5iueLwwvvlBizv5
g6K3LEdgn/10rp3qVSfY8KK7TSsAKpcgXFI2tOrj7C/7dykGX5x4x94tJ//+DbVp1LiLpzi+E9RB
YpOslQDa569U+o9X3d6oTrV6vcPp8V4tDtUjeSBgvI8RpVZcZwDPA3KJvhpgwbOBn7+h042uHA94
OdC7kJOPKs2Nf3yzrUFvIMTkv+wxI2F08xmvwx8Yar2lSU6zxPG1777d8cugP56gBIlgwB+JjWs6
MFOkzuAwM090Mt/oE00JcU4qkj3+3NCgDkTbdphekdsKtBbMaklJwaByp2auJ2GE/RGZamG3kYgq
hwOVhzf/ATYEvHL96wT+YX0vb2KIDE0D+eQtbrPKW1FdfzEPcGtI9kCRT9IVIEW4bCwbXyClknzO
iiNnag/5LT7v1ZNf0Ob6NwPIzl0Z+6iGwWL+YbLI5tHw/09adPOoV1wNY9DjBwZy6amJHfl59PjD
ssKsAzthuXhWdpQD9F4eDcPGpJIDJvp8EbO8Eyd+oQIO+ZPjSjtm0MWB6vDqOjrzOGtuiwE0cstS
gZgSJ1GRvvKni11beaww2/8HQMg01dnkV/1cMR97Z4r6q4vgGRBf7spF89HY9wcB/68nkTHmdoib
uzKQmJmLjxW5M3c3FvS/GfvU4Q6ea/f47Y+R4ZWI65Fq38PRl2W7ys1WsXgFY2cALQa8YKRpUkqY
7z7XQzZZEAwOqKoWRs2WiXKrPuMbnSVDdEbBc9kqTKCDs1z90haPe74XJXG1hLzeEVToXF2yIxYW
jV8oACtWbn05OJbj5I1wM8lATwedBMQ55O2cqrIXtnNefwLahNOishAveaOi6ruwgmAfZ+2LjaNS
MXwW4MGFxZq3VTyd8fpfO3Ma8lHJR8fP6jpvs52bslMqK/V70ukfz3sYUnWDomztBztNk37xfL6+
GhYJejB6hIZyCZKvJK1GtpZRW4mes/5ZYCGAwuOIY9sLPVyGdGAhFY5TZf5xd1oQLrx1VAwAG7v4
Osjbfdh6IgEnyMhwwrMzzS9ZqTrJvNnxSk7LdQ2ayLKdpjNJaPSWianYmCD9d5R+6BRUqbr9Lo1x
eZ92kniOfDBWGqPwn4YvI4K1RYZ+sddBEVlLBxN6AKnYlxzifSROMwwrC0IU9aH/GbUlpCxwMukI
UB7ktpJX4EPEr5gJO7AMzaAii7236rId9b48ShEz1KY7K0qDDb01bcmeF3QLDM68fe7yzPqcP3ul
zjgJKJJLCiuzVsXQ+33WCcr/BE4kmuQGafmQ1WS6pmtIngkhbtGXYniQQX0DGQgygorIwNBL27KZ
9pe9fGqQg2Z0y/bdQ3LSgehdETWOWN6xRfn66DCAc/RvQPizYUi2RymyyVftx/QaQmqy5lvBnVZn
FD3mNpirNCvTN8oEUw8n9Zqwew8CpWNf6km18xgBjIqYk0c+w1CB5LdaxrP6UYdZj1V+qtkQmcNO
0Mo2h1eWB4xysAMZ7jdk6APl+BNyVZrI8m5KyN4UatUVbCG6zS7T8aZy3aoyfoI9ZwAIIUFFoHJQ
WySZOwhr1AiQJBWelxB3MhVIYz/0+KrHJ665d2jobvhkVM0O/gPHKuHVJkcdDtCTtjIj6XFoyUzB
dAtYyt+uRvCeaZs21bqDIWnjy+ZsaSjAHlq8oCV5w9nMdgwG8gxXnJWLmUTGhiHHnspTZlg+/ECo
TWLACTbTO0+XZVLA/gaKudJy66baiM4wvbpUE1UibR4wF8OR6fnD7sLAaZqNYxwL2vnaNyCWwYKK
hv96l/BWATP/RX2oLBe7YMwDtdW9r0C70D6IfDoDqHlBCIp+MEmbMaUsI/S49AJdDjrQFDi8OnnY
xHK+dYvmnTaAOdqkxOK4EFq10ucwN0DE5Ki4k+KV+GayomCjCRknB9Rg2zRulzhAILUMFsd2OSbt
DixEaGm8Kc/sB+lxyjaZ9Yj2EKvbA94iiCIcCMZ1TvzuJguRJhgz4wXOirafyAx1mbnS1XicySdQ
zjtix2d8xrPji3JEUopuFYXVYonoytKDg/D6nU/JgktjcV+M9yDko7kNIuBD5xIVZxgtkv2dsblS
DTWKv+zYCuoaDV8nt8FoabRp6KYw+qQUTEN7vpTHE9MH7nHm3h95NS5ZCi9KMUK9sv+hxfhceyMy
03zZG1TSdK5wLyjOezSMjlaqSFqd2NQTf+hafhNUXnbENkR5vjUuKE36OkPE4/ssy/c01tpBq1lG
ka3MnKrQVFxA+xCN4H/lKPMS2wqS+vPg30bTFt1pwqLwPdZsmOX3MDU6sYwX5QcFasl1939/qEUs
+N7IHo3F1Yx+e58oyXKg8Jrs8Lre/hcbdeX36GBX+VB2BCqWRGZgUG1w1k33m/bgt4Zjk0LtEK0j
PWQ1ALTzwnn4K2FCsuedy941svpDjvZIG2r1w3kFX+1rMo6ZlBWNihFrh8RJu4JRFh7oMUHwLCmT
E0Wt0EKGTQt+tlFKqjF8Sxxu1STdO5L/w/TaDazyW30iN9bGAIS1gchhcZAuSpzwHxtOZ6jKHJ7I
p0uC0nKo3OCitOGPfDDqyVNWNGq0g9F9B/hiYLSLvMu4DGBHrh0k97bQ72Dx+R5xYRtOf4/r6nXh
eVtAAxh6pYDMxxQHNHdFbuzjBuKevckigEesU60yk5X/UzdzrqOfflBFkHTe5xNcz+RHN+o+Un1N
8tkiu7GgJnfUmbPsXzS9NaLqFCQ5w0c2WIu3wI1EXhyAC4ejVac3MmzrvTPTCWkHZmTdpHae9FmZ
M6ebcCVob8Vhfp81jWo235MS80AuFuLVFIhHWaoLfoPUc1s7qU7hopyd5VBVOmFlm2wwDKxhgUKz
m0e7vzegrPk7R9jKbJkWQyQRIA7a3PpE8MpWFlSqKoku1/KZbvg0khDJSCgtkjaW9H2pzUY1Ue3Y
SEa+kr3GCjo559l/7lRw1DX7ZZ72fgh8l/B6oJL0LouMDP2TULICbLC/w6h9BkjJKKETwroYAQgg
nKo3BXwWDgP56m/RdHHCYg6ZpoCfEGLdvQFVPmTTf3DqgMsO3AhR5qiimR64TNSo5mddaEVgMqLi
3/iVUPsJxZLWijdygq5UdRJh7eKkmMdbsAi9pTA126oer4TWExkcvQcWr6theUrRWBZWSHfEDm6W
S/U5lZJu1t9oyJDAUinnaLNl/s39k0mbA8x+3aIwNXXM7JAYHXQ28BCPr7o19aUwwe4hIK+LomPK
r3n2sHAkbamwYM7WjqJvh9NPHC7FkCrCjnSF4iuUrLLFqJL0xcey+L/HcJq9R/fjCQt1J3d0yGUm
zRzpY6v4irHw6LOjD3NyFevnrqq1okdrqovU1X42qHYs7NIcNk7S5SNyD26nE9fT6VLS4SWEXluO
xYyNsB+OT18TmAlFmPjqO5gejfnD3InJK78qrIwWlFs8h0kwN55CVeGHZCh8KzuKmzAOEJ7Udjn8
SK3w5JhmM7dL2WG4gt+J113KK+Wr9GCwLzKckqWFKxlvCNMjaE/G3vAKPkqqGf3AkC+FxzUEOqRe
s9nLdD+7YtZaZukR+08LK0VO2Y5d1DOyuPi3pjiLbipHzXgI2YiMLRKzQzIIdNasWhxt9ygVPWI4
6IDbBIfQpkmsmPnO4kN8LV1f49FXN1M3zZ4q8k+EdtumyZm2r8VWmG7eEmKJ+6EdH6oJufw04tm2
8SFY4gXcq6zmVL1P+dwuvtaOA6Yxdk550g+RshBPPW7EhS5b2+iUGtlw2uKGVXjYh78z3FR9If2Q
rPeuYmp23s2SkAL5H3oEnLycdGWY0G1QGSTMfYD1vflc2C87RJvN3G1wDvzOG1njhrm9TWT+x/ZW
2ek3bJ/WWo0zA/24nIcsbZa7YXqIZ7VPMKnlFVoH9JKaJguPN4LzYikcQERc/AXsn7sfYOftNPbJ
kTnoQts/MfTYTkv+GrL3qLtLwxMiitFn5ABxkXVS6L37X/IG6YG7OKkWCDmLt+KTSQVVCWU4UVqI
1Lga+020gfpokMjSNBm8afxXj7n6IxNuKDT0LuQBrTxMB+AwtnDvRABJvTDStZGEa3uUuJOh1/sk
PPpzwOfDHQTYl+iQjOEm+TD1+R25/FCTuS6AcZLDUW7k7ETRzYgjgLz6Kxzo7QtQMEhkVMZbkHh3
/ttaLkZ5mCdXf65sowIyO8TSHppF8tAPpnolW8rPQg21AMu1DghTgNlCV/DeVQJk+NUoORLb1Iwy
nbx/6qUCymwKHZlU/QTsW2aFJuoW7Bx6gxpvG90QDUEs4P9G80QLrKv3P6Ndk+yMi/yw0Oc0HbxZ
/eunahlh+UHWzJR5DlVhOaoVzkAyVXqLjIXRFARgMIAe3JHv2aotfRQnSos3WuI98KJMzdGe89mN
k7sRiY6F+dmbOlx/FfWdkp7Ve3QRaNTtanYTzRlWwdOyCMSHZc5oPQlhsDko8zgBRqXKK5gTvTyK
9t8P4bL9YC5idJMvzo6e2vwtEftDbSAcmEkCdHlgNDT6sv6pNwBMrNjAD0slntLxslBqCrRAa4m5
d+NhFEBWp9QcDzv0Cj3/kBVMatLpKzR7U59AfVaR3swYuH4UWH293uDlcsD4YUtdTNoQXM2SAktd
9sm9cU+O4zxC+m9mX5mtc3fn7wnQVYskUT2/1AGMWULjJ/8PAw5X66DBaybLsMNEJKE8hCBA+hKz
1SEp/hoQQeUS60FlPhYpbo3aCXqUYbjx5ys4UJcxNLmxojDCYY8jbFO7jOFuW1HrZigUbprIulxR
FcW2mTXm3ZzqTtPe3R+AF7wRmsLdpdbfs4gOreAQ12MBgqaOUkR0bbfqkFW3X/NiKL1kw1rJrjRF
3aoVVj40G+7i8ubUMY+n4Eh5vnF1tvYuYX4BDRbQWvICh2UVfP/IaDUTJ+wlNbBYgSYGQlkQGuAO
AOd4gZJKgP3UqLoDtNlVaIrRNj6AR3dJqzOAxFrLAdLYzmZzjhDqMZGO8kG2mwYWtsQiQwANQ7M7
mz3lFEVEWbeCL+VIfmXeFLkIJj8mOeEjy4FOHplYv8vWrNwMHjFMUMxuCibKhOw2n42EZrKWK4Ub
EmeyLM3xNXKMDtjhBzEDAJj8UYnyrOyvmEu+e/ST4oHQhmRaKguQLjn5ERFcsEciJo3CTuSZZL4O
8xR9D+QFxPjxFVO2fajmOYsTGttf+GCvJTmEApJXTqSsCMkSBtpk9yVQFU96ttzWlwSk3/G3hb0A
S8dUwH+EM6RF34kCvZElkk4wMvfC4apGr7Ot6ok25z3yV6gACCjk5qRnN6ALCk/Wcb8174hfcXsp
MIqPKgYzincrRklGF7pk8BeUaP3aXSNID1eIl7C7mDBX9IE14jJdtGJA3MmFScNzd5b3fu9Y+nVM
GEDfKtVZS5mzv66h96YeQ5AuyGX4zXSCvHdj4YoNJLBnctoO3p8cflyhtVnf0rFOqSpVmoaFn+ND
m+QhxymaGxZBae2b1DpWEveB2bE63C2U7w3n4TJurVnQayubetV4YQ+9Bh2ZwRdkB/bFZfUsT4/Y
muK22TliQV8A12cVEG/zCzZ5hijh2zHZzxgLqhah5cPMNqAXAF69ENAFR1ic1HYq7iT0/O1ukIua
wkwG4kRy8pkMB/sNDgchQywtN5ifCLb2IwiqkjcA+6WaydvcDpkbUoW0WM+Vcg/zWeFZlmu6MWJc
5HZ2M5H+eH0St4P4cIgo6ZAm54llm/+xbqky5s+EVbca65talVjtYpfK6KkCkstwq5OJE/k1u2ny
r5H1C1c5rY9f6cxn42yUq7XRcuXhYwfWy7D6FhoRKI+7k64hGlhxxIF7x4CWCwicqXUlZI4Irg0j
TuB//vNqINKUIudDSsAb3uP1gezvLhgvb3MgyIXdCkhawVsbVpaqU9tnQKlK/aT69DZ+Htt6d3M2
iAowdN6HAdRY51ffluE4v7QvfOyiBtsKvPU38+eMjQA5EguCJyREBRC7pdoLJAAeGNY6ZClV+WpP
MTrPs/ibgFi3EQ+gLvk8UXh4r58QTSwbw201IvGhvz+tVSxjhA21m9ZNkRuXX1UAGk9GgxlldOG+
WbZrIuzhrBASLpg5iSlIcj/3NASVt8aYD4OLlp0eEhABPSoNMJ4vwRRkBGAaj6tlw+fjLH5wsIsZ
rfCSKMKhY6NhG4Z5Uq8qvMEgrYfU+QNUfLn2MSKkxaJN+zU9qqray3Tn2BCtL2+jijhzsFXK3gF4
Tp/WZwqkFFJM8aNjQSF4+aNLRAk+Nq765GgNkpJx74N+GUr6oOGPur0lrvKiNaqHNgDYSuqvSuRx
PaX7MUtoSRPIUsWiBTQCVdGXTy7Lo75HiH9BVwqFSKV4kFA8lZIlL32fr2JYi1FeBp4k2gGn6+rG
7g5UCMaVxO3XFm0k2EuOSwCIwi+tP+P5z2oO+61qrwqNPsIHRiPFim4sX6+VsJJhyLmA0MWe3gE5
107/VTrNK6aLdxPFaK4qtRUtj6tzY7EF0hxrailsp4l+qoFinDmuAZc5pf7ulUogky/bhAV3okan
2szbQg3gRDb4UFh4hAezVMB7odUW1A7hr//6EJK/F7HoEItoQKjoqqAlP1Wm6jxLIhDuUlTOw8oP
cTtmNCFJzsMOjso7d5Kc+bUGDI1us0UY1Rj5l0kzGk2iVFJrvVBsQAEdCo6KVJymnnZTfbMZwp45
63YN1IWA12IeN7QaTkb5MvAOsqcXeRqUWW6GSqVVdhg0PyMU04+srbmvfMAT9xlrSPK0njOLAZmF
5RxQdYgeIHRs2F3vdk4EV8Ln7WAvntKJEh0AGXJgf1JwgA1xMDWq3hU9qhQTx2GMICz12Z2215Zq
OZZns0UZCn6ZaUyT3KfrqkWzQo0USDGM9sjN5vUNJuQKY0UmEUkd6xdHb3EYIJeisSvqMbT+9ONt
Up6ASwH07kKxwZ6txqGCeSIdfeMetO3JfT/PFQxHM+sIiBZaQ9AORexgY0zOxUuv9L9v06quIYC4
dBM9I8A9uoOZh+9lWGNxHE2S35C/WK7EtPm3k0v2QZviE6oXxYJshDl9RfgQbXzgQkbuVjkO3aIY
/nRMStiv0fnwgTnssvzEqaIfFulXhxlnwZZ3RyoUh8etEC/eYGmi/iGBQI9t84W+2aq/3WQhMnyU
Q/retg5oxo+Dw9XM85fAKX8zqte1/7aY929kddj7SCMOJ2+TEvIVs2xLkHcB6PO1dYfvdQbawLYJ
FHfYO9bn5DuF7R3+tG2hrlllVanYw3kq0qJj2h/WuH265mDtP9Dwf4QRLB2NsbRln9BIkdvrBOAX
wUPRidlUsibtOZOEiguDzVMep1SEQkfv49/SZXBybtQmgyPweZcw95M8OyrhYTu5LdWAP6ywLLRR
R+aUr34ooTK+RFXSOjN3J+XH5zizsNtRSOc3AZ02HY29Rp9va7QrFpVAY+ZdMtS5iJn2K7U077mq
+3c/poIBtwBJO8UiBHKvfoN3hIM+LZp2EmcfegBfbahv98vuMd1x8eurxfnhJ2C26PfKpvaZ+52a
lRYN/yajuZEXqysyuIduVDVbc8IwexrlbNyLImp74NkE2WxAfHN8A2M+18lEV0WDKlKBGMqeUthy
oRmJKJgJ8ZCwFEAhPkHpyJB8rPASWe6do3maoVqS4fFUzQDZg90IgY/imEgxYkGrn7yQUNLyS34n
hBNMkFQezh31oYBxso+gK+deHJ4sBAzNSPM+9aCYxgbotOTu2Ge3evqzE1gUYltUkhoTI4hoe8qC
VNnw4tbM4fJjTF4U5UxuHyW+n4aL/Uihv834mWb/BnQIExvvJbobVg45aw5vzSE/5DgGeBtRYM4H
CxXlH2qP5ddY6l98dc3yz6itSNnB0jK4NxCjGjtH4CPzFnqpZG1sYwigc+4bZXbGryTN954f95z2
OGxoVPdPkiRyU03VRBRyQzjfuZ1AAfbZIPjySq8lgEzk6r2JbeXDUJtLbz+2F5ptjXYvaeMGocnv
8NNQF3Zp14s6d4ZBIiBG0j5ufuzw5R20jTZlvG9aWF8Jap/tEfTcL3Z3J+BGbeTr16cVvg4uCeDB
AOM8O2xFPa6y1qNblM4lx151CiY0sTOP7XLpZH6iwBtj/hLehI9gJ+W7mpe1Lc2OyW8qvSAedv+b
vSW3LzsEUYZiY7SOHGGf+2D0W3WYdLzug+d0L2Gw6abTOIao9Q9jijGD0HZcDMtZrSqXFMivug2q
JWZ1v3oVKXK0JNKhNMuJIsj89SrQXb1azLOkeVSggODhSm6AOS25C+WGlt+rSsYWqrX/+V6Q+BFg
xsqlZ7T1pJjMODfPyDvVzntKh5Z1uzMVndJU3rX2fghTUSZgFvzEdnY1+WLSqec/pjzlWO2cgstW
DTYa33NEfk5Y8ca2+zixw/L8OGb5iQFeUe52ONdqQpwpY5e66SMIJNP9HkzpE8uBQ+/+5JMN0adD
BqYwNdtz5ujLJqeRd7aaB0Ceh4Q4TGJNP/rRJG28Qw0jqP3gb4gkpVe0oieMMZJIlsmZtrIM5cQf
K9/Ne2f5ec76nvJsSWd1CqaRspHnpNdoVw7W77vSV3LAxK3muzXUKAjzitlZ/wB6L//xKuE8EUrp
Wnq6Q4McPxxSdu/8jTdrptqH+Uxp4XlTUYF7FKQfS73Bh2/wlHoSjTWl2Hn/Xz/D364iF8jmh3gy
L0ZXbM/Xip2v2P2UckviMdaQN+4RHAFImyNx1+VgjNSbdgNePixuJ4bhPpwd56Aogy3Ud20tYYWh
s/8Z75IcxDPJKHtKKBR3x9Xa8MSAkq3bqTBRx4ImA+FkzoPtfsVHLRfOmu7UIN6e4RIUgT0niHRL
ZjF2QUSnrJf0XowKlPbBJkcvJy0nNvYLLzTODAyUAYNLtNFhGQF6Wf+F345nGWe9aPtW7uF9mSqn
7vF6WhMwMwpGZ+NdTZGWhUNsr1OzcHr0gY9I5LtBgSuZWgi9YBLd0kN2qPH/L7M8UZjrnkUs64Rv
lM9C+qHJ4XrqBPLg+QP7cdpYdvN/4ltGR+MNdzOqtSBA1P2AUuAUTOoQ2cAEMMBWk0P6Xgs6JVSJ
D2EJZp7m39IjhA3YeWjHJMnUlVFxPsW7UUIo5LBNGmMB9oCMmvZXK8fJSHQVClVp27AIghCKcyy1
k+CH7GcgFsyuNMvaHoSfad546r1kPJcNW6MVV+pPUQ9L3Ap857dORpHLl1bIA2HWjgJvbal5KoYB
8wnJ1xDmq9Xy8nTCRU+rnDuTpPgfEhu4tfUG3q1AD7YVF3VUFQ84rT0DnjM40vP13dnHnpOLGT6U
kColgnlBesB8M69RVTRejzTOonOyWhI+7aPBcT8YuoJlVata19GYlzaxSo0FW3H9gusSl+CYKydC
J7LoZmVa1oZX3o3LmYNIaj5StRBQrers32uK2sOC92cfEUKIkMsVY7vQ/BldoxUHa7wgYy0gjxEF
GfPZ70IOE/0EnXH17gp3z1NXI/JS57jkkq/OoV1VqRAPBc6oUQtpiQT0TDxte1kb5j1uTOhRITDN
u+WlLZZpQvfd6fWIPhHpLgLAMgv4O3LNeMZaI1l5QM2jnwnA6lWtHLBPc4TVmGbD6L8IT2DEaSGi
Kdr264iVYPDY76hjhSPzzlnW487BQrTOfuBy7wUoYc+5n2sUl7ZZI3MjghELJy3ceG0DyTBjPvVQ
2gnl/fCSk+wKKEgSxQUo6zJqlF2S3GjHlKVp13eqzG1lxGvkyOVjGrhDnI60mNgPUZL2Ic9yvfEA
abCQg/2Ynvy7sKUyRdOLZ6v614Y//NzVzhQZFD5FfPhTkJ9y7/ugtw4uGQqStxskOIj0DxFPYdCK
EyZ4Adx1NlENHXTv2cbo9jZinZi5DtQkcdQR6RvqCRZIV2TaUjDf/b9d6GC0btf0euFU8il4JBup
2zpfvhsumqknW9jGDX6n2RYzSWimV8pbj23PAqnH34HdLVRLDpRf4xC4IMZjFT7AmI8TkiwOVbsX
z7fhQBDFQp7prC05K5wIdLrqhNN4kvfmgpJtl514mCzMkIf8gUMD9x7j2f4CzJareWx24gTBXuS8
FRu0kiQO6nbjwF0vgc0kw+aftYPy9xr5V9VR4MUUHHYgtkF7l6tKNoRT68vb3vTnyDzUZsZ7l2dt
spqf7qRTHRrESi6BAe7d1fT2t+0EWp5ZXElacfJF+3ooutU6iE9/w6abw0j/G9a6/Ec7WkhLwGQ0
IU3fMkikA6WKKEw1EF+agPeejsaMbKbW8EvZxpe3M4P05+k9ujH5orOKIupAo2jG4b/fCGqCUriB
w1Z1OA7dqVGFW1gwob4qvkGHwbOBxL+q6jt/sC/PUHW+jvzbxAMGBjDhYm6UUK1n3GHa6aWCepKe
hNYFyJCH+0f6G9F6g49RzGNjxsxuf2S0l6GyhuPoeEA84zbqmsbv4tBdnWqw3IlbM5FOD76Ho3qo
mMpHNf4BFnJ1Sdsz1CIVIsdmcv8+REVhheU+YwStzlH9qwsYW1VlHMFhdq0BbNLtA2xUDEORStGK
i3ba6D+fRMnDkO7k8n17RvoZXN5+H20a+CCtzr84wIz6lZRucnAiG2qWYZ6EhDdp0Bbgc3Jg10h6
lV4fJcGLQt8twJ+Epd7JmbNqJZAxCuYHR+ITX9J0hAetmJM9xekpojEuvdkVckAHCWHSHNSZu056
vWqt7kAJ0dsJ+1AuxoEC+2UAXz3WexI+hg+tFZ/vHH/9SkO6JOzUT4d69a+eBCjGeQGjunb2M3hR
QJPiup4JGYmr/1qcKpfOoR+PON+4+lEBYi/FPeF23m9fpDr2fLZUof5HzlKIif9g19syBvhhV0Rz
5sHEAMB519daynZ8KWvoM/Fe402QWPZDUjCA0ccuxjoRRRLG6iml2xPj0idZS6k/jKQfyX6Z7+bn
yVEE/XpoOGwuZuBKlpIzEYQu4FDwYwEn0KZaY3+QfVRPy1sWDNsKR4lfs4JY6pBSZbP1LK9ASNw1
CK8c9NUei9/VoKBQSDTA0mYip0MXY0dhDuxOY4+OFDXClO1u8Jb83qFFATU79B4jZPo8FGBq/E8R
pzGH+yCSiGRNypLFwH96k+lZjh73waPcjO5eeIvnCMWSs5po4SP0BZonO7tVmpusQkJJm5d1tGyQ
18RDb8UDTLbrGln+5XCQjhffm1bt2qZjAaSkRDiq8mY8CCIkl+QPUGuRWRm/hOmafcVc09hBblC6
bXYgqM+ox0QUBDUbR/jpP+VromLKAyzhgBPd7vPbSBuIpX/gFQzdReunDWsEx4SqgBTgAgW2jMA5
onbtTTyXxBssLdzPyYrgPlMZ/Phb0apXdm8SvsH2l5N8GdGC1nMaGMnaKozs+UOsCg9sz6iu8fS1
koBEKdW5DwvSx1cKJ5ol7hf4qk1DF/9lR4QprnboFTXt9lYifbswOL7sPlmVHwwIxbbdVVGyOQ3n
/hh10PJcX8Qwp/eCVlrHXcEJNa4VIP37GGKiryPm7KpcxUd2K0N9V/117oSeEj/Evic5OybL6qxL
VxYNmhh3RqQHB8+eWAQEK0qi8E9szNGWpwO2bNf3WluI6C9FAcHfIzUrasmoLanQK8DivehL1jUq
aLNVAz/zHm5Sye+2dbaCBz3TIf88xMpJPhAnSybBcQQ7lnrvylk6iPJAIL1TkcAuM7kYnUHr7gs3
6xzzmtdU7skRY3BkKd7fVrBmFo6BhrWk0f9z5a/l30PRo9ZD4rROeM3xLw9CkW/vH0zFmGTgvwRk
5NB030ev39qDKg+lFsjDx48Az5Bz8wxuHHe+ffMBbrEcwLqAIiKrB03gvRv7ozDbffbzmJ5dk3lm
5ZQTdiZWANmX2I6WMROscVm41hWv1LtbCir1pLYVFXxC24e0tDFNMerC9Zo4FCrficFgPsM9EfiW
BrZY2tnYWL7AV7RG3AS33f5OlKauajFm2U+tF53Vwokq0OaqUI9XHmT/NiT3pwnDJRDrA4ToHT+P
/Xvs8jL7E/zuYpHspoLD6HJr0TcoqdWyGcN4IEPc4TbMKAvp+8iMa4S4Budw8GNQ4DwpFa+exjTk
wXhoKv99PtOGZZ8HqHcXbaZULjzbWBS5rNhlvl/pnVC768GoNBji8i/DihH4Ihwy6t0rtXxv9QHi
fmKwEEllZr1OGn1/klgl26LZxWsQj92ryksq4j9roIpfy7dxHjLAvTSG02l2Tki4ESyU8GS7BJdQ
gOsL3UDMqkBon0FRi4LoFkw0HfFFJmtHHV1zeg0Lx3D4Ak6b619KZV0V/CAIkNzNb5SjJpEielSl
PjhLzVnbFQ0EMlAaeQJURSG2Z0yTd8GN3KX2htw+N9Z1q8kxXCES2V8zWAhUkLJ4CX6fVXzMulfT
fBfSY9LWB6zwJTtZOkiquQIHpxxk1o96TunbMC55cm9WeQRJZP4R3rAl6rNAOpPbHYiYuKkF7rD+
UBPAC9PUTtWDsWBvtCk67oHZw7Svcx4agsOOx0fFe7atwrzJLKp2QWsxIDjSyTtzMsxEz/8veud5
QWQ8RO1XEZKKG3rPGTtDgWJHZXBDGc2hjLpXtaFG9H3GtS1L2pNC8ZR3mYC946BXug5hsewz6XC3
JPYCJv2WfVbAb6KtC5NVpudzfVnVyadRFuQsIMH2GxlllQB3ybnNffKEwIteNKgKIPW0jst9iKt2
qd2Tc6cwvjEOFw6MgWnXeopdE1ZyMBCdf5kcksQc8RFz03m8o75TMl9nOGamLuCpf/ozfyXsQN17
z0Z7YteOj5/1VqOWRc1C6N0JCgV7kUEWJm9EGKz2bQHdgC4Z3zl99z9tk7UZZyrVneQvuURyrkZ0
56jOgXEmTebjCvmXRTxYe3AQHTIfo8i7QdwkEzICa80ddoQ4q6eCJB05U28gDng8ZXOQd1ZA3Wpf
yoxx5MnIE4HPfW6oH4TSd0it2cbyicweFrBA+KVsw2+56MV4t41ZVPEy4QS+nQ+IvxvR0hIBYHPe
NU+jNt4UfMoTijXRRI/sBaFZ9eNSYuNtqPyrJUWDxbHpCLCeanQWozN3jY2W5yRI16mwYlU7vEkM
Zx44I293rIdf3soy1O0jOp9dqr2DZPS/N/+sdqSqzoXa3jNMn3BuM4PRdIxhf3vR58Mriw9KyTKt
73Zx/PKXLDsmvmw6TsKb0xxAxnxCRxIXQEUe2gdbux+adntJaGMQV9rjnzLAsbGFgML4CdZNIgUR
niRsdgK/0F0bxw96UfwkK8MpyGLHYVWQHay1UOOlowPELCLxRpEuCPtwg73F4nL8B63/8toAiMeV
R5tkl80aVX11wdX3MmsOJ5CsJf3TKEvAsvMwbjzmEWRXbaajawusULjJn2YLs/cf//PS/+sOpbZm
H8RMRDPXtvaKiheMoM+lofxQa6i1sdUztO6kxORVl+IaX/e2q5X2Ed+JEuYOjg5Cq9hjVo930LAf
Ei0g2lR596WhnHAsiWaHUDBFmJRmig1KprA/Vyh6ZaZX6FNYutYq24rqEnaRP/WNaJwrvlvbE6/p
WKLJ/UtulGojGXmLWBRyQejgZZKWTfG9kICqinPP+IM9Rtyq1yQ4XxPR+UFBCFbP00DauGqoKf2r
RqNFZKvJxMLIo8Tij+/6AIkZ8F2Tpe8G1Yk6htVu6deUbwXqrcOqnlfsSgB97kV1oxybgw2dWZsX
eZ7R70Cj2Wr3qRLbLyrU9Gwil311ILlLW3LAfA2+fm59IV6421zqVAVnq5Tb19GLYky6B0ZxDmPp
MiUoLRTp/JcqiEmdIkL4J6PMfgK4quNL0lV4Vi5+8LH0+AGBa6/FdINLHelvhh3zQO8EL2x59+eS
1tr6pr8Di6E8TUI5X0fTWeE1lcN5YzKbY4Ta87sK3q3t7xYCw3/XZ+CWEUfKHV2LQArHeCWC1fRn
q6v6XD0nlA+mpOlACM8BBAjlL6AoFzYRXczPdJ+VmqcGljPnnh9JfIw88SR91LHaRwxi23Lg2cP7
PPCGRRnq08+h28czwZjRX09OY1J+17EJMTcVY3K9TCGqazd4E9qRRjL2yPgV8avJQ8VvZU6bH/pJ
dvlUOlhR+H2LhHXsP7Bxp7gxV9FMT1rdHwhqbgOhs9SGWopnEYvkLcF+y8ycm/RrhHtb8/vgTrp6
2RaHrYRQ7MXMo6o9PwhNkqeoe0P7lbb0kt0vMtpgZe15ge03zcREF/GKgqCGTcte2bnDGOCSvh6s
9HtMi0V621LBkncm8liecqZ89+ArIpir8QqWqPBp6mL4ZGXG7QGgEV19YkhXXgzNMkVI4WdNuZ1M
tycDAet69tucJKA2CtW3zFmjMmOWRE7YW4jDic0az2f5hQAJREFrn1yzxpwW/dpCpzNF51lFYVtg
ywatwgvRVymIRa0zUOWgYx3ii9F6XBnSJm03JWJSMk/O/cM/rQxDMv1BlSzayVQPz8cwJ65ZFOeF
VXD5FCn40wWpg0kG/JJoEmHfV5HVAjazSt0NM7UkIyHBkEGmufYgATU+PyODWv+oD2W2TBstuDeV
MR/fH9UcWXLYGKXTEibs5egI7OsVE0TcCcCfz4qPA3UznaQ+1wng2lvN1/Ud41cy7cT7Y+22Eu6U
yfeFQjuWpJzDu8eTmPXsjyKn9+sRUO/DFExVmyKiuHxS7G84/LvB9ZCn1YjXLthSPr2mbRm/D2VV
/j5a//y5mMeog3OiNs7uQarUVm7sznoSBFeS096lXmRoDnn4EoxHvK1vgtYk+PIwJy5n1AxCkHdg
7nKFwfoiQ3+8EuvCA0MzaqyBcCMT/d668SzW8GwlDhIsI1O9KEM53306qVrMdx8QuKZSBS3+RCXD
0UU3R1Lnhf9Y+/Hrcyb1722hh2MqV4ydRJv/HLSOix54oLyT+bEFrI1Pu9iYoDPlIuKMCHM1FMyt
kEr/GcN1osdTlTlpFR+5E0aPk4lPYK8I/woyfe0XYQ3bZwBXKRN4/k600kGYPeA1k70S8K5JQ1aO
BWKbzdD1r/7E8RILYGboJ1WNZci4R5HOhv5SlspVMkX2YQy2DjTLhyt3tlrj1Ve2/T7XTMCT4Ldh
+p49q6dNx5nNzxOPO6JjheHleXhVlK4vQeWRIu9eyyYxfwlzGSN896HNXhGwmjclUd9rkrwcNjNv
kAGICA0VG0cj+jvH2YbT3HmOb5EgmwZhsZCtvNmcg8qqvC2u8ScLs5eaxl+ER3R+cBSCGAZjjb+4
q8YVAygn0Z8pAzp4S3w5RsNc3ShF7irZVDlAJY7y+i8zixM0sv4OTidq3QvSQDukoYaldA5xr1H9
XCDHZKgQKJTlf8CG/TyLquQErUhd9lDcYhwt7nZdrIHdpO+EQgNFJNDQvsuCf+BC2Ydq63AAb24X
Ss3JXMIfTdeTdTFW0zlPmM2ZGvncPIlWNklI6HZl3OunJFmwLyzjYQnwqf05pyL1YUMXbjXVvpLm
1jbirr1a9i9j0qwbWP1HJbBxrjCIhSC3k2d3eOGiiMKFKhVrGqZrR8KAH//z+XCHS2IfF1VSjdtV
Di0+di+B/ON2AxEGXWBA/ZVAkT565nYpa50VItEoDqgEx+oYCj9mEIDIP5xNLdHheAHFlXsZfR8h
FdrUlTiazh6vC5LiMUitLi0jbHdCdJvxRrSzn8s95zHMXc28WZblbmzKWKp5XwFf+0ZnnavYbZbR
dxYTttFYOnt3V3ds2fDVP+qghd+hU1ussDLulkd0tl2slNFUDPqVYkwtGRrucZ1YklRID/8OIyjf
HMGCUqfQPYWO1DCwCLD4uFEs8iI1VUMY/J/PZZwJyFXnP1vbOfkkr3gt1K44pcK6LPpoutWcsQAP
HjEFgIucSCgpCguz7foDeG3UtQBu2KFnMYNCe58JtzeySnseGGxe+kPZkTCsnDjxTWIHZhsOcPIi
P6FCBWTGVDC3LQXZVZA/rE8fOF4TZa2sDCDxt0rRT1uBPIYNkhYRPbvv7ieZCj4iHg0BvfxyJDnj
7EQmYQ39u8dOVtaUJ13mIihUAwjq9xLXA5i0OsgDm7qhgdSZHKc2LMiGmapprK0D9UqMSVXG9DUx
vVTeSvCp9VlZ1lr5XrMKbhmQhlPF1x3b4Wzn8UkFzwuCM8YGuGFsjwxaPhixikfWYGIpgCnU5Dw/
yAFbI4G4UHTXnru7y0TD4ksBHuYO40SETSTvlOPXVKs0EjJJmFnCRoDf4X9zM6ifWDQtNVVigQhZ
8U6DzMUJlzZ/TnyfYRgXXS5xseQ/auj0Sbdn9wpsrOj0w/o5WvUc116xSWoMSv//SG/1FszDTFjc
zRv/t1NWcqkkOEpvVBNn02HpjtKFVHdvmSSNyeDhAM5vMchhsd8YsRK1giYfnQue8UEEPUZS0OWe
9bYl1vqoBAYFbDcXOF5b2FTk6PZ7BMcVh9kqL2lMujwX1BBWv+a5fXx1DX1FlUHvpD6iVqgej1PX
JRumVkQ6103U5wGHotGp5o5kG8f89nnZwVaKBe37c6y4wo7V/Oz72nvZL+O+BsUxi8tYgWMr/bdS
VFkrck2EBak5U4wQP+BaSHOmd1BeSFltlXGh0jLmyGElAQ7OKy3shlKxqN/8E6dSq3lX6/U0smmW
RR9/z3KaOMhrwOumyiJ7je0OWe9XqEDUoa3XLyEQse2ERSi6l0vyJiPxOm/I7ZeiIsBn4eQashyt
ZVoZsOlyAHiqLAr0eiW09Sd8C7AbBTp1SkfNRdNRgshttwWNnyebAEcE69Zh0RUARLel6goPRdi2
FCeBWYctQMRd5UNyE1sWOVR88qhE7VV4NwMnvWWw6b5jd6JDlbAJMgJeN5GRFSjA36Y8kZjEzukw
Bf3G0KKvK2IUZTDtRJw+dN8bCjOBw1QnnGFtxnqwL92mFByqpLpMIGW9k47zdWnZec79RAmFOJQx
//pL1cOHaJmaAGRZ0G1KrwrXcuX5pW9k2YA4+A8kqGdhOYIm5mM29hgHo8H3YWAtlmX0TLZxM/a+
7JHN+QB8tmIzfWAr1wB93w5VOE5PKByHNz+9sWeOVRzI/2R3yKMbNMGVhBm1q4UTIeQqPz5HaBet
C+Xo23/ayMMi12qxL9Dhj8qKyIRfN55wlzg6y/G6fLBZvQ/dddcqfLYVXG7B+82bMuXYbWXPyBNx
wCO3CGtB9YJ97QCvVITlBUls/gxEwR+1/W1xj/3JLC4Spux+8iy65WgClyJ0z15hUdTw0R4n4Cq8
QvmxYGgKYLlb0UvIG81s55KZhj2Y4ts+fizNDkLWljiapXIK68tDZFORyqarnJlTCkjkKXtGzrF5
awFJhaI/gF1dlZyk9H+XCaSwUf168WWSDUmogKXMj9UUUWUK0QPbewaRTVzIq0QtPju2AnPkKyNp
eBpu+IAuMIb+cOurknskvgSUYEtJW31aPQBy+9sXuQ1CZyWCCplxx+Ge73K6IiJNwadPCpF6N00L
vLZ2R42hgk0Wpul8Rk2Um8eYW9yIP1QPdu1wcDwkpWyjrgDlmPaAVt1aHyMncZ+UC2l73poH/q2S
82xEUnIO1SOU3dlS9TWRwYUD4JL0tDNcZ0WJmQEEoSjXexvBL0i9+sa9azoTykk0s6ovxmWtbXEK
c87pBEQqlb4/hy9r/EAY93tUib27GJ75FgR9Yh5b7vevgSFzsnY8SU+zrVCoNPcGV9pPt5aoX5Gx
pUWo5Y41hQEUX2ZzEoDODKyf3LlQ0Y0t4NvxVvjoH/8uViDXCMo2jmYwQGfAG+oDCljeFzTzbjeq
Ro27IwDns46w0XLq2RE3RO63rG0RUZCky1fO0+Z1r/MaMkHpieDttv4D+K+bwdUUJeU+sQ7Z/y1s
3oIyc+rppHHMo//M5179bTytkq7MM8U2UuNIUgJkgje6mzvjiamZwdwYekjuZhBdRO/Goi7Pkn24
E5nfgtw6Jxkd+OO9nv5ARiW0HA2IO+oALPM7zOS/CW5dHMdLJlt70kc61Xc1WUcFQjINcuKa5CW2
KTK4MbW3460+dNf/tfTaVsjHpsJjmheyBx3tN2bjaU2/HJB8M/OZVM2Q6qehpxk9ZfcsU3xmAt+x
3P8snZpvVQeFASsYAV0sPoC+gHeibKTNb/SUVejqXtKdYMcQiF5t5JvQB6cgg8YG7CIHiV0FRFc4
SeX4pdgPf0VP43Likl3m5WHNTHAiLuvQz/ajv17NMYp+YqlioBtPdNhN5nPTHFnRlE8KX+l/bqXJ
ns8mT+Auni9XOi7+TbtLNHkstM2T2cwC/H+/9MbBYdVmv1ZoSw5aaFeNFvXGUOw3NXj55cLV/d7e
tQvdCsFBkBzxK6jwmM/XBYJ9zklmcltp3A9syClKK9m4S4HIC8myBEl4zbeSMkwvQS55nLOrEdN3
/XghDEo770VCjoocCdiRDXL722cPf2TbJr5Vk1EkyuRRKTsBDxOBe0Qr+yCCYdlWFiHLjjNuCyoL
iKZPf8jj+aCQqnNSOBq+9F4FvLfi1Vkf5vC2jF+KgXx4RIaxefgnRfqx0mfBKRktG+d18ZFaGUki
Pk5FgSdngyl9uMKRFnCQ760Xa8I3C+6PdAUWsy6vvTMDSTvHdKiTOtubxBsDPNTU9dlcb2gbApBl
9bBPrc4qHu2RR2ZQUcOWM8/Rjr+ZoojfRrwBWDLtifX5np0FvC8l9bqTONejxKpseoAkcBdLxYiC
owzuJZyD5CI7BGRRMVRvmP8WHyVqa6OEX4J+djdlXeotqKOIDzrGcp40Mo0zs6eCawYcmlWhd2GM
W26IUzCS8IFHskwWnBCanCf0wD775Zg6pqoSTyzSdyx4gjL4R+4rRzxe5AjPo0Vo6jptO2SfwTq9
ewd77GBopfCMt5aqFiw0FTwmJerOkm5tCCwio++txUCdSe/drO+qVXrsmH/q31fdjbePZkcA9X3Q
BUHd3ErvJlizusUw2veQbWpZSo8Pg7eYnXkL0I6n+ILzL622WJRgJSVLZw6WfFpE18GNdVRMEZvF
PLgJpLwzmAMYkqnmywMybxiTxmxyb/4i5Kxjjy3W/9DCKpcUME6GbmmgKEoEVglVDgUN9Ev555Xt
4ZwKUoRvuxYHAxANC07s0519Abx/8LYeiEsA2Xxrd4J0rzn2rD/RcdaMxKzIlLGkIMl4Xmr2a8Rg
p2LWkYP7LGrEJHv5YQVPylNdy4AgDnWwcWNaga+BW/9hEelZR9zbEN9VHFZ6PQY8Llm3OQAkb86q
NXcmr4icaMOR9hgfqKXxZvm38toBOQTZztqPSt3Dstt9JA2yXXJOmayLkQzNoR+Y8DbH7sMOmlTI
dPWcMfFiydOzzNtjk20GzhQxqO+mako67RgI+VoBLZ//DjUQ3cfEmW9E2QOZ4U1lypwUkarq9tZF
DdeRVIqmAifGtvc7CmiVnoO6LxvkotXF+CSGWzj9WaAhGtOTDOM8dBr8yr7HiHgAoDRg2SjCOgv4
bDvnLRk//8T9P/AgnLqGf7zk9UKp8KdDt68rrSUCZW8H+8mg9qG091QdnqoVSa0Fij3YizrVm7GM
zq+6C+NngB4E4U2kvqG/G8n44ks9nMhqfmwfE+BUfj9wuVr3SHrgCK2eqRVcrHV6KvbmjNYL/mqI
KKEV/+aOlEAhza7RYOZTj88UDOG8PQHSFNT84yXeXRGW+AuTDPPbVhmA9WFZlKYOWduyCZJZHOm5
sEQPSiY+7u2NzPMNDQTUi4yeCibb/X3ep1MGKc9JzI2rYxST72MFzhpqCSf9/sT6Q8vf6c36uMEe
b/eerPU2mSmlqUU5DOZ4aOnEAVRuNd23IoYFYrWxFQDkghmUn2Mu5GNXIyej3ZYkmCDyMvcEpP97
LR321ZmosHwxgRuaeOXQjp6+XGNQEbc5yBXCY8/yzEMt0drDAosRUPUVKZz9HLhHVSk03ST37fzE
HoKR2Od8UhEocOcQIxMmqic1qeLoZW/b6qLyVAeqRGiAPg7iQ3c1jm4txb+oaNe3Slhjki4y510C
PAc+JyE+3SAdeUZVL/pGn2fcwHe6BmikKG3GlZykP+0Z1iuoU9feDOKRbfYyHgjeftuuNmicqbVR
l06O8F+CDKK1PZk+UQs+eXw47O/bNRUMkqL5tUO7Pqado/t+aWgHOfD882Sp6h4BTfmnLLyMA5eR
l9GnuLXuMmKjoJ/clOdjJ2cRd20f8drejRi98oLHxrSjFh9B3fiStlOFnEl4vcbLs//Dloqr5VvX
yUYsjd6Vd2Zfqnzddrp8H3azZn30/MaqIT6YKihqjg0UA8DrEr2IOEjHhEX8QWrYYUERnIrDqTml
iMqxQPbOj5rXWNVG+ibsk2tNoE80vzIlt4GT56KuEBIVf7Pu8hPdlbJCo1Ajz8ANYsHBpxrHsxef
Z+oNc1qOeOCM8vinn/ixtowpotDU4Zl86c+C+M6xEyBYrZN1d7riZQWTPs9PGUCgkjGGIBYTmTdq
EnfuTL5JdWWEnsAsc/nmj2CHy2Kw+hPD5pxQrnjE7ghgFoi2qwRP/EWJ3rOvLEStL+H7rWVnLN2o
h+rXQBV6Zmr3J6p9Ijc5uPTkIlevD0fzeizBWI1QDBZNWX6e5//033BiVrHd8b118CMac2m6vEI+
/uXCY2ln8cgULt8Lc6VKj+VsVxzFPv1n2Q3PbLt0H6RH6SlcCMoxyrm04VGV8ydFBCvJSTAid/K6
sO6rkKWHRAFOkfs+QD6jWEpAxA6opNEtlkQKYcmcUPy+QL5KXHjJ4bACeW21hySmS8sQx5FXQeVz
WzxcvUw+ljUwMbJZcTmK4VMpjtadPeWfTbVq1C/bLK/I+lu8e7YOW0eigajZVQOm1uxm/lQ9xUOE
e23vJmhYI17tGTq7ONfdalJ+mz5viVhOd4l6oFlP63n/p5/GiL8Fx9GB7ZI4XQooKMKt5OCQhAw3
tcr8wjfdMSUi70bGyhtMsc7V/Dx8PR9vi0t/xYR08eNDYRZ0MO/54d/3Sy1cZI557OFE2b1J564X
SiwbwJq3JqsJZDD5/sGQFNnNQ7g7B/d8VoLjeIUZ5u8JCYt4z7DYkm8nq1Y2gjuyYVCyI2sQEvrE
7HoAi7c2XirfzTbitVr5TqjQ2VryA3nbXlnJNIbsfZLiO/e2yNHshfhO0D2gxl7XOg6MdDoI0YoQ
CV5l3pgXbx72svJLmOQT9gn3KtqpKb311W5CyKGkw5HMygUBTdLOpmRKg9ZPcbewi7ftYfsR30e7
LKADQmyeRdppVsE7NCQkrB+e4VdVjgsMkegcWCX8KBguHQ3WKwOqg2Ps5cKURuVskEGaTn3pCVLL
trbZUmc3e2XbcvPrd3LE4aUzvVmri85glllfg6TwWkd9fNo3DajJF+/CmLqjmO0LtE6WVYXoazn9
VPgfB1b5jMybaCfyFHr4LXARhsSEFzifi8NRGX42eE19tIET1Qv9QBh/YLjlGkxl1tU2k8erj3xK
31TeavB9FBtxqW16uoUztiCewvsqFICw1BDP+1tTyIjX6e0CRMEF3yqMcgzaGCt6HLKPm4kDFUVg
ch0ntXOT32DtXlj6LFBIEyYG9magoC0NibGcA0in7Nkw/OeQbIy03qekBiY5/9RwVvgVitM41nB8
QJL1zSB/fYDlMapZrTnlJFl3n8R0TH/n9KGzNxP0DO//M8qXVrNKQFI9D7gGpCRmIkB1NVOUYvDi
doWfsonfplJRv26DdiNtkyGiSivU3Y/870SkQQEfqHqpSLX/7fa1AFC6hgq8jJeApkz1N+CAeDxk
LsS/GMzhz+yHR3H6nPjhZ82TXox3mhF0sNEuKdl0Xr9AY/gggxSauwGHUmP4ip1qo8n1Turk16ho
FepykCgT3JQtWD2Mw628wzrtAiyaPLh9W0Bpk+Gmg+FjeMLFPqH3UV0zN3JW6P3zvbbrMc264a7j
v2SDuJA9phv02qFHJcxz4YySzAcxdoaHKZ/G6O3EwosBeDAc+IH4L3VPm9icAhT7gYdTFwluXXoD
FgyoseORRuPRbCGiNie0trBMfmzW1iCSV51LmmRBzhe+/th6Pane37Fg7vYPlFfHpnvIRk7ExPy/
mg1JHch/SdxPttPufMiqL23lo+mIIcDTuxpMtx+1N1d0H8Ge6s1HxuEcQyazlvn/B4xifSb401AG
CUylvoWggIFIuo/DdDFon+m+9pf3Lg/nMShuS9Td2mgy7rTAsO77MUceTK+jccALTkCMEAY8VXma
qEiD3YOOG1JsJ1ZwcYS4qRCk6saTtmHQJfsbJDJR9B3+2zHw0hfatMnGdrjWmvW5Pe+jH9ge7wcs
aYBHkBYcB074J0bBBYb4dnMd3uVKG7r9A3//zrq4NlUSMeiPenCmX2fX7yjpSVoZ3Q7u6Tpz7iv6
gqyOKKwCBcExxx+SE8VMLiQjthANI7JttcnprcGACsiFEgprve7PnmBxrufnkMMmOnSisQ1YxjVy
QHGMY2xojYANZM1P/g7dpE61HQaMEq3Ho8iuXewpiMhXQrL6lLgV62i6oGkn4aWeP+vgOLeORXHN
DGC+5bciFKZs6673jNS1YHUx9ENpKpUZqdLUjEaTkMwU7tROIMbfI7g90whjTqsG82Sq7GX/jrjC
1vbj3ebVKoP8rj+1qS2k8NyHhpgwMRhqcLMXQpbWtw/4jQvtJCrv8Q39JrRQAOzOxqRrnCEGczvN
J7v2ABGFy7EPf3Z+or7JmKg2iR5X7Zh5RF3+Tp58MNZmUkRpze8H2Z53OhB5qoGNpB/PPtWnAdTZ
UBDdXv2UY94HgC8Y/taR83Wz11M2SDPHm2I+N472wokX7YoZbRzUNfftyroNfcOyFntFSM2Dkbuz
SlFQDngvoEGzTYPjmv7fKb0iu4etJQ2df+T6aL4R+ZaVTvBWMXzGh37JTB1PbRowTKP8uhTjinDW
l5IfDuxtogze7Eq0cKEgIH1JrK40y6Bhu/bCVbTO+ySXWwiNa4UwHILcT/p7TNXK6DDcl7N7n91O
3TuuE0ozDRggZdNKtN40Sbdt4Eyc4c8AFw/ukBebon9DMASyki7jPjrkfAs4k9ipD/Z1ExNSjWnS
UbCEqVmE6gmOFZTFeSEtgIZdsrJCCcHRIaB+IyOkMW5z26/FzMEfSxmDoo/BnTb6vdjE/WF1kZYR
c0Pt1O8SH0EEH0L7en8vTlm/8bGboPJyRLkr87k01ZtQMT0J1Rfi7rjqzuZadA8mEJFGrENUyN78
rGWdslYPWO3iXHdKYQ8aXYvZgiM2XuKxHwD9JA/+4mpCBnM8/j372yXOu976A1tTP58NgOogREkc
/EhD0M2JGc6Gqodg9nHDPMwh+KNsOgC366lsYzRso988FQdBt9pvKrOWT0X4XjvF1u4gqmFGvyMw
kOHf5cpa6cDMffTm+yZ/mARZhEbykveuc32yLbpRMLGOOoS1krMLZ04qVTTV/VO7BdCBltjdRIU7
ltY3Vw4D7p2ZDJ4tnWUsJEv+M1r8aFNfhljPvy/UiRq1N3IBpRmIFr0L4jpB//7lJlkPfJbDnSgl
UW/D/jNQWuhQDjh/hVaEr8VcKV/rltpx8Aj43l7ReXdUV7qPiBC51H++xrvYOQ2UcnO4D2in+Tx1
C+WHRwqUWSVgt1XGyqnyW/ANmQ8V3W3uxP687DqiltBBP6f0D8daqRHfeZ9fbr92DqM4myDPAeew
0P1KClbDBi7Rs5uQnebw3wIhSFwG4WI16GvY01Xcy3dTH06wlAvLPNad9rMek4gqiPqxmD2rxPEC
pktYReEi9DORnkDSvjhTK1q3kcAGHKhOejNHVBHXEz+gEudE0O4KNHwzBlDzQE0l7HWEruzNoXn8
NCoiK98kZPBCW5K3t3Cd/lDGIm1jv+pvhRJLoPveYaK5eT2FNg/0tU5djvzQyeGi9hBHo03WZY1l
C3xS9Vo4LRjarimuZ+uQNIHHux6xg1gjwIeXyH1QseW8ZmyKUWyEDFXmzJ7TQ7+F/Ui45zPDNSVO
zGW6cbnVtjhg0lvjQwaboGQd5CoE6TRXzJuNNcRGejA7ntIjRRPbJL1oe0fWS1T4I51As/qmvZdz
H6GB8H1vtWeeccNo3SjHyOgMiVwo0kHbBKA8uX2TqWtNDYWhXwyRcjloTlSC11kcfbwApoE3zDnt
EoCV1guP53vhu8GjD73ojaf34aWnTylBjhelD9r9ohpdCpHAgerS7GZnMbWKhQenXuR4yAO1wZGL
k/qZVqhZazW2Ey9EMkLcIMYgsTHaGzZHH1wnfXKB8FyiJuRu8J6Fs0Op/DrkJKJPVBV1MispjHfD
oe2rWDf7KNkjsyfNXS0miMaGBiX1PJGGgJK008/+ZBSeNi5+iuWu87kfS1KZiDIeMh8OYjUx/qz3
81Pjjb0rsB80YJ+5Xz/jO1NLM+G+9oNOXJl2eNss7Ar9dJOo7zzt/1VeXIQ94ZmkbiA2/84WyJh+
yRyrx6f5f5yzoZIAHagvbx8trnsX/QXFOwcNbcMi5fNCerBpqMH8ZNshYHUme7+x0nyVx+kYUAUA
g/Tv/sQTzg+RYIw8dGaJ5FJph+YRqPdkwQFJ9ocxnk/ZZq//eCBKvXscd9/Z5bgjk/tAJwbmjedy
wyE4tVibRFD47Gj2RolaOdQhUuni9cYyFthXm8fgUiDt7nmWnxZZb370i8m/6Z5F4JLnK2m+V+5/
HTz/2nk1q5a2b4k4efgK9CHz4DPVye62AH+GwU+YLNc9nkuzBt+0la8G6Xhj+VV9QFvtmhkk/vvK
klPudY0Uk2Gbz2RLeeslJOgon5iQP08MkI3KuoM7sEGw76VcEFtciZdrIE4etmVJHuHC+8pIQZb6
yJzNMLO4zlf+ZD1o2SkAAj2HPpDD8BJKQNvKHYqPKZnqosGTZAvGYTG1wtQOq0YjkoPyo1qH7I66
rq0V3kUp/LrS/s07rl0woEHEvvGzSUmIB71+HQdCKPaU75nfpXqXOJoFVOmv/vC9B6rZqdBnIMVr
Tj5T76yHK0iZDpDT7YepA5WMJM6cvg5ZC3Yw6ppThJOSeBb0/3AByirz0cECsBZEhCjm9gC6vVQ4
DypBiyqAr8Tsrru4ZeNrk3c/rYP83RBzZk93BBb4rF7W4zBAtNkgiiqaO0V7i+O3+5FEUgIE2amg
zwoz/LKLmSctifn90eR05khwVBkrcTB9df5aObMZhlV6ZGOQ9bMNTsyq1MgZPoxk+AxqMK2DnsCj
Z5fMkFYDzKkFNidqBVrwsZQMDTfWRRVO6aDAAjIvnyZgnGHBtvN4y+TIvVc1KgngeP5eQobOcQYh
GKIJtu8ZifnQPuFYtMvMe67SvaoNYfjGsfh4wf/f/JTqabNCo67jFAIuPiit8IRfs+gR38TAx7Nx
1XVKuIJjU+1Oyl570DDmU276jNQqNErGeK+xy6Fi8vqjJSt3Wds/R42Pxv12QZ32nQRTTwuOSRy+
y+kqf7DQzs1tKx3fMZsMr9uyOWt1XRgq4F7Oo6YY/vTRStzgEhE2+1TnLfdvaT6ZlebbdaSlPAbq
t90tieRLVA2LFF+RAMQOTWpHJPnA1+Cgk+hbRsTBgEbZJ9dURDBFaZM+kH/qiDna2VcAkuQeLSo/
65pZ0jInjHxoaljAC5AQjAMkTe8DycQVNocoADarKZiXPtqfyLjNxmWHScOxcIQNlT/R7jBIroc9
kwlaybZcOqwSHI6WJQ4ISAf7cDbhZATmBE9satqXmFtRxT3m4qY5iEhm6UmANINPzwUlcgmhH/oq
oknbpHrKjkMdCkq8V5i8vzn8mvY9vF54J1bHeIsWrkvfXSRdFOCqlWNIVcDYnJHHvAQw27D4s+sh
RfaHYl/PGBgBKPMifVNsjVqaNkCO0sTUpKdRu+WnoV7XN7iYmUfeO4dULwFjhG994Re8xkDvl+LC
lUw+g8ls92EMkSxl3yBoQ2E9UIktlgsRtOwMsNrYSg0MgDPR8qEad+QPaieGaPSPnuSwlRVTQuGi
3hI0g/FsKDPIjxbP+ThCwIijf/FSGo6nA+gIHnce7u6YJFsZh2/kNUNtg3XpJfdF3EY4bndMP+Lz
u2KIh1U+HqE2B5WX/nYk0P1M6GtL7hIFfgHhDypKFc6FoiPIAyotCwSsVg0Ka8zNsD2nyel8v8bQ
0eLo6Zh/8Zg9R29tt5/7ZlUS74vDOLL5hIunKVyUko4TXn7Yezlb0UwYtsnpvdUeXHjUgskXPk8v
hHkhc8wzC5lPuwrS2UgrlkCzaOCPofGHdjBQKjg3YmNi6cYUEu+Td8L1zPqAt6S3pWcX2t4AFL4V
fu6LD1YWlEVZNzfJ9QsprEG+4w3MT4Jou8hFIA4VDYzJz8LiEjKsfDkFTOUS5KWi1T/D1Z6SrPxR
DwVLtxp19veWkKWxsu1tSi0F53L/V5WbD/FU5Wn0f0wjtbrrqSf2eUIBEB0fiqKZrefuaYrju2mX
Bjlqn+b/gP+qa0uAI8BW9dhBqjr5l2O2Vmf8fIiNFj/NLRvId3E7S6l+AXJIOrW1OBkt+vpG78Jl
0nFgcPxCcH7JjoSiIW2ybXb86oN9i6auhKCWRxTGgW3ioFoW9lCUlWtyeOtAh41w03HCvzp4DNUA
vMV/I37r9ZaXmn3hpfMwiYQHOl0rNCm9XBBEZf1A8KF/Cvl/NNG/ysmcca82lZdxWy7MGx+CMf4/
ZplykRwoCynLduSSNpdLpPPZFYMSE82XQlzwSVs8ycjqsnopnttuHfP3xSmcURWZ5urH41AKfH9z
GebVILBYWvOtt1TC77rn/sU2p8vBmaQdVvJYqY2A5W+JDCBp8heVzTU/thj9F1CkjZKvUORqaQ6M
aFncB+LC/gb8FDb7dntfRGCrCN0ae42eBlkfi4bomniD6oDOcFcykkYuEXnCzMDPe45rA7BsxOJ1
fOyR+hv8PQtW9Tc6ztQVZ6zLXkHBA56OY5SmutTrAUkG/QbHVg7rDzmiq4O2fji1PdQBpa/vaLE4
rOU9UqjbUVY+51uQe71f5cvOwRw2l5bdeTzSJlLx9PRKexicEHWu1UOBZknkseVtOQjngOpB/DeU
L0RKT47wp+m61UPFe4fvDqFluFlDAkV6wiagZ3hhANAe+F0VIlO3QfLm2pN4WvrICxYkGHsU1cBF
ohOpuhIaBGS3Y4bfNwBKy9VxJSK6S1vjd5f8QVeTTXLbttIWqRt5M4Dj5DVU2UU1Smt7VYzo8Lel
QcI5fHFTKDL/St1WbjeH6ge39YiKPunytDSQeBOlehAfLgVPQH4tJDufQpbE+vk6UgUL9FoLB7hi
oLjpA8GzKiILvvdrifPe88xAZWhrXmFQiFBMpJwnOYygwADBfqYSk/NRL22VsO3InGmL+fCYE1Tg
niqsQTUJwtI8yrh4ORvpRA6nVzMGF3ZFI2G/I2fgzyIkBIoYBSrfdjzRlo43CjF6TZ6hhgJoHvh+
J+8ZQDs1q8q6zywbWTBRAxBJLjfyipBwRzUW24vJy7kg/l+RrIQhTelo0p5J7u5mv+Wp9+LclDnY
zKdwFP9TtXjgY09DG8DvNC0h44dGPrv9vIXpLa7Sm6IDKgGDPo9uq5yrnI2uoYrRYXiV8L72biRf
l23lqEP+peB9dsIgKNSoNPLBgiN/u4pqpX6tSWVbkK7VcnLwBOT8j/W0e7NPiJ29laezKWC4OCmo
/r/0JMbIkbWMbNjZjTA66/FKqbnYlHzzWRt5/znc8OCLsO+TXp72P4PA1LFdtoRW+ND9f9zHy6BA
jXBA2Ga28Eo7WlEmqk1Jy3NMjPsMyVbnzVsr2vWbxK55meqpZdJTR8W4GefH7Uc+0ezjKUSEPpG0
qkUvEldnFEyPkfsBWMd/aQ5LN626RAXEK4P5McFbnceChuy1Z1fC5j/0fj0lUjg4ixDy8T8SSJVi
SE5YS+Cc1a/QqFZae6Pg6jvBnvPj0tGG8gHdHJZsZHLJe8s5D/pxoD88Mb4D2hGDtjl91AIb/wkh
PgMID0wpTKjnUPwMLY9bae/Q5SWWRczM9lLWOKtSOwAwxnLNzfs03oJgtd8dwEMeVTfl3z7B5yqq
9aT8a8nRoYLguh6unX+llW0NVuDMubHOkL7O816OyUIHeKky25pPdJEsOgePGQJ4P/pWENpsl80R
XevxiaEqNSBptsrEYjS+kMco5OSObPGKmXBJSxnD0stbQmSqZKW5ng75J7jkKSG+UeDcSe8RnSfu
T/DCml5xmLPWuoZq/BTeh49VLyHGNCjE1BF0hCYUmElzXNy7wfZqx9chK+uQf3HgwLsejwh4l3wG
SNSbBIC2Fofeo3b/WDJzLBfF/RAHTm5BRz3hnt7sXLNRiRQH1d2roCemiD+rEl7a9168xuRBPXQ6
2ZG/pYjR/QbeXzIpbeB5DqgO7avo1KPmLsfjge5ktWPDDvI6MSjUiJmhtJb+bONk3HRdDNlVvCIC
mAPxj19tNZiOLcojxF1j/fsuvZSpMiWhesjtFGfJPrN61rH+ddwNJItm26p5su/PQFFD4FFcXBGd
okaP1RzuToxJO/GQ1ldoCjYfioraw532aJcVrCNnG/0ygcgDWiSU1cN7D87MQLt87atPp+04/iCz
5LTMcJWFq/LvTLB8iHCQ8dY+6oMEWUosDFTVDpBX46amm21Zo2U68Eauhkj2GoobCPTr0oK8WmhX
Pv8zh9W1O9+9EzHvbOWgBgYrjKeg0T5YSh0CeUfSZsqkKLfzCRCwrqc3ZTCLaVf442nwaOGKhHEj
TQ1v38bMHc4Bv3WW8C6SsRZGhYG17p8DIjVTdN022meli7PyaH9YlZxfyB1LWXLuKqgrO9GvMimX
Cc5ZN5RGDsxrh30F4keXiaJVIn4kUqdYg6YOlTzS5EqB4niPE5coG6jBBtMRDqOT0aO3J60lwjbL
hmNmbEJB8XmdbRaoSzgmhiySlacbmynX1mY4CdbFBELIHO9L2xnzmwq4VWJWQqKaNEWm458e6Fp4
uCedG+EI+ln51dQNIVsTBAxRt1nE2gVVTt3C9GL6C4BKDTJPXrthr/rVU6ogrvlR6EsOBgNwjOaD
ZsnUs49EKOXc1rvgEqeEmmVTM51G7MpwLUZGBCQPtFVXz3VB+QADrDUyBgo7HfOb0rq92v1n4pLc
NyR2TInV4YOZUhSCQ64Bw0un0K4sOgOEFORIJmsCQo/b80zqJ6dNOXv9Nvvrp2IHArYGhbySMfGy
v9XWH5hZIqBMON8xnmGafgFywOynBy6XmCbN0tP/7sJlAoo4pYwx5OYqPQ0S9iZ7urgz/2z3XWgJ
FG/uJDwRU55+LjFcJxofhWDGb//nIG6YbZO3WrkUiSHqqiypS0aVurPW41hU3BDDxZ+XT34Ix+DN
Tsqv7aj2ulhXj88Vz3o8gU2Ha9kkm637qgh0UcVwR3pSwsowZchBtSQv9jl6u32VXi0cZRg4bPTU
TVSFpX+Z3/gQ6dmVUXZTJDfwEg7IRXPL9Jh2PNAwoKsv//Dsrlf5iZHIFCBnroRmQQBfEI+XWUPL
k8QUG9TN+pETiM0tkEfGIwP8y316jm0lLfog0KwoxOjnEZNeHF5vbkZvdRyH869OJeffpVaWJcjx
KFOG1V2GUqtuRUA4LeTKkJysWfcfgndgE9pfgvnqkNsgVUxziSqyG9tl07PadwXjhbhbdG9ltaHN
OdqTksxL4iho+t+Pxmvw9OzXpG4iv+HenW0hPt5yygAvLk8WFNdUXELNp0j73U/YxuYsK2Dxu72f
2gQXAN6GLIv9K39nHDHP0kWAU6na92/6XOWEukFBf9FVq6PtwZWs1AfK/Zzgs+m2A9qgdz+QWGmY
7udKfRCfz33O8HvxiaEaZpJIlis8JyTR6ZdF1sG+nuPPUk5T2mdH+GlO4qWs+JFqGavrjTElw3wT
gDEYcarym80d6z59jfgoU1W0Xu7aNlo9ZLrLEEY45PzM8Vq21N/WBUVmEXCQukZVdaBlPvVl2Aop
cRoA16MUzPM6JAkXqDzj8aygPTRWOv1ZFxWVuCjdYacfQdQTgfNzBbYFnx/gPAKbSjpA0UWz9ujf
v1Tq5LkfBWgcghD1ekuxqmMNaEFbj0FU7rsqMEaucDZwNs/KNnvDu1YkDOVk0W5Xdeb1yEsWCZol
v1AXOM31lOKhV9K/J0x2oz3hY29mApL+EHPXARMoLVWlV9X4LZSDXF/gU4FObZ1yw88RsOxoIg4S
ZKTt9UzweYeTXaeac0u/qoqbO4QxRjSFOGVyz7ckIrCUuPWbXOSYkWqnHEgA+/uXirJ14SWSKaBk
xDv7wcbY6k6mk1nCHDFQIrXc9QR+gf7xavvbLdFR8gDJ42f2z8q6KOfm8fopQ4VwycrhXMSkXqhJ
3OvAFHc04kVBCCOtaRwx3KRN51vkHZHQYX46Yiou1hwMCEQyYvBjNdsfu7fTgFaTAocw3wxKdatG
/EeL7dE/IDAyF+2eD2nSqh6ZTcGCiKLCLwqoBQNVFr7fs5MPzWFTV2Nox3fLfyscb5cKPguFZkxg
vXIfGaheeJCXKyqMKEtpd3Dj2nbEtlryhgFgAR5Ftyd5BotZ8WOLQSM+/GnvzVB1eQuAKz1SqMyU
49cxZgv8RDoMBmZfLf4fMLFKKYSAR/hoLzBkGiXxUWarZ4IiVhbYs5UwP/q8+rfYh1m2fyNcq6CQ
Jbm1SQgKy2oUvOhtFzbosdzC74Wcuo62IdnhH0DFB8/kwUdPXoHFYRgU5ae+2XYcMZSX5TeMfs1x
lqv9egAh1dHmj1I18cWuZxHp3pV0Gu+3xYw1Lvnqq4V7nu8eOWK7b678vLllxv29EZLXW2O/K+Jc
k11EbxD1dIo1/LQCY/qxC0u1siKrqxKzksV3x8Ek4il8zcLm4jSkdOQfPYL4DEP/LR/ThdquYn1w
mU+2C5WTh71DfznRpb+PReg73/J8GqDd2xtABsZcX6KEmJbG14kZZpgy0X6aNolxgt9QPqImA7fx
G/fwbSlyo9hsKBv6ih1JED6CXgrr+Ud4r/balbkfs+tRAHiUGbArnDcz0QgyM8HhDMkRD6xWNQ9j
sURbinSuzVk1m9zZYPJ751KzHs5/wh3TwdKQsMOCfdnKQHjk6AynT3vga3Yu1zdu0uesp5MxF6lS
lkIPKNvb82E2H69MjFSjrftXpTWitdhUeTlo5XejLqWVs0w81C8Mm3D/v0lpLsc1blfLdrt3+vC/
zRAetQSY+5uWLsGzAmwldIvDrk/PSbzVRGui3nw4JzIb+u/qicr3rOEgLGsvbkbt4Pfy3utxgJbv
ovmfqUVpyaw1o63lEgIMdcYr1B0cN+/OV+5+7phaJ46FxxwwkRBBon1sq3zyI4xVF5j1S5rzl10/
QyzWZzdrp8WIvgPk9X3wrVw+jEPGK+5iXhLFtDOjaI4tvt3YXcMuIOSFHM+xnbSzqzQa7ZpagHbk
xgdpPdkeU+Z8BSkH53CSnhNYkyqwA9RIo2QhKoHRNFTIZTHVOcXdb7X5eHeGSNqL/3aXMDtuuDNh
h9NUfer2VQocqRJPzgMiPWJQi7FHjLymAAsUvpNqzB1xD/2FOdU/24PvLJA9FcSqdG0fJ+5EL8n8
cDZlA7lpRO/6lEfb6iYfgdSeEyLznFqLSJqbvHZPmSBwzUTl6QeaR1e8dpOu7jzzfBeozkjR/mwy
YQe2UKvrtfG4Lf42pGbRnxRHOitdkjD+g34DUDAVF7AsllgZNl/lt4Utc1OzVuGH/fth3vOw5Hkw
x0K0POkUMou1r6JcLpueHO8X3yU75wIp5ulqqgvXk2RG4iMMrIlKBsjy7z98plALrGlBQ9y7QKUw
X3WMHK8X9MkdtEFEyEw8eZl5r0lG4mOAdPJKERHaqBrpUGTUHE8eaZX2yO7pzBdi4cz14sKQlVu1
I0DrdI+IHGohV/dOTXA3syX/zDImO33ciesURVMrJqseEZiCUYa0s3Gc1B3V6VUy5qoVIR1kqDxi
rpv6TB1H0SCUoxaNdSF6PncM/MP2IzwFf3pxEjKKIttiQHXkKPSYsZbLLOvDh6iITNHN1gm4ZLYZ
JWh/6Ld3OcFtegp6pN6TiKZLoOhkEEJ4712+BuejKCcxFHURKF8VeyR5gxsk+huwn6OOtM+cKKsW
aeTFPGAs8QclKoRX+sJ3n+IUBW1sN894Eh4TEvY8T8eUqqWeqf2am4d+Y9UeCpW2O/C4OVSVDSbE
OpwXbAnezFl4+b2f5QhV8bK/R+LGrulJ2npP9FBzlvJyvQC/OzCFJk5rnG8ZoZefeo3UDHjoE6zv
KBGj3gMyrRNukkf2SY1n/JyMN5hSyugRukxJJ3HW1RoAwVjXxG3ECWOeJpvKYhdyY6rSCTx48+ft
jsMw2ZSba8zbJcrBW0TEu3kxWp4oRDU5jxwTwwkN3zQaGDXDTb69Wkaa2d19JwdMJv1jox+gmv+t
b/Fm9FL7zCd6RtZGpaErKPIXgxgw9AKMYzQJVoNWOO9qKM4bFhyMVd++RE7Daz/h8YxX+tleV6/b
71zmdcx2ZSuPOvv2HfviYHQ0nxD8Zf3ZnI6HjkegkzCVTYIdsf52mE8+/fWEfBoaiIb6braY+AAp
DIV12ZqAogy5DTLOtKKSviV+JYBqT0jgysmkN7XRShSfdkm9iZbr3I6yQKozrKsJd1VYdi3Uo7Rw
+xpcqnEajyzDlcXsnJjZqYjNo/glvPRuQasKvIbbsO4wyWiUVo3NxRQKpjOMYdL6fKuokfDPyvWA
xGGxGCdKjizswZACZr3CqWao35A9clksZLChB0xlt/dxl2Dw7YmHt0hulrIYjjv5MFo1II/TAoal
IL4fNqw55BzCII0KeqRkIChFch3DlRPcDFrU1RxpiievL5qrx4lqn6Jh2pFzdrtaEI4eK7ryCh+n
LiKhtZ4nrAk8jWKv8pLeQewgIuMcNRX4OcFyHI7sDw8iTDUG62PSrijO9fv3e0of82Mw6HXgxFNJ
z6dsgcWvCa1ECPwB5xrNsRmtmslS0Hz4+N0Zpo+PYjyVE54tp9w+OJ6LGZV8k2OMjtCyNiOw1Bex
G1hrVFi41zMyhPZsyugEV436MQvuix5xNBw2ErDLlVdc1a/2RX5oSx2DWFjpFlQ0vmoUsAVtEals
ArAvv0ojddynj5HqrfAas75JInsp8ejnrY0is1EuL0W0yeDspkR4NDLKJfFVF9fHyietUCkBpKVb
tJdQtKOtO4eP8AXlmakUdSM76c2aRQxh/SX0i4TNMa+AgI7AtTilwWiEisus4RxR0gRQVjro8q24
LZurqM353MgEk7DXWbysqHtiFMsB6+MOzH+2kL7vTqMQb5Snlv1Od/YKcfjxZ5u1M6QIlLwysn9c
z2S/l89Ri9xXpBKumt3CEVCbxTVLdfaiEi/HZFkPmsEk+BaR7wMamRYvCYvq0jXmVuUmBrFoX0+2
YwKOgYDydU3sMgNX2X6vLwFWfM+nLnV1uBN4xIX6Cy6zH7pC81qa3mYy9ORsFfWyvOunZIRhsHWl
iysqUGHNA+Z+QEp+GqXujIuUyfkrmb/m4qCe7wyZHKOI9xPuOUFz7ZimTAA5DiDCHtnFWVyLcNii
2sH3aPsRs+xXPLBHo8Xm63KjX9sBeQ2XnwjB5nK64FvEvEHPVrMzughARmNE5dYTBgVPcafCf2C0
eharDJEt8yh59MzFdogWfSPg9gVJrN1BiazwYcIXvX3rhRjqEI6KL+SazPNcHz1IGbGgTScneC7b
Jxt2omG9W+ZAjLWvxvrOJ+Eo97fQ0KFHGhFQ5/ifjVLwIT+ec+n5q5tE3g3aEv3RdM2Sek1SCBRL
5ajeRW6RRyk1EPLW8pJrqNCUvB4EPzhpqztcCfeB4+F3vzUDOjrsHAyT0pI5rG8wBClwITXOInm8
2Hc1CEuwFmF3AB/BtLLZWQK3KDys7slHF0Y9NHiA7u0ZUsSE2pcbx108nHuIOLcg0IggJaGoI/zC
wPgXCINa9BZDMm4asyvuJzaaaFXIXg68egrZizl+CoBBJVTSt18E6QsBcgNRRYQGQx/dUmyMEjzs
RSfVGG2o3K6oRAu8wQZwzwFqfclWnzlB1NrzfYx2jl58PwrbIAtX8X1d6NZRiBygu0kapzPRIq0L
NcXAs7puH4qHTuX69X3meFnP13+qgh4Sifqs/Yq/C3yz0yl9WXjWRaFheygQOKCb8Uy4YW7qHwX0
NB/fj4xqmqEei8KhJyQqi3gX4wj1oxUFEZaK2CGDhgWfyCIEyBd7TCCjaknq37tOPaQzWTcSqYsD
iMXimDKHtNvP1bgbGwRBihZ+oaIqtTNw1fkvZvMj8gx6Oh9EQ22FQpWt5RF9t7V55l0m+9wOjYsk
l625GsmVYTxdUX+hKNpSo97w5hfIERm5d9kSRgSlkel4LW6dq45Q0foknh66q6qjkNjvYeT0PTHa
Kw+th9SjSgQDuZpYNVqu4RJzEsRs3suW52n3LWhtTXW9LvcvWItEk0jQrow8RViBnEf5YbQpPgGP
rLnWKItmGRHjOGkoK0Y93paIYhWXYx8AmWVoyiH85wdCXpp3yvtt6Y0G3InITxsAs+upXiUC3xTH
7dBuM+kILOnQVsbfb+V2jSmV+hPRdY91DEiTDIMtX1PDYZz65m/gQ5Om6pIfFI9XD7PrSQI3qo5h
yw7iCK7C51jlXmg/yxDkZHyWsGFDrulc7Q4AUykeWCrUNmwcZW5kRMT8CAbfhF2YejU8MLZjggU5
fnA6Xf1f7cgdL+qHwO08xxtGxXlJkkj/LQP1h6lfVY2iHOD5jHRml9FIrU10TfIAzFwQN5bgd1Mi
p2jpJEAjvjz1lAvx3P3KANkQCFD1qK5yoUlzu9prVT15zHUpYltcQg6YnlCANaEUb0Rrsp1vJ0jb
LXs6x8oievXPizr5sjVMhWoClh4qqyXq6Xr/NHYGuCVxqiqNISFOJ7ii9GjZtbR7gRJDDs/jzirH
Eh84aCG1tSs19viravkVwgqJ1TOCkPqB6j3AG6IDw3uKKKVM9C0JpC60YAuz0LFaMBds/C4ouOpa
f9Xi8AAcU94VI2VsE5CcP2LVO9z/QGzG/KUMgnvhOGNNCkY4Mlz54/i54u9bsNObzdYTBiGBsijO
03tu6aenHxSzztYBcn9uNiq0qXu61PHvm+6gDVk01/CoVloWJs1aqEkNxbgKwVWLIMRsjxSSD93z
cTONTavgFML4Yl1CYDdTGWo+Gtg0jiiOsEVyTqsbRBxU3l7K05rvfgDCxpdRoUbPkQPZMhR3vrXz
TDht5//+lGrGTzOxh2mN4mdzsfjt2+1PH7+rOacxN690yzqY7uyntqoDiUqrCpayRlLExzDsV+ys
o470VXn8oGTdZ6mwgC9VO41KFbbiwqI1wY+uUgJnsxCloI5VDUvr6/f1qfCqzNcJylRq1QdQoeSp
pv+YKY936q5L3jCrariOHV5hR0UQ4+MO3XRenx8Qh6/MZ0+CetWcDMJBydk0qMwuGAQMPLNxD80K
cxx511V7u8czMTTXTe3WoyBrgoi/BzT5CJBDni9glwuREsklGkpC+T+HsDh/DOLXPY6/MmZFE6b7
ejiGUS5qPW7FjUX7n9uvoWYdHjKKor0z+aX0Cj5TH/qWQwUCMBmA4dl4DvRceJZp0Riyki2h9hIr
3MwG4wi+Rwo1dVNrAvdHP35Y9mzNuyesoMhDLrsZHwoqOnsNP2Eyxm8KktntSGFUosmV8c9c3oy1
daWpvWBOo0lOhd9pH37HFLttLRITjeu5Cj7BIaOaghsnfELa1w2SnKBcSIGXtnPcxspz7UTrexdp
njDd9JX6rKafrxEr5ERIDM9PchxwxnE0IrmUqhOXFHQvMefpS+1qmoYxBveMAm4xUjiWCGzqrQip
08SBE2/CXTdLybNmb276cQyZiqsXQClaWkEYTOb5ffeh0PxvFPYUeG6er3OBhz1pKGemw1ceMztp
mqQHzu2avnl8PnBy3oojqC9g3tViZtYmUZXPsUxdS+GBeWjqP4rtOjCgBGoJhbXMqYl3vJ2yCPbq
mbny44UYes7dLozjudg1VxFlqxMltiTPMMpoI9v0OofbTUR/j98ZPPpW/P+tQg/Lh1rL/eKk7qAc
lwVaRKt+4Vx9dXUG1IpTkfWiofB9tX4QnRTZOzorwpWM2BFrw3mhWPzti0fln3adBrtN8r1ibyeu
1DZwo7mf985OyF7J1wLpEe1o/E691Ri8tgx3NyBtch6sUNlthUGhUnZkoSLVbWuojKNcE62TjFVg
eL7m/iR3YnR6Lmabvqgx+p70G8Hk5oqq5yU/LON3AeqPgkjGBex9PKMhJS4Ed5AYaJ95DjGbpgFT
PC/DIAzbkvGpUPxaHNRDDcAvfrcuGql+dzweQGmzAgaVAHQZHniDnLgZyoCmUUgFWqWL/Jrv0iOM
dWu6TA8f+hLwcREa2QSDDF5DFLLGeLUbtwHnsDw+7KyMcng0QYd8tQ+CEsPAlC88ZFTwjQeU25Hj
2GIpXS+ts6CiiRHXIRy/zJUFHI1dSf35qvub9mw4WumIl/3ciGb/nLxUjsGOYEsU+4bmsjjZ1s0h
RB7TzUf1rfFrGconhgzqLJC5MyEBtwRcFZXH0LOvFNHbvDv42BvCK+/+5BzlJlwSx1age+M67/1m
ezKjFmpJY++L1TQ4VJMfLzaibvjVlwoSswt/GkTSe/Tcjj4LfFLAzR/SCT8XMivmTK7+UXv+9GeA
As7g443XSEmRom9v9loIcRsBl0+3rdKlkEX85IlQTI998V1yfMsXHhcHhrRIwXGuBHoBRLTpPrF0
J0NsDPR2T2/j8CF7SvtiRXBD95pKStQM4EqUcqDPGpyVMaWtEhEbf3C5C4bDtgDHZGzOrhMVWmiN
XjBCAlh3RBeDwpPijmpFQ81mt52Mx0VMrw7QXOcnkC8cvp34iTToltN7ZfJI3s09HlTVA5yXDeqS
Yui9TbrnAhcb/FMr1uJEB0cxYBMAt6r6D4I7kHVLg1yy14cxEmp1AgPQMk9bbhXA227CAHHn9qCm
+65KjIZAbgpo9oa9jHXAnQZvfHzfooJdn5Fyt2YeLoKt/fDyI7nfsnrfC87YNyCquKlRUc5LRvbY
X2garRtHiz1jOopq08iT3tyDSnE+dK/W3kZGPwl1AJ4TLFfWbZhmcYFLjLrjM5YG15jbMemnMHEf
wr5VA9t4mDld8H02Manns2gwr0pU9MAv2CuHJYTKWrDBB6ri5Kk4mPUCvgWRF7lARlHOrVv64SkS
i9wpyvsrpeVF6fk3a9dnaJ53nXajuW2zALx+RJEPwub0ogxjijtmJpNjcxjw3mzEDaSp2hXKXq3C
Ob49+QNaMLIwR+IPwkJoPosDHT7NqIHs9GdzBf674anxUabbnzDb8AlrioynnYgJC1F2KBt9I14R
TFS/hFG7kA1B+Gof0Z1tD1ybF4O9sV6rAAM9hwGtXFqAP/d/WxH4kBsS5STRQwELtWBqptgIA8g3
rwLPQhgxk1HXZANBrqp3nqMKWSBYffnyC9ZoAWQ+zOFBkAv5dOTE9Tv9DEWPm1STzfyryuSpIzGV
DXdo2MXRtpOjrvi0y/a/hLqSgY8hMw336w1lOeQVSvEpz2c5q6pZQ9z674hidGrb9U4S0/RWXp1t
9gP2LHpycyAJvDLpOyw9cmfl9zAdEivFJAKxQ9hjm+nIQ1YOcEP3hlxU1JJtXUisBJ8s+eLTiKko
XIiFJ6IUiTpkb5NnZqOiCq1K3iix4W9pQok/1CltdFKgWVCS0o0+jAwZw00tw495YDTiJfQlrGYo
NCrnABwCPGUQ1KJamAbSuakfSPxt/9gJNy5rTQNKExcgHKIK8kq0bzKyvyMgNvKYRqD/Om5+D69d
Jjec+sUAp62YRGqVJLviXz/9eXDH9i8oh4xxf0Lh6i4RfVakvlLQ9gjPebfYiyxjF3F6BH3+BsZG
xbE91+iyb6ogiuUfXb0Vly/3kPTVUxSSh0NdeqpPCAQuuBzLoEVks2/F/BUDRqO4xl2Nc+9eleK6
mqWD07Uk/6R1gyHioI3VC1mkXDno+v+6rhGBzAIN8cwq0VG2fYrqge1g6Q2Oy1DaI+QKpjkPI2To
V4rd2KhpoZel6srCPGUU3LmmWi5uCm06bQ6su0dMtmUyVrh5/RE80Zo+balh349pin5QRl6T1cWC
rwjAPwgyn8rXEfpG+opoaYCp6ZN+ZWquqqn4KzVfv14ixlpek8NM3hoyeb4lW/ni5yX4dcsiRLja
PuiWwGrOT6BvHIL4R3NmZALTysScEXChgVB8Huzu0a/53WFKK7JHtU5OncNcNWTTYhba2rGjZbhL
/CFlDeb93mMr5mLz59zPa7nYx6q1vFPTkwfQRE28+7vHOeZyF8/QtvY8JhH7pfsogoJf14F2k8Du
BtCpcoWYFDFQLLo4ETdJvwAgimob/961J+LJ+8L3FJ04n7MlVBd7Ht2/O+oaceX270gFXZfuA08h
t2kCNaX+AnR+OzlH7sGiXtKq7K9ZElzx1RLe9FPyZMBxM9nLBJOd8MrdJQGpY5VU9G3rGV12EtPs
Q608EOQlMRWUxBm1JR624c/Io4U77zZe1gLTBDyHLKmOToYWTJWR1OpooLcFhGni2iJ1kMUtgdUa
eDvRWXs8YTydNesxnccP1EvP/VUbj4oxx+48ncDEFL9AWYGxTPfggeBDPiuj9j9XkwyIg0WoZJDh
lSWO/5/KX1kKU8bPAR7X34btoOdtYV1ltsqrpLcS6/E/9nA9wWk2WOwDDJpkrnr0kp6C3I5brBE/
6BCtdd5INVNVn2kJqlHJUqOHaZrbUlfjLPWDH5WUdyq0QORbrCNdP/ii8vyzNUeIqZj7LbSwURiD
bQgOA4r3PLwDeCuXIa0BV6LYjfiskBsctO17Ssf29JMtzzPiVFPZ6RwUM72kZYTVSbgpnt1lIV1k
CKr0losK+D4iDedd8nTziRosgapg7/koYVbnGrhxozWWsx/K1VIjyARkWrnZDoMAONxy6h1rDgWN
jn8nJzRlx4ACmX3qlJ7qmyPDKV64HwoKaZOuAhOqEEuWpHQYxpBoiYLOeuFr4zPh8pgoKTC2vtXU
3O9nytcdm+FLTGpTDRaTkxrkcgaEx7jVc2ja9KYIKr9EazTXtXjzmIqRQ7sfC0d0/+SF4r3Yi4Wd
dWjAZ/IKGVhyKMpeS3SJPGDGidVrxFr/uvLuWrPyd6lMnnDFZtGI2g6r8013lLRoB3srQ1NXtl5R
NyBuD9qY/WAzSRDNr3uN5v6xI1/JBgbajm+3DL0Q2Jcp12dxyRptpA/r7tIUK2iBpn/81aXA6b5P
kQ9oKQdH2u4nFre5c5xuHMeoKkV1URCE7kz/OjmftrHVI5CqvGX1p7+aczHVERExONx63xFQRI9A
GVfZYwrlizYCldsJ/Te7S70UnpAP0ND+M91eJ39n6Y1d5MNidlJxtbFikldw9rigM2uAyXhv0F62
fnkdpkQlGrZXcMau9kOAyu2hiSE/BstptbzIPqf9iyUEgsBSfgBhjSR57wH3i/5+8kmXr4evXpg7
kZTbc9ufu9NU008Q4yaztLF+nmaZWF9OMe/96XuclnEUkoWxLAk3zYekqe1D5GIcKbQH5xocn1yI
bwykmMB4b1CFoJ0HXC2gZz36YH4M6088JuKPdoVmo188Nks1P3Hu8FqnFZ2uGrdHhHt7gI0I50+S
v8NrbdMDI2xZGekmsz2rzeVGiHLp76WhScK/qlWzInP2A/eapRhlIRqdGgIvAJOWrxL0sVXxg0n6
F/0SD72yDMAHch1RrgOPiUPgFqxmNpPII7XfcL6kP4a07hac6dXm+RIS4/b2Dib+fPNwelAvo0sh
4UyQIpdILjpUkyBjEeNn/zNF2LGAAWA7y/p8Jili2f+g4oVteXusTa68MDDjhdnA0D5pUJ64JPZX
4tPWt+A0J5TZ9eYXyp51vlU7vynkTBVBnl5FTkTKP/c4e1p8mNwsp95qnIl4QY/neH5J5AyDTCiO
dmxd8LP9MMPIsWdg10XClt+C8ySzK9EA03KAc6BM0gZH5ne48cKCzt56OUUGDV0C2l65k+4hAipk
0Z8V7Vneb1G9p36/24/ot9sJZbcGUta/DI5YTWAwJM0/wPRbRtW21tXm82Llkyic9bIewd+o6Xfg
RumoUR5hvjGcvTstIMT8y+WeIhgrWKy4klIsICLEsD8Q4sw3f4fxijj//1WNFiKjYvtOQPbvbWgP
egrbxty97y0boahN+yFNCXuLQpFjijBlAeud+9wVBo4fX3gEE1girvo33g4+d/cseuMGM0QrW2dc
w/Gf5CPXxnvP52JfUPRpKoobBqatdWovGPK3P/wM8uoLsousKW3Ja/69MxHsJB/dZf9KTmWr40z3
5/MMHVngIuQmpboVRvQflSKxXr/hbTNt1rV8hwps6+yelJx3LyH5+F9o3kvLzmNl5I9WqvNUrA7R
aCoihwMKCG0EbT1UPcJwyAEeRzxOxG2/muMsjW47INLbikR+9tBJZPl1ESxo07HdmxfzSGshNGF1
xIck9DqdcT7rt50e7ZR1w30RUuGGxtPA9vq9oDmDm1jbDYgrSTGfpvdF7tP6ZPi079H9hNMpdH/Q
cBe7UMiDec/IoXwBY7a2nAuqp1MXE2rEDdvxQJ8+e8LCs2ut2IefEsEkr8OJM/kVL8rpYYLwMv7b
GPkg+bvZWr+5EUTHRTJ91VTsP9GnHBxYr2RZSIXu4h+b/t6Ncz11kJYUeKJm9TqGTg+pmkRqi0hp
Rhj84hZTA91R3hTRmBAinYem8eDM1ZW7c99TBPObVc3uGPJ49q/eMkIz6gbYVQAEbDStIuBQbVRp
a5/UgYKANARQ+776wVmCP9uxGtHCin/eN2GsfQ+BGxbRQlRR6U/sfwhAUvd2+WjoaYLp03/OUeDO
5XkSwHnOs/ND1IsA9X0envMIjSBUOr6LKAA8ky6fPZHpJC5XN0MfduOe/DHGPR6Rd0z6Y/VPT33N
bnymLEykaspYB1+K6IK2hw6zBl3zawhr8A6JIqDa3kVnU4oy3+UaofpW/ZHbR9PfMcsS3kKJ+OE2
UbFLzGKdLM6XvbkCuegkuupRNETDVODjDP7yMWljRbYwZ7AtnILm196cV9LNRSQYRgJbzGUZAWfN
cZT9f1kDGJqPze4te3ylx5r33Oglk8cfv3dGtuCmyT+UiCu6gmv3S3aw2M8FZ5Ra4gsTN5Z74dJJ
kZ7nJVwfO0322ZL2q6e6n1nVo2LzPmbQo7Zx3bx0fijbJn9lZ+wjtidAss4U3/J8WrgRbbQo5ZB3
XmxCoccwDuGCcUhiL+gKcET1m2J9LvByDTklEY4oldqcFw7J1RgR1FcTfdKvK8ncKWuiCGMThhzB
b9br62W3mAW+mMKsmwbj3bYb9WpZlHa45aaXTKI7Gq0goTHutXr6bA1OrXbMrPu5OMNhY6fpIW0q
7SERzklCVjCiTIyoPyXCqi8sDgpM5JIo2TwSyw0N9HSZNyWhC61TPuj8eChq2p+NeCFs33t57bYU
bR0ilO3Ru/WqVfhJiG4Tv5koTCuRsaq+DpqqDyP7HdDfODH4BxuMH06SvPvljz+toaHtg6rTA40J
uviI2DVUaJN526xJ0JyasQnQQras7CCUXVlbmT1Dx/JY4LO55aAncsaAJs4O829xFpMMPh45hvES
x0OwSxM6IPIHUGqi7HjK2xLUZbTdhvkQPtKsIlfmyWecRBpk6XhoE65rXZXa2WoOn+hO799s9HEz
kOp11waB6Bl2dBbsmfFwv4iGWcWrCRnovrd6UpqJweE5xLpFBezRrBJ9QilAWXtizOwu5XSIcKO4
Pa54s0WS1tbBTChvwYZr1SiO5GgzFlZSgfc53Yj7NcpBoPEyx3noJWuOkbjAcWPimpKNXVbACwKo
4/BzLfYnPnryT6KeELRa5qUvHbW2PwAf8ynX8uWNm5knpg6v7HnlYV9ByPx/2ArV7+BrldJn+J47
UrNnM+c4meaBUIBjf+wrlylAQEYYkSo7lxlU1znP5SvVY7JWjQynZ5KK9tML1zRDBpo9MPDcoKIS
Cz4eQjiL82jVSDo0hoHYF34GZ6BFhgTF4mB4bhoapFR7npt+1E+mz+pf6subUZC9X6WuB53jyUtF
i0p8RZNHyBojXYQPaLOWk4BFQwUUQjbFb8hxZsyK+yaXwKKic5JkiXk+noa1/o48PYJFyPrZRMgd
ui3PIKcDDyjDI/8bLzArYnMWnJlnSVGXQX32KC4DjecDo/GyaYd/pT8fO4MgC6CWDxXRuf/uMRiK
2H49tjoUo2kYjabTVuieiY0nxtDyUppaiF8UZpCa9G3ZLwmayrdlBI6pHd2hApBGcapxe9BcUFCv
AZ5Hh8iYdkxJKQBeSTbu2PFAiMjVKnlng5IaRdcA4nU5KHeUYUuVPzwOHgkvWoi3HqCzDV/Eh7bB
0qkbi4dmSu9qNlpGqX9zBEf4WdwYZf5+vEdePI7ybbUDqdChDeabwJu6R3/G3OtDIGwmSpoGchiF
fEcGrkBFOHkB0vEAP+b13jqtDeppruJInJT26IEur7KSVa2YMJl89KvlIIRVIC+84UXLEMD3q7to
U1Ugetp2yITPisFsFHXxrzmA63jkq2foVjedTLSgbqghIgj9BOzEoSYLsB8Gj01sLHCquefiPOa+
eLCK1wEZYau7vQhDm3yWYq93WsMGI5zqQyjwd69iiBTJJagotVZliilkkTWTt9+ooDbxXu3n7owq
L4owsribu7n3QlnEZoP+KKHZMe2Px+zpyo6nJOL9Amub0Rtf4ufONaw+FbBRR0fyRfqSvb4V5nRZ
uMrGBnINDz6m0QU3cvR8KL8ROX1lKA2EZzhbu6yXMsS/432yKVBS/HEscjJfILhLc5IF6FXc9PpP
Qi59X80y/d7M2MKXgptY2JPgrH2FubkrOz8s8k0Q3KDOtdu8PuKszYac5pK5y/RuVY28J4Cj7WZu
b/ketxnN5E/GD5YMeBwVXzIs7nspkWVOS/JxoebYktxkCA3XuaUA3jo1Co7Tcw6+taeqh5+0kVyV
RKwvUi7mckzveBjdZLPge61PpQRvUNWtR/h3Ae52AsyTx06eQ9qcDKTjnw44Dm/w0w3WITgMkvN/
E5Jw9JREWPPqOM0b01/N4nY9nw+C6uxZgXosigUhOTA51g9LQC0ppQx+iKVq8eaFcm92J1CUZxLX
jebHJraj/0L90tVQ5Go/aV88wqMRyx2m70BEBlVvf2rwANsKwWKUT7sOraMUzUPKxh5AMUI+1F1T
NtpeAvJjS7powTAPlRUYdYy43sAytTroBv58tK1r73BptMXWP48xuCaGvoOoVu8Fu+zt21xDQ+BX
bs4MZEMmp798uxcIEqznRNSm8TTFl1R+IG3xFPS9PRuP8TRk7IzN8q/OnVerJpfe72r1sDcvjr4F
9M3iEAXLz8YL1RfZx32Kxgfk+wd5Kv2XnxVwI9xUtTrQ+Bul/OANAtEZdiAtMw1HTzbLduICxMf4
9wV/2egx+vVMMIFlXT1HfC/ynK+6cJq8iOOz14xhEjsQJCYOoOmxhSj2v7YlxNxHGkdglk8MbKBf
tDMzJEVoiW9z/Od/Jh5w2BBRvgs8GEJsLERegocDtAaK9p3WQxlOYGiaGdMgNjSJlpVhb9Hz0Eln
wwGPezPReO3/l9m6h/vGBNE199CQQPhYhRZono+AGaaadqsmCL9X1G9mDoGC2aM/IrxSRT23X13O
+4rWuaMFVhxfoU7jtb2XngQiX5l8D7WCURO+4lXaiMiHV7iqbz/IQflgk9TGHnZzwAc+GrVj4lLY
0qg4Vz27UaIqHxmIdtQ6Ok4ump6AKyb5iGKOk6QBCQztbi9pbZY7FzEyarjmQKBSdQmEjytCrJML
ab82fORXsQaZed0h1BjrgcMeBITKwjrB4siXWxJ5G0r2FcRwX/dxiLQE2GAvmBE93eoSVzR4gEEl
2f85QiLmWS++OwCXRm8BOQC4MqvOdwfFiSjh2+sxD3UQcnzWjPrYR+kbajlX8F736X7DitkaxH5n
vnZTOuuOaRiWPUI/z6pN+FezM2T5L2RtC+uaP5jrgxPSuDPLbWs7cSmXX/jbQvd5a4JAx6bMNypK
LhR6MjKg7Rx6ekX9Q/aZ2DXdXxUPubLaBd2n8exgqvaGo7ofuzs1p6xQc1y5TjnrHvGtOi4fAgEr
l+T2fsU30NBxAAJzOc/BAgOi4Gc2S+mg1O3IAjuHdCbixj0ajH79xYgnPRhuq+8QXbhXm4noHDyf
oc4IsCE65U892TmIEwugmxIQFe3pVFTWz+/kjLUn3qD7s/PMIEZkZnpE2tBEyyIbXpXzJHXI1cec
MaU9GzlVP3/pXCieLsQ4aXls5501Peo5mEfGjwIaCV7te4NmM9z6qDAYrpyG0ED0NmanW85eGHvW
f+DKLp9o90864meHDWjwJnsuXB5wp6+uyNn4xLzG5qwN59X4wCwXhuYmdcSeMzCUMKTMyRMYAkcH
bcbbHayp5p33ZbOjw0Z+2km9DN/t/s9l0Q/7XM4TSBfEvK4pd7Xszqu4fPaopO0XKRXVaGjmZ2JE
j/oYCJmEfgbwLrLx869E1i0gB7Ovwv2N39gc0LQQLfB1tMHoidglF9NV4MlAi+Bwn6UexDaUwKKi
AfeewmevlYUJA9KiEmZa+w0i3G3NFRT8/8G43f94GbDiey0Nd83ROPon78xbzjhcJgHKts4P6sGJ
j9zvqH4Ljy6CR4Do/9HjNaxj43SVV1MVhB/T5imG0ju+XnpYlSWJMzNh4TVT72Q0R6AQXZSoxRjc
YqrYMSK2h2EO2rE+6VX9A3g2/t4wdLZCOGVRdpBs73+dviIcAtb/8zDOcCLInjvXqIdY/TTbT7XJ
LEwpsQNZXNwq0xLljHvxlgaHaajhINRLbvOWGvzjEwPEU1MZcPLaH9pL4nahmtL2KHZgzP/OvoJP
fmEx8jdLV0cfYEHLWZ7poR7u5HD3JKY2VFDDswmJ9EVAfimRYhj2FscaHgKnNikEZLDB6LOSxF8g
SUAJtPr3FfROyL8XWmo5SxPj9G9wsuTwc9nRaSCMKgMZTvqzkLicKyEHCsvDP4x43sgvVXrRHcF/
ZHxh4z0O1VlBF7pqZspykmv6e3sejWVpov2GbbBK2mlBNmujkOPCC3vvLdz8j+tC5OE2rdujNCxX
RPJh1VHsLI9TEzBp79HKO75SBi5YzFXQ4vu20WYa1fx+bWILfUYwNb47JPXC7AbMKmfomZ+d9cVO
3sBXde74yvNkF/0lVKzALc/UosCXxHg758xmu62P8wftt+nQ237Az8VX9J3kbd4C9WYbZNPMoBkE
DtQ1Bkm4RbJCuYmPE9JOMblA7O8o+lruhrrnjd31QCdfjusCBH0Q4Zcd2hOacvyaOrGnNnMs+kVz
uKKOZ++JwJbC0pEZdh/dcJkM3C2lDi7GQMXk8lngW8F/SD5iSliUYh4qHzNAfHegIDs2ZwjwDlV2
BTuL/SP3hps1zpetN5Ebr4ghufHT6Xt60VQbIqaX/CCKxCWHbUvzMlBNCzodwYQct1XoOEb6/uGJ
iwb7hQ++HHnIbTbwGQu+fNi7MUIrLTFW44+HIigxD+cDQ5BIW0Ppj1GSrp2CloF3m0KUU1Jphe9E
1iP09kMD1Sv7aYl59s0S4+IIn/8ORmCn3t1SNCGtXxcYBByFK/AL9/lHz/6hNoVBpKlTx6Clwq+1
M0nyg4P0m4rnbzmSs6D5gIttix6dE7QyZzk+jXQm+R72j+LWjQh9+kB36q8CBGSPgjgv0skX9lUm
ly/pil2r/O7EUyG5o/RHJ6eVf2+h6qR5cq3YYwnmzQtPHUC7BUsLEu/TE+ZUBBubQ3Icf6y7+z9w
8HXWs28d0MinjBaQ6GKLsdFhLUvSNoWxv1k2z0bW5wFZotlmtWZwpF8jLXhG2CYO1xlvahNb3VU3
aiAfpJJbvCQycO3CO6o3+ml8ulsYnoodRc3EeA+sp5o3k5ppfax0wZ//wMx5RAceA8IDyzcx/ITV
UDOzHjkUe70I8JvjkNhUsIlp78fF2OS5iuxBfBzdPWWORMwL0Y/ao2v7vwBPcW4MDeXWguAWSRTR
DXV7tlrkzm3ErZ4LLAvOopg28OaMRTUMHxyJQjuuRZTPoc6W4AqbIXqfq6x5fInONMNBOQdbgiJ1
t5dQp81szhSJlcSKj7l4iu7FaIV6NuQgA++THFyNjFlXTfPBazCL7P/gQfyt+cZJ5K51LixL45kc
xRnPn4Ka8NOA/S7GQq09q3IBF+BERmy9M7/qYqRczWXuWB7AKvb59OoSWsnAQkIa2BIYZr8dlYPe
U0LkL6rlr0PjNd/hbL1N+rDYaBmTYooUaWR8PmR1ibS0uyy+R0Myv9Vz91RSp1Rw3TP1ZTDG+ScG
OeJA2VU7hBKNGHayzMVh4nP+K1xDJXnGPETuCSSYlGA8Mkc7+hZpGyfFD1VMTfC9h47isSUScnsy
YHG5IKThiOT45MTLNO8+KLcLmXTSujCmE1P2F5G0Q6iAfQW/YOUQK0za3hSqsn1llPMFZQwE0fWf
e3Yqg1qC7ib6lCGYNcsIPWy9H61xQWy+xVEO5Sk3h38oF7y1pqs2otJnG3H46aDstHZTmLPwazTQ
CqyIhLiOAfrw4kVW5C8biwKXTr5ccOCqVfT7FMSovIJCMkLLxnG6rpZ8K+yJzsB7Gm4H/YOSDm2C
LudG6teK4fgS/ey9bJjg++NanS/WDRKAyjotIFhhWPqDQnkYELPIjbN4Da6FPPu+7eJOf6CyI8JB
AIGETy49lSpSTYtJkiA9k5jMJALgt4qGwhS+jMGnshcaXFfJdUPs6bydV3PNJSMDy4LxqLy3+QaE
zZDFiG7iMTpYltVd0wO+4bA0KNnNgT8nh71owSUZOUctQvicA12R29qr9xpreyd9q+Q8TmituDc6
WZh9NauEClL1z93cdklqhbZNQ6bi65MUrBUZrgwGIRhULO2t4nOqpOS7GOt4E/deJVUg5Y67AelY
lbUtHKn39ZnVm9Hx1pttrKwlaVAPHHO+EPTOxfvUWLMr1you46O7H2SUfaus8vestVH6ngOxmRjc
FfB9ErYQT0a+jl+OvyFocfpN3grDQ3/S/GMyOH11x31O+Ibj/q/uo6yAsRuOiRekKBdnR2CfwXU3
k1Tz8O4HCu1KT4sq5DG5lpkEq6JHDAIcRLXyL+wS64//w9n+iZsGhqcY7g5FLTRFbC/2fvqL2XSm
gAtCw+MGs81oaCznOvT7pZZNMQ0RGLJSz7xWa1B6rF/oOG88O9qF9GSXrOCf+rZ5Iu3Wxx4FXGdr
aDI9MccaIXGbLDYVEyqwCU6X4YwWSw4piUUOIh5ZwiICaqSF4jQJt4azixEYDYPfL20IbxnLM6Vp
+JtSfYPRZssCaJZmd6itFyqTbyahx848pPLP+SZUZoL7F/s7ULYFN6VuSDid5vq8wwrn9MaJkYHc
MiGU/Q/LqiJtm9VGFGt65ki6f7r8fd5h8N9neXNNNPzgcuQWSiCmfGNSk5w4JMlZQyJa4BjoDgus
+ia4+Hrz10DWOJvQzlBBMhJkkYT4IO62fMS2ji46lexc9IYw8j1V/Vk7VDegtv36biFn+3XycRhn
mC35Np/Vf0z9uWbGiRBGHTpK7fmREYDTU5RJxpD5vb8wzbBlrHpkJJqRMh3I/hLv/42tSlvHMPNO
ma/7+gbBs8KaCj6uX8rBPh4jFvXlgRb9tLoqaf26oU+yB8MzFnOH7r+SDhoCSs0fFiF/GrBGIpmi
tckKIC07j3Whe/aANyu4qOldNdtFrdiQH2uLS/OBz5LnAltyTQ3kwF7MV6vL4V9oDeroDRDYjf9n
CHCI99jEiXvKsAcU+j+9RPDFVyBWuJ5OMAe1As4s+OI1s5cAKd0pOAzUH09sAjsUQKTQ9XWebqmn
O9RbWbXlM89EOBnbXFn9FHItsoEGkmHQ4KSPp2UOOztUmE0fNqLtvPChD0ObEqja6TLXR6Ut6VuI
6eRkD6sSPkaI1xpQOWUDvce3WputSffo4cmnXxHN4dU4BcIWnuT8bCmX9gVHDJhFgoqil37cwoV4
opKLeXlEkbT3uRy46xW4LPWIa3bYl+cHTSsKkeXLv/zpuX76ydPJcZXbZ66JY0FRve83uRVAR+5r
UzhQlVAyhixGFDyDa5fpQKJJDQy4f568nCaumrwHmGW6iFDVCXeyBQWeGA5JIj83feBQSMwewyzT
nBdsEHxG36b0cwBQbvJBVtAZQfe1jGv+qR12q55REddbF2BWE9HCCe4dsMyQ40rUqgcWcui8rOny
khhgwT0XGZAUwSQPCxUw8u2DABC14aBEPoKn2H2sAX1sCC88PjWKhpYtdFt8hgJtOpdAzObktIJ1
j4qwxGEQWceSBGooc5HM42nq9nSzvcoIwHHb9DR0XyhrL6FetSGcysx6eaIjTerkKbOubaT7LRol
kyMyOWp7QrE74diIjS4769/IKNvN4gh4Es9Ta0cUVWzDtuVbpITptqgYLr0nyrGSkhZwRekz6If6
zvGlvhU5UTKiOKmg/cRo4xE0Pz8p3BAz4RTpXQvw3zLx9FDuAKc3HogIEkpgdAiaBqZN/PB5kswm
EP/MkfhrmZtN7q1SYpFOD81OYXhyavw8j4hh2PzyAGkyG0yTyPn2kAlDg0bvH6liJ8bJXjkRMh7i
CR8zkbC/kkHiM3eBZJoMdJu22IqLhl5x1XwSt7FttSZ/kCXuO3RGBTA7P7qR5w5Z89kMc7rV2sbO
D1BMqUSpV9eAHQmLoESGXev0glCWKeLDZsLYneXiKbhQ7dFgJ3N9Jvl/9c3U3dL24LD5Okh2pZaM
a4sny0G9T4lzbxp5NGmaVIAlEyiZbySSx45Avudbzlmojk+CgV2+gyHnfqhLaFQWm3rJlmyzsWuz
gG2Uu+xMmeI9iSONS0kHRrzExInLiaf6ze/lpRduH//TJOQtvI+tYXbuWhaFcOy2aGbuPLrtI+IJ
2Tr6mCxzfukckJ5unUDzePZQ3/ljKRWYxmi0DasNdmFI7aAyRcVF7sfz5mANTF1jq/H+/lsdAskR
6Lha5CMgQGq1sydfy8O78Z4cMSd4V9jZFwN50BaZ7BYhX7nhLCdrTg0cQpHv9D/zGFjt600py8pM
AWt4zJ1OybVjF+yEDPNzEXDVsEb02u22T1/0/gLaOAKRmUQEb8P7r66XyIMQ62xugyGesyR47Gvb
uaELTbAJpcRWQHObWpr/zT5AqhlbQWW4UpNAfaRr7OcERV9LkrvfuvURtAzSHZW85MQRMh+5vw/u
S97D2XcOYbDENHj/bSXwu5hEU7kekqYXsrRsGg357R5dI0VcW2ygXuWiv8gwn5FogTLWx5JOCVlg
A1sIB3g8ja6osrY8O1PVWvtw4RnUq6RjcTvvWgvkgYTDWV+HlFFIEWg+C9bl1IzkWt85z1zCWN6Y
Ni7TIbpEi1KWHILRTixOlNGHK+blyp4GZGUrSQyABCHBedLDjrnTP5Pb98buGprWRfiHPTQj4CvV
oDn4jNQo1l7a56nW6hQeYsdMXXy6IBB7jNhXdJC6clLRAZf3ArCCvscpyWtFYq/5emB45b/L4qr5
I2tTm48kj9w+8MCllORI3pYXWpCz5Chj72lZCwt1DE2EoFmVgQnO1CeG9TXnhLHDbCEhTUHIRsCI
+Zt3LNtxnI8yxFGf8WicKVT1JOKLr6H1YzBnJ/3onshY/Q/GNLfDB3n8uSSluTDTvPDfkSKysBfX
hJuFHfdRe1yGfbJZGKmdKppgfK+bVJNUEwcuScycgMVunfhPD5l5xXj3ljMOxMVshhdv/Xn0FZzF
+RTnt42/8fJfP2Ji3QxesPYE3MdI5cfD89otiK8o94HPTzqXwP9BVoAldHprtMVLyAefcH1GUhJm
0e5z4DSlTBZehH4DlWWpIqb6JBJA7UCmPhtVgmVtT4hB5j9HqZt4XczOKM9O/yYV71nNXNEcnj8f
VVef3yZcWzRHCer8IlAexgwLloyOxvDVyh/z4eQONKFHMvCtEYlY2I0NgyoaIy1GrhEFWx5nSVmA
xf6GJbYKvNsORZ6ecDmFKCViYD1mCuUApFMP6K9HybYTboaWqePcydxADjTra2w7s2eVShAA16aA
FsFVvC3B9r8+7l1zPwuO+hiKY3wf41OAKEjRb7wOBmvyu+ccUtRnwXIHgYnEcTBnws5/8XCIWrmj
Ikc3yeKVSwCVymaL5SMO1fSVEclU/nTZ3KxOCp+GrsJ1T0pQLeGP7sKyqjNL7c4mgFbcFo4C4MbG
0Nnd0qJMMbV3jR1x7dWlyuvdirPoaF8MfnkGqjTdoa0fjHXEAr6uhKMXDHOK1pQG/accAyE27+oE
UwJCQuTxcljxwKVL3UsmJGf2EogOPjFHHygW1IjossHU7wuRrJRRmo/k70Q8TATTsDF6TRNvBW/x
PuJJqfhp9L54bjs46XyFXxox4er3VUHpvSeVv1yiX0HDmB3XeOOt3apxZe3kpqEiEdXreq+/27R4
xCBCu2WwRnjl9wVwvPKOkCXd/PnN7/D8/TXFbis+chp7w6GQHR+6oUCjcnptd9r2m6S9lyQjH7Na
sZ/L+x/XErRDq0AdBHsYMUkxyXi4ExCR17TgXZFR+3JzQVJ1ZdCuOBZYBQBLS/dQ1CkKDjEqNnrf
bYGOQqz/Xmt5ObxTuQGc8McwQTMi2ZrjyKCTK72ECZ4rbE6Bsu7TcYDR4PVMN9mstlFV7OZNRVL2
6S8kZXoWbZAMjDga8Ck5AFu+qRhsbCO1Iod4DGy4zzAo/17nHiZk2RbahEijtg7nXrk50VDjG1On
wnK91inyrtnDw+PBp+2HTockw2dJ3lZP3uqj3ImKnW+ccoK95TMnofVbuFtCS4iWSRcHK7uaCXEd
JjFpr/t4Vl++eFak3Geery/3oUOuBTPN+7TS6aCgEUPszfZNxBkqJhNamIr9cl9nTI+5WIEGISIN
JBMLJU1xbumfdYg6F3s55do9nSoQS+9t+RXTSyMLMi3d2Z0g2SEYr45Jx8tzQHh686BwWfErDMvT
TfIwabz+6dLxyRD1vVNvqIlB9pvP8fX90HX+ImTwPjsVdRasIReGX61P4UELFERvt5LCFbeikYT9
Ej+kaVwVL2j4sdlVvAXNhpXx9CW2IhXopYD2pBH1JR4p1dnkQdjtZuzGyGgfWlmBlxs/9QkM1mLd
Qd692X0y7MKUtJnrxMhZezDEb7aLfk0nCyFx4lR/vDfwiAW9poJSKB4qNJmKhX6rM0+32KxtCXK3
RwYkHo2XBM3GBMVqBNR49wq8zlOXg6R+Xnq6dJW+oGBEDQ3tfey451+KKEW4DRQcQZ6KBTXhuYbn
5XqEJKn3+sTZqLu3ELeaKrknxvq2ROHEMOXmOiJoaek/cXiMPWyFU0ZRgLzMz7P1x2o0/5I8eKT/
EMjrNfKfu54QnT5b99ap/cN4RlLChOxv2bfKECHZYpqMYV6VXja639duoFWJkRCUKLHpkFECAB37
zM+VHXIpZmA7rBMsSLs8dbM+ibWzyEvX5oDbSCskOon5ROf5yo6JcKu+OAwoajw5XVMoMNKaUH7q
3hM1U2LNY7d3PTXxQJ1FIqS364eK3UMr5hlAKvdAPqteDfQsJs4a0K3FFilyGaHtd9TniwuMTpEj
CpjY9Ss0jiY3v1VTW4HwjTE2scxUB3D7n02wH1np5KBmWwYxg+9ZhUzkZiv7KLRG+Glwf2hPNsJY
ka6FX5HVGdl8SrA5u5xzzsYUCx75Wpn9nOs92YRPuZsQmoNjhQ25etsxb5Qnns52H02fSIdGtnvF
lfNEvTn1yYhdSVyqtY+7jSHoZtg4VGN+2BKQ6bDm2nTZK7omJ3hEUgYSf39nIt1Duq5TLTgCMNpO
AsFluSaDt8FhX/LPHqJqZ9MpDzEoZujFdCLTprq+SmYYcoQJqQuqDgbXhFNh7gBvjaxk9EtjEfmH
bc17cg5N82D8wj7Y/jztiAdagU45/FW7SmP6Ic2sNa0rnaHs2oIwZ4MF01pg/1tJA/j2SOMcYsq4
qFPpx4cXLXvTDloKDhCk/2wJQ0++PE4md4zF+0o5vhX+0vt9XSoYiAs27evGnN+u/u8xfYiCu1Bt
x+++rimE7GqvoZi7mTm5Ss+d13mtn/zrbr+0SPn15HKi1l5rwALlTXbAcy2NpYRzDgLNsUeMnI8R
lMm4TMaVSSJXvrbVQCBBo8BMFM3Ivp/0vnnyGTDWaDglSi/WIRbu4mJ2c6yBw4QFo2q0GbMNk4kq
dZV9p/XwNEZfjrq1A70mIS4y1xgbesjHCEdZ2XPYnG+cKM6ANFSQDbh95G8qzdcuNKVLUS0yNoPh
b3CLqJedsHNfgVLM91MBQfraeW3wdd1DRIV3sfyp4t5S4hH/c+VacQAOAY0KVDK2C8yOQRdKSlTW
qaD3LouDjDa+VUpoD+D0HrjHsqfSINryzvA1+8XzoE/DeYlzTHM/hos2eG95f4MBo17dTrtx7JYb
t72LOGyb1SybxXla6M0rR3urRh3YnCCDQtxVueQYzVw3b2KDM4ajDJ0ymzsw+ZZ221+FWZ0P2UM0
jHXKLE12673P0V/c4tGbDV4afCpOiW1mXXtPwln7WOYJap+/KJA2bt+TUguEW8OOKB80T9kdJF2z
AcmQnmASOHi5pw7+ZOtbfakW0yF4IxigP6FpmJVojm4EUpWBXSzpvljDG1ns0PeriIfbx/o10ys5
fsUaZaS9ZgJBIhV0DliF4uLXrVG5/MjMPEXDqBkXbjYErofHEJG3O/8ry/V7FKQWPMY5V5gzmfb5
xnP3Lo8/5FgSOo+B8HGitvxixm7r4a27AUhXKb7chai1JKs8VCVUpcm+zVGHDAqYIde4h51t7Pf+
INhcUYKK1NpEzyVa38pmU0JHMqAFBeGs7jGplJUo0cjBspi6WW134T69D58gcHlx5mLKYxNRf9eM
kDfvvLm+j4pMAAuUV1e2tJEesVDHKD3g5wSgoo2XC8A4GHUB/TEaXsxPjI6infzuCxQAMBTNNB1C
pdsxC4ioCRv/50q/mR/gd7+ByIA/GxrSMRo4Wp2vfcNxMYl15kMFBkorvjCfCLULf72UGP4RRpmm
NpXSVUuv02GVC/6FL7B2Jes76mieqlBZRJXmA4YXz05VwhWJ6QpOEe+GQT+SEu3kuL+NJLDgR7Db
zPOjusJEugGf1QRNgB+r09oU0S1KFFoGHL5kCtmUnlKkVlrgWJxk+Kl8LofuBiKzch0PpIjatCk5
lf9jCUlNp73nXMIr0cwD02TCCIbTlEO/7kP+B9laapo3/98j31SSXZ+kvOYY0fjEk1SCtDIC0Dxe
nX+rni2BtSPh2wji+eQFDnu6K2jZz+HTxwRqHJc8+rSVs18CnMBGxLYZEMn2IeUS8FIxqz+HLppi
SPt3HWteczPr4aFCbRojoJhYNsK+ALuF5DQuhyP1wS5mh1uoZ821/LpzgkPFrknhvOJSyTbz8JJQ
GMEDVe97TWV/2xClnCweErF2Aiy808kbJXewxlAopX7BEqvRrw1LKJmti406IWgvXTKxh6bRNFnV
ZBi9hqdVHudQGNj/O6xFqWnb0GnGA5JomiZ/FcEhUaboVvKqlTbKNANOgP9Ub+E9SzsaMmU0ZBoE
xuW+VinjHR2DlxjwhHyZEXFHD5pl4H4IWWD3xy0TSVTLLIdYV6amT+CnFGN0gWAc2cmuJtutN6OK
mAwSZ9MxZt06e/uZR1Fve6Yv27A+P7lWGzBnkkzMbQAD6Cq9JmLsZh6tGSYI9idjUTUC/sbu/RBh
iLjD+PIR/qq1iATlkLFcxOdSr4cySgKHZ6Gg5tjuuUBtvho6ECM3t4LO4dze5qwBO5tATqnRR6m2
7aon+a4fbL9LxpfIJFJCeYMK1L3nIBZ8l/i6hGGAlv4CsZ8Yv3L0hl/TIaSb/7u9OsE+4wlFyI0K
xwOLArFx6IYduxZqKVwxQ+w6J2Nq3IqnAtcS0JiR63EyIchVvVkgA7TVQoD3Tf+iFjjwSwjtLfti
dwMMjOtJSGAnu+Ae10NAYiKStYXN4kvXNhmB1yeNtYSdgsjN0ckaoGSmArSJGVb5eXcaXS/mMP2v
aGov979PPuPj7UdawnZl6r80Muri2O6Fd1DpOESlGYN4JKbGs6HcUZn/6bBoxTNVNaz0vGH5Rb4Z
cDaddvNV7JbAnUw4E6A7kk5ZP0DArihqVhdx7KX/esI6rpBveh/fdttStbIWTzV7OI5TO6Tjon0X
/RORQtLxvWZPv3LDGALK/R+OaEzgbIhUqp6lCpr2S2iqSrHSXZBTFRypXp9Y955To0+9Fesb4Bil
hQ1E65gG50uMAh4a4laH98xlz7wzIZGo9xhiT0l5quUdhQAjoxrNUEV6mx7qnpjocid7W3l2y2a8
2bz9nEVucZS/EIIdQ7FjXauWGG2hKZXZf7lDyoenO8dsrzuefE8oB1qIRfrATOvENdLYFd0AI1Dx
Uw155CVIqWdEEZ2qusDXFkIq20yESw5iyGQ2CsvIKuAWUUEnBfsMi7M50/wLh/0Z5DKTxYrgqrg1
0wzcX0Afcv76ZyRl5zL07kD+1kj0rjw5BPwNLzom5lJG3WadPWH2Fr5aZ4rtotT0jXi36cTWCyOr
8I8haV7EOTuIcqC7Y0ILXTNXU4TISOSj3savW0SMPkLTRoTOf7JRbnE2Ef731sRmYTrEkmgMrSnu
ir2sdkyyG1Nx+Ir3PMMXoywiATz59os3D3XZolxCjHaMZnYbRL5sh3Y2hWnxa3MVO1qYwPwNxYyH
5fpq2yp89Fzr8A/8DiL8BXbFT+/BlvL+dgg5qst3ArJAp9pCJ2co6A/99RjkVkfxcZlIEPnegLrr
xbRxLTZEizywLNurY8w/5deCt/oE0uxpbQwP0GB3Zi2CSPgIBdhTrTB1pX5PwrPsKRaGS9RhZCri
5uCODKjThEgDmQi6Q0EIYnTgTLJ9gJxDiUw5HBWDZUSkUKJivOMI3X3ou6DVfl3CVwSssgFGxCN2
gaYOvyhMoZlOHktdZ24g46lRmqpH2jsrJZaB5PtY2xwi2MBO0fYW+UE6XvuWQoMDfsY5I31FtQW1
4k/ZSrUlKuonpqbzmJ1sp5s3PXxAE2Y9Rt2FpEAX2LKb+xSDJiRCk0SMuA0JR1/JHRDZZVHyBbbF
GK5Z2l8vi+zbCu996uqQWmPDw8H/2UEln/Y/f7t4GNKRf33lwS+tsQzOJdHrMteTPO/iALCurrf3
TKCQ3zObPH/h4u8WKqYrnACoLYdw5BvezW3PdPdA1CbK/vIQe6aWTa1dbKnkr/2YiKEaWcl0P7yY
QoRQZt773tPFPwVsScWWbwrI96ONdtIc+xEZk8muk82gmEpMNkWk/X2IEYJVEt59cBWt+qhb3fBe
fx272tY7JZ3IMdnPs6zwA3ILOx0LT+IKKiiSbeFhJ8rDZTTFIdZqTxRB1kxonfLV9kIKTrV1Jwoj
t/Hqlt75fUqOpsfbQV63+vp20rE0/7tIyaXRPT8ZdbT9LrmleUntVv2VLLo2aBjC4s3zz4x8Kt4s
cYSEI0o/zBm1BYTQHN9IZevznspKggjpCdUXxngD6ks0E8CD8cHWHQXudogsLIL1X/TblaUye4Os
WD4nXfnSrhK5EzhQ+bmXflzdYi2X/utYZwHElwMP+4jvicJmLa1nSFhoVi7Pd4ug1rSGMHireIsX
OudmIczHvjYn86vPmv6WSef8Ah7UVRdMhwD2UlLEF1RMvFOV4y7Emr27li4Czjm0U0uwRYXJ8nMA
Cg5lKeFIv5U6q/GcGN5MG7CHwT9CUQnZBlOp8IHTnPOaihNY8RWhi2NjwABpzzFGV0pAV2r+Q4/E
ro6zrl2fBRPnp4V8OrIRyaRMOtXCP4rKtyE3gO+Ht8thlaZG55qn6IfjAHIEaSnSsvTdsY2arLjS
VgBzqRSL+FI6nUMnqD67VSExMPHUkQF2o61cdGPtnEUBYsMfvjzsMzkbDlPdMeQFGsJ3iN9dtIoC
jiGRE9zSFBS686SHWJEi0ka1s87H+h+uFHTkKxWmeQdIXrHMVYhYO0Um1EmTZ+w+puPDqxm9/vxv
VYRaTwb7JUYth0mLUOqVnGLmV+KciFGcnmoRpln0YgqZ1XD9rY2ZfgiGkVZDwelwUin8BceNXf1J
Gn2qcxPUf2qeMOK9iFVSUKbryoIg5csxf8KtN5e++3DTegKEnFFqqrYwzt8mlrJz+byAf2Rsvo0X
4cZrJ8YszZU0QD4D+Edi1m2HpxVD2025LH/LhpdM2CRSfgPhonj1RctmEdJSAZ+YIvphvIYzeuuF
iNbMmWM3znjJRPSxRaFZuVioIqnqlfVTkNZqHvdy+6H0fTP1fXQne2+k8uEyixQkon0c1wYaScNi
fyWrz5XYqDLmaG5Y0Dcg6zKgvv6griudWZ9NH+WtudC/XMn37sgcKBQ6HGNJq5lP5YNbl8X7vdmX
3ySvtg2xgHO3P2Zwv5cl/d/V0VM5Ci9nEhqBFl2EKwc4ufzprsQVzOCZQzO9zcnXv+3Gfc9h+zzA
kRGjjxN8TjAoCAucxu2+nkGcKDFjsquxdzmrdeVasxNIE8JEbLJEKBoE3TPBX408N3H2CIICVdoT
c+fn5isBL0xH9GfNmk7fRvFSrTLienaVy8wYig5Zs822tsyhZQzJtd6CT1+f75WrGxHZYsZfYdND
WEan4gLHYRTJ8zK/ceFYqQUQ55aUgsNhDgs/h3nKdKN1HVtiG2jWDE3AWAPAvrf9C1gAGaRHqGCc
bKcO2+stBQdj7tawLkaDdMPkpSSnOiTi8bCQVW9HWMa4kt6M0ui2aZzxL5OpDWbZL52WYhC9/DRI
bQtFfknaaFoK3tMXwvQdbPY1lPBEIc1/oTbuah0E1dvWD/ZH5v3geA+O++3s5pKqZOJUtkzwJg4N
tkl5fGitC6LbkgplN4PdWFzLUy/NKDF7J27zKtJv+DCJDP9vXStzQKS5Nk6lUeEVJkblsphIQzp3
NKrUfCt9BNEoM5LXalHY1CYD6c+/YKENJrMMK2W5HzIMMN0s41CbepAT2menjCQVQhl7rbAIAAGc
Sqlp5yxJokZmoA+dJZ28t3ElUNt6rvFlECyQUrQqz0Adc+XeUuc4ej0s/aFa8zdXYRqxFrdxEAnk
NjwUIijckHct/2pk9zudfo2OfNEA9rPL/zQGJp5poUI5MODsvagkXlhFC/gj5R/7BnMGlCSrfXiG
yV6npwr5euLLHIDHWmGml7oFALHxPzrznJ4IOpNaFTjqgL3VcUMlHsTiQb6eHlQwxHMM5NcIJgwT
p3J6JiX5X15haqRJyEMTlNon8kffrXDr8lHpuyl9yaieUo94xEN1IizoRaypf5y22qccmXAhTlyp
7+TBRYh6Tj2KDg3tB9j9BU8EWi4yxt3u8cBetCHNWen483KgYz1ngPvmI1ETrTdfIh3X5XZcNd7p
yUlAjYXym92ckhyCsyZX3E+9qZBw9yL9AJ5wOIn/gmMFj8M9j21nc8zZerpWgSYBPWAgmSwyZxn9
sebMf7D2vW0H6XJggaFPnS1OD+UmcqijrF7pM5M0QfxrOvNf8xm4hGfZZBLn5RQzlKuTjvtZN1qJ
vsFOJnUcZ0nexZyA/LpQ3t3sqHZuwKkRkP8VaxpfUjajqeszfsERqv+oD02rFt/bYcAnmC0WY72t
FZqL4TAqpC6BPkLQC/CmpnRbCP7LlFYkdw6ZTI6dawXjD6lIjUYPAJXPopRs2v0GW4Xf2w89rd31
OkpATPpRRDFyQlh6YPyTofBZ1RCz8R6RrF1l5yVk3E+9ouE8zaIQUGEG/cRhNaUg3hArhc9JDXSt
+Wk1QPF2FHu3D/qhJaQHmfsOWEct0vvvbtm3Km102YCZa3kmyBoVQDRbbBtthJFHW+OS0Z4I5zUY
7QPQ9S9FvHG1PelR8GkKyimMsS1DSJkXHJCqBJQF2Sel33vHw77G9LYnL0aWC1Kg8UrXTdTz/zpR
aWA1YSEYwS7jMWbEGgNiK+i4yU/avlyS/kXC4S3aPgER5I6rCmshEwAeulrX195nQiTnMPdrYAo2
dtF510chnFld9tkd+b3t1iWXClNCYSvn8uSSL5dkOgY491H7x92wp6VuqQck3Vt3aXBdRCrinxK6
r6cOsV1LXGkdBDLxxBpeim8LEu59GeOnw2015QZSVgUwMufu+oAVRZdEcUwncvCQ419bj/0cRtXM
jsuf/kLozArTl3cOBfafo8VCxGseouj65AgooT0x1GBgjOMuZuHb7SRNWkCopLE5x4aAw1y4AeYE
XPIA9lZgcLSsarzX0oJQOp/a7tAh140u66DqE4D+TPUhKBVwPIWU25eOUqDyVZQph0+XVBo6xcgA
+LX1sk45vy5musJ/kxxnv7uYZZ11uOGN4+YexImiS6ylIZWSepdmac3gV9YXHnzhyIDX2rkpi4WX
HPWVUCEQr8lW7qLuLKek4e1ZhEmGqR4NxPJZ65q43e88quK3TukCQ+Cozol8Xf+XDTnpUgC4UZg5
KfS3a3KxpOGpJY9wmr/5GtmN3i6A2X7NjVm0L7cMQ6EB61QGmm7cwlBqRgU8BlXcSiV1cDve4xx+
QgidRcj5CRi+RT7+uIFF/XGUtPzitwEKlWq3Oh3fqClPDNHqDIdnOe/Q//U4bFJVcnpxeHyaXYAc
HMqiaXkZxae3KqbCipe/TkyH67UHAFDztCpkwq6GIwtrHbhGAdhUvczbHor+UQa6KXt48WYz1JiB
e7j4/4wY2cg8hXAgZntNRnQfeSOF5ZWXOAB3xh37AbU5lTfEkfvlbEbndt+tAjNxtO+OwsfQ87Sr
5ir36nnH0P+8GiFO9WtLSsqhqsyjPuvhxJ68cKypzbQKtFuTW/Mm51xDW+KFLuvNob8hvyMo6OOy
l7WRbHGZCw6IlGiZzmLNXI2qk9vPBortcsi0SbmieLqk30OtEjZOyKv0/US9+GXFASxH9H7U5veZ
zFtlC5wLSQ84wWRaKTOZ6ClEyl/Q9QmYJVMCelrbQsFcsmNNFbXQJN8zF6+4jcGOlIScik5MXi2L
uEOj1cJIliWY657jcR3MGCmDf/eqMi8pZxCDriStflG+byrmQKTHIGr437F6Ug1jNnIKI6jUU7Kj
dulfB63hI+bFye46dofUBcLv8PPjd8mYJuRVvYWphV+RYWNNKDfk9xaGokG9/Q3UJfGGc70oY9x/
ijSy4fAJ2pvCH1BXPtkFebHcATzvB71bWP/AzLz3LUTycQjUk33RjJw6FYJZ6UViXNAEeNPTZlcW
4nzBex3KiepNUrrMnDRPRnZmZNhXYgrhR9KQOBWJ7q/oEOonsO8kNporZbQqdAJEoWm54X7fQ4I+
z/7QAN4fgRP7l5EZNarARgDgx9kx9XTdupJfp7xmNsGmjpZZwIWTatzLRy6Hm13i/6N9WLuD1+GL
+Es1eNXoija0mKobZg/qkWcBgG6laxc+59ge4wqbIeRRK7SggogG4MpJrxxsLVLrB4DexT1ecrQ5
hxyc4vYWuQf7Z9WTBSqMMClhpPKP1+sb9/67nJe78q62I1fCs0QBu98yGB/xUl2cagh1Mb++LfWm
HuGM84wqEyd3v+AgE2jGUOKi4bg3Bb2vE8yOryB0rIV7R+tFqSG9txXqqyEcOOvW58A/ktPqcPWe
fHvS7wVD59LTxxUW/AxHE4cj2ETAezm9pGZ8il7MCsLpHPpHJzG8zuCE9IkemuLGGO6CAP+t6lZO
XtSvKszLKV16D8WtFdzayt3XvsP17we7MccYfXwL30OqrZc+Wa6hzD3E24uHgvEF91z/3xRncqd5
YwBRKigmnycCwTDcuBmefS1WaMNznNJRLKBVVeN94l3TfB44kvw53ZX6XPPOUAO/opUE7Xq4cuO+
wcznGEYgb0UGJbIU1/0vwiIx4BEgkU+P21hVslRooNSShPnaFQvFsraKTOLHehD07U4LatqW92ag
XEkrVL0pNDXACmvsJ/emDCLv1SY56hroa86A/TgYTqLPmgRIFfZoNO+aoJWMg2HVmgZOYsEW4cv9
7KftART3WQ/UuhARrYTW2eCO1DX1UyZfuq7AeBJLHetkZaEDjSTJh1yKstZEDcDxpPzr9rj9pu5o
aaiuFFWnx6wnxD6KRNOOV9nmBe5zWQ21uB5HCpc9R00NoPg4fT7gjIINE2bNOVo7M7JArCDCSNPs
kazOsj3nkHUW2USfu70cgbdIZwag4HdsC3YF0+IgT0Z8bTqlAopD6oST414klGDjKVw18JVesoli
iPtfuFqU3H3lBmLB+m+tsYdKzJ4bEsKECJq1t9urBL7/ysAk19mmBCGeLMEwPeIGjL8pWx2nnptp
TC+ptpqGwtR6pMM7HdHukv7EQEm/1Y0sgRKwpxgu7JUqzObUq8ThoJdyvA4AzDWySMTMJ6piAuIq
27FPrhQy8kN0o9Mti1xSJJb35o7aOtDJB22GNnUuEOdxNHfnfeK7iOCJG0jrrq+zKX3szVISucDQ
Dqq7GFadELCbUHNmt6dxuj8RHj+edgHkm8utjxDnpg6kMWT40GNBB1rJUOVSweRfo8nnuj0wcp9T
eO88G5v8zkv6XtW7yVIcn8hE8K8v9S6umS3eup5/IXZ2OmMgV/CS218ee9OHnAGXclGzcjfjEPvV
Tn8D9qweInMiVxuaf8l0T/cX3B/Imrk4M5fq71N5TJ6rVk91HN/g0zX4HSEoDv2FObKGWYDD1Aq8
GCTLLNwZEwhgZfsOX+pakyct994esta006mmq6KufcahGSEfZHP+kmhCdBoqs+R0voFo8n9VwYF3
bt5BqUhVn+0Egbta2hyOGEg91emoJzXnGeYXFUFW92Nz57DJbtokkaWEDy69/tBOEtuyS+7ORCvb
CoYHKojKHvhZ+bF5CFv+se5Mx2EOnWkr8/1GsaDurKoh+XjbAvmVXtMmta6/KOrEm5kWc9Roe6dU
6EvxfiiPAelGyjFSxtdBk8Z6DcogfxVQE0eI4eDkOXONEQ8nBf7TBTMIYRVp/pF9+aaDc8oKG4i6
OKdDq45lzAvvFkhUk0crZrgGLWvUfNb4wA8N2tC8Tcth9UT4qUTk4wnEDZ2VLFJT8ZwEBmq2fglg
Q2CKJoRnyIKnCMyCS+mQiCVxT3xXpiDP7yLrIZYeAa32OODvVOKt69/rYFJtjuvNi7khvZqZ9RTn
lzS32JE59PZUGfwD6cAqFgZRZUJ+8fKKi7eUalXIk22w/flFiLvkmV0ZhnyFfBv1YeXyY8si57Rv
GSWZxeOeIiffLhPCG3MKGCsylgk0+PxyiXUBiP5eJYI/LlwW7kSkRMY/vksg4r2BtUjL5SbyvZSR
SFC81ouMs0pPUVmWpmQuGSljvstqiXOJRHDtqZFLUdNPaktjYjbSInxqHsgavHaQ2vOn+P7NBq06
9h10eUnWt/K+IV2JO03/laFzdjll0ZONPpRQO2MBwHIXmipbHZ1YzrwEwnWKQyNcJHplE49ScuD+
yuWRprUHu41MjNxVEO4jYrnFPgyccAzOws/59+fns5DniOFLlXGDfzZM6l1uKUoknQvioZnA4xA2
rtbtOYLay6P8HNLpzgpn4rhoZeZmXMX46BJjkCC5Gs1JT2knqCIAagJkn2MN1nsaQZDsszbRoSiD
EabF1JgbSocr2qGofYdVf02qzz3Y2FuPMcynxBwSQOpi+ZEL9KAH72+mnOr7ZmVPlD/pR6G0VRBi
vKA3uI/kIS6Z2pDQ4VkiJeo/RICkJa5kX05DXl+pDUOmljfowfu0Y7SeqjXWFB/os4qoYSW9gKYQ
NfS7zRkRrZlpkb9fId6U6Ux99bs/uZ6uodKqIUgU8dpHO60fcL06HynUXZVf5+iDbeeqPSR0i9+e
zzPhP5lbv4zfvMHw0GdnE7WGdDxFW5Rv8y/zMRfGeOK5eajNV6pQoVEVoPmxEWMMejJzsU/j5WWl
pyVkRSEe6QiT2jfap2ByWTfsTwF7t9Qlizv+YlYUVPS9QwofIa/i/7JTDnuYTYp+5KiNMnf17i5X
gnmpPRhGlUGXqJlmn76Ei9Wet6dgPNgWQEIt90QY0ING+PUexQcfMsy9i2YDLvRNjjZyRux2CYY0
seYj5AYKTWc9st+2RxNtywhMCdDN3WmIz+3bnuf/p0jczoSqA856AcX7nCZLhh4VrIlgnSsIj0Rf
vtjAyF/mQBi1+7XJr20s/KjeNfTDQFYJhDhBAdzxu7f2NN0wSV2r5pyaG7IT4K6HqAtKoinmmyci
4Uzx4bonxHIaNSHXAsYmi7XLwv28b4CZg83WEFV91EpNLGqiBAiqGaTK/Hxi2fINeqm2HY46urZ9
3IdXjM56iVhDalcEaG2zhMedINaL0A1s939Nml9v4XgOtguqLKMMyx41TwJiAg+mba0KuOCOw86g
RC5Lycnz84fHMpwPzDFwsMYDqYHSn7RtjkCDfS4ilXGLtrfeZLtBokMhhocNp37YfSd/scTuK2oX
hgn1yYPyYczbmtVzErdiLUpY6fXagVZM6EP12WC3il/qcZBnpvqHibedtr1iBt3NkqWhmPn2ERDO
LEcwXdPkYnbJUXXjeVnfWq0yR5K4N7xlRs+T/8EWJJfHyngXFffYY4znAmaska2ThJ2+fhRZ6UFj
D1J+3elnF5nCYiPWsfPxvG7ssP6kLjzFBAtcbNm9JFOoqg5Z6n5EdyXqoUd2exzl365rCVop9vDz
WqmL7A8q9nH6wM8sUSREQnBIdqiv6NDnwia4FIhjiyc58Gn2VRRfj5radw/hi3QaxBZ+MbQjX9Za
DdT22oTP3EXXi8TjUNRhlUmhCeM6HqJSWmXWfW8FsHmKRNUG5gZKFFDQns3KgLUjZlv3z9kPjNjh
6wB8pRCcdaXDGNavXoNsGeaPGhTXeKlkTDGYlWrz30MN7Cv1puX4vGRzJ7O6KtK/6wlz9+2xqphX
eQPXJ/+ltHPhQYP3qSB+OvHspp+br0G3hPX9t4WGGKF12yBBSdf1EEN3xN4EHabW7F61Y6MCy9Ez
zD6wRIT8t2hFQPno5jJzd0kKELGNytuo54/6mJ2iCPJVM4r8htvvRDX4chziPkAqyKkDOL1u5Pz/
AFJHuO40XGTIQRWMl6NVQrbIGjJd+mdUXmYVyAmFu/7Mqdbcr6AjSNNNPQmIG6I1cNzLV80YV1Vq
IsIg1isxj6CPCamibuA+n5NcEYNAZHqroZE1BS+Rjl+L0TxVtwZ0tmokS/qEPGpboDZoHcIFJ6/I
Fkv2FpAY9KI25HqIWZVKnljtk4CVZb9/lEKXtjrLNmfQOHO/yIw8Sq4rIUFHe2Qi2cUC841PXuG5
UCC/224Nj1hZnRsd2bJank6lZk1N7vtQIcs8TU5pyFMH7aQFxDnxQIb9lD38MG0cEQruNNkMa4ae
xTmX3LX2ydIcd6QbyfGwKiKmu8sXH6P7hftBvki9iO3ICVMvCpTK20evCikpCDXDmclO0FRqjMy2
YyG39EM0qv4XbdotfjXznZLy0Qm+krOFeKUxLuseqqPocJBKJtrDRCuZJFNVt60Vf5buP9WsIr0+
hFDpyQ7QN6i9ZWq5OeWMDK0cTfu9Oz/POVi01A9a/S0MsR+jttEB1N4jmyrMCKwwzS9YBVtileqn
SP9MRo4bLe5Tc5DLIhwDTyNlnROjcnZ3q8zyk2taQGpCDAAtxSvP8Nxdxa26Z0pIFvRNNGIYVU+t
8LA3FwSVQth++JMo3tPlSKGzr9p2eIfn3O6UkUHouvJmbL+vh30eI7+PbeMEVWCrOyN1/VApYg6b
wXhVYvWTAf8mnhPQOil5IosHHt+WD1oPF1GRdXjFloyzCdJiP8b2mYY3tmgO9tevJ5UcQUDKQxln
N+xejo+bSLvn4pfDRyFkC4qTUujzJejCaZqK1gl++qeUu5kk8QEvqITZuBB0j2S7bpNvSlmgLYbr
69iBN93PJ+lsN9MVBe+GuxVmBcCSviF9MrRxcPFUZtYxwq2WClXB/kpBzYjHQTujvl+bDFyXHJ9p
U/5PCp6xAhu7u1pXPRrYoIRlCOWiA7aPzHYWQCYvs6q0/LxpLNcxuVqugDa6dfxE8Rk+YXa24HNc
OqMk9voW/kaYwjoujhTJO6Tm0OCWvL709E7hESzOJ8F7w+wiHx3WeIr5mi/nmVy2kcTPR6JX6Tiz
kYtuSGDewOdIT+yIemVRboLFJLPHBYU13hoJ3L/ad+nM4xfnikTFNPdet8TsGEAtyhSev7iTHbGf
WVZ7pQcwYNb+y6SSzIo1qHpZ2liMqt4FTwfG5dCR42wKQNLi5pgmSjWuoXYeuRfP/xgIaFF1jOZL
ED+xk9c3wtN5Yo650TXGusDMKyQLIYGBuDySCQ7b3ZGWw/VYBYvWRm9wln3/Egq+uVmFzOxw02Op
uz0b9uW7+a4a50blWKbVEVoaVwyX+Zluf0u41CIyAgW8d1SYKQiXrpLXgo2ciPcB6inM0ySoFJ+b
6VzZQq+KN69YGioi+71dYjsfWEW3lwbvxjVY6PFlcGiecrGNUgAzd03F6b3QYQtVAJ7P0JDdCc+0
o33cxI06kE63DijPiIqtHYthUf7wzJg/y7NcYsNHPIOyzF7eRv86FfOJvjhbrXx0vtS5RznAYWGf
LbSZDku47dQqNyVDOohegxF4XEAbwOFuttfWnhUpQrrEpORUCcBrC4u114CmOM0MnLK7QSSF1DpL
fOukPYZL4N7klzOZcRKKrM5k2n/MeUf3TGYrGO8Z8fyEngRL0qoQp7nVTrF61KyoODLzl5QWg3FF
wFnKJsTeQtB5OlRtAqfNc+cpH4ncyw3aY+ZiWG4gC/xn8ApqfMkQESLBd9GvGjMcYNc2XIaynVsP
2UBnzARnxYQB/MxTRraYoCNoIKe/qB9+UzWKZKCsstsNHq+HCwfi5wfr0NBuxfMMSV1OdW7Lx7Xb
Zanj6VEkT1847j9k513eH3bTQSYC5ZkCNSX/16KY0kvcwzOy1aISttxni31CKl5MjfmXHncDykXH
KOWxB1QoQnaWvRgI0duOco89DfNTSRVCY0B1Y5sEpIaXIVbEjH1vz910tbysoECaj8CSE1+Rc9SB
n0vrq3BsVYr5jCZCh9TBF7EbPpb2M/6zydFcT/kCXzgod2PJMgXqiV1yRS3Wb1cySqPNjJl0obYj
e1UXf5TzpPY+Ye0dGd2XEzFGcNQtjCiw760Iclng0HMyy2rU8LY7/uEZEVzbEbXNoqcv5gBb2a4j
+ggHppKido9BDeVH2na3+6YWciQ/bJaUNSY6nO9W/27MoedPfYTtC34Ive2FFIg3w4AoConlSH2W
qegUOeTN5IHxyXrSPNDSPk/fBBj51W34JaswMHU4CVXEYvLKLEOykLY9z4vsrb26/lSaUcEjbOmt
KL6yOKe3CdRy3lPQxDasUXazbq8gCPN3PBPd6Xs8EmpVF8PxPXY+MSiH4nglqzis775OjLWBZmop
L62zlalNy3UJkH0PKl/ca2kQJEpNz3mY2oojIuCcAmVizbW1zj0g4fM6FNL04ShmpQ+slm/STO1W
6y01P/32jyHISMhKINQTph24CAolhkLt8VYbftUjLtjhJSsjBAH6BS/tMD4N1ehY01MO1t50hXX6
ao2VDUYeuGRGCQRivHOQehEv3kG1GwMThuD8XEqDa8Jso88SwdqXHOg5Vc3lC3DRb90NTNhEaz37
DhRQCK65ghKRjZAw1kkz34uwBRBVJ0thHqqKVxPhJXtuikUa3TLM3wM3kS5XqPsgdt8SxSHQE+FY
/9GJiKK8WPd+FqalkmbNzZZvdMNjOVsNyG6wBqxC76/MYH1AQ5ugd5Sg/gAM09ttK7mNO96xI+QB
cd837Stq/QjhLytWr5sqiqv9M6jR+B/lbsKtlXIX39pwj8VGoQ4hR2n7R/isb2XpO7w3yegUVTV1
vEQ1pHIxLH2VTjHOdgvElOcO9sa8xpzBPOQj0buyEGVLfVPS5xPrLY+8B57uitF9t1M8DXGOby8n
pg6Dm50hgyONsDDDCrT4ekBfFgZr+I+cKR0ipeY6aSOLEg0eURxzv5FPLuanSQ02lthQLNV6t5+a
qWCRihkC5AawKzCrcIltVdVHhCBOEj9Cx2B9To7t0HVjpNg7NfZciLH3/sxIeBsLbASUZmNMA3rq
PuBCj0MjWZQO+nklXPN0KpQB58X3AgACcIlOWQZdJhYXNayrxmDMyw8BgsUaKQVbfLloyp6RuHS/
ByQJnmOeqFRF5SBM3Nc2MWDLVPG/jdKXjzM5noJpLWrvB4VIL+iwzBBPUBbfGgJsrxvZ0yk4bI2d
abR73FVWbDCpwEwcXv4IUgSs72HylsiFosckyQYI/8NymBPinZmcOHS3Ja1etHquxQxzrDdIk4Wo
1TgSDrxOwWFNwos9km8ah2VJRSnThYl3xPMBPoqUYmT/1FQIkry9l2ccigK7VjWZg86yl3ReDlFE
91DVLQ27s+tHgD6ZYZNDJa7+zkvOaW5KErr8RxC1L7NLRWTMR6OwG5yOHcdj3wiu+DeXDhC/31d/
tRq8/tNwiTSIm1tyQl7sfgtf0JSUn304FI5nVewi903ducjy66mUXXuJXIWrRD4UkE9wrFp4nrwa
p1HYRXOIjzlF4HnPTsERqzgvqsAo59SuFi/5LBnPQg78xcph6n+vhT7lrhRC7Trz+TYmaMNglnvA
sWrVVrkaMi2w/0IDFkSzyEANvIygVU3eSmQxTMpf/8jXlVq3XvOTunfP1zIwcPUD51SVkmkEizHI
TfbWKujX8adrd8ic/XQBVbT2wfJFnUL3BBE5b0YDxCG1DcdSSbD2rzD3+uD7bJ1tOnUrZ63aQbSs
t1Ag5hZqkJql3YF69aNUN2HlVIxjD0gwUtMJg/uEYRetep5j3H5a1vzEVqBL+7+aMMvhARHwJ8oB
efKDITyYaQJEczsoKZzr/tQ6ohu7zK5HrDpKkzzwO2Fvqk2PI6ZfxmT30IR/7KI6JWeXMefkSgBr
dzPUrXCLB4RA1r4SRAdpa0Bv2Mq0aQMycSWixJ3yDf3IUhH/oKn7Z2L9xswhwKLk7Ba1Bi8Y5X3q
EtbB4dYzY2n9nfu5HdNONkzGArqINkmQH4PvYVIi3/cmht+9cI0d1lQHgNJnaNzw4VE/yJaqCeG0
tXjLaQWAm6062ny0iXc0wo5gTBm/a98dZmVTNVd5xMPeVbGMRLjXVSXxtepmCWYo0UP2O2fDh398
znVOYbwdEcVdRYm0Qb7vWp+ts+WuwWc2T/FLwICONUfEUSNK5NEHFSk6QZRihST2wQT06ceYdF3O
AOjsc3zWJrr62ITOCjxivBZMDeLyuXYiTnOWZiDXWZjnVpn7AAEUL5FioCg2mC3jwpYNS0UhNVNK
e1zuxiadQj6JMfjh+rFYR85SN6Luhw4NwCZT4vFsZ8DnP7Fq9uyNcnIZRo7Ug3XbZjIsizbRZDBh
6qd9YjnEKXKnIUQA17apihCFYWX7tW9Fxmp0aGNepgldoRb30fT9svX7JWQEwkhpWXrtApQHRATX
lCI9LUOkC4OnB8z1Uj+EKIqmqeVj6Bgd3yjDrbRNyx6U7bwNGpqBrRqK3bIg6Vbvpwr8gD8GiMK5
W7ltOSMIvtT21ogMpXBGKhRlCKNfr85BNLnWKp24PRyy1YqGkusTrZ8rWbKB6sxFx1b+oI+j67nk
jFeA4+yEl7ZL4XIBffOOZCL1dvi/3CrHICBPEtStu9QcXVCp2timOHTt9x8SDbFTmx2CJOGA4FsG
8ba+bsvmghbhvoLd8mFoePWfMXzJph81XnwDB3SIrKrfMpyr/+SQPuVjkBG5n69zVn4B99mHOTqc
eV7zNC3s0H1d4wnRR7zCKURDIZZR8q5qPRcAGd+3M1o6+sEsgnSCdIYyV6YifJ3jxlq4BbIdWMSo
y4pEdY5qojMHSDTxos8cAmppovkFwjh3YDz4fktmGhCkOwpZk23y9FTERBxKOkNmWDac2/tOWUkY
2ydfPpUJDegt9LChUoZPNLMUpCAjKSiOcW8E8aaWUexu7LKZPFZLZn3AhMXKDIzEASNBbM/js7pR
2YZh5sT5CDwCIOj0kzwqBRl5pUjlyuWJ/IkT4lYuGyu2+s9odR7YWfi+6YKdrQMRG0aY7Ds7BKUF
1f/o3WA4wBHXhcki5cWCjiMq4z+6gUpvDj4ssPgHP+v18sHNZmuo1xIWisnRkgFqkZ2cZ2j2MISa
3FopgMWLj5HNW8HQsTs7LrStxKKQNuSrY0nNk0DjR3dd7YjbjqT0Mr4ZmgD4P19S8HB8tjblYtMI
gCq55N49NcwYJo/TLxKMOZhXGBL8EXp0omPDjbEFam8IhjL8gBpLNQkUSMuisDdA6mAFNxExaBIb
nqKXNyQ4keRYPrpvLGBtQ0m1Pi/OO3fqcmC2WMGCl55KLwykDDbGUERkzBW+C0O/WGFidfRDB7xf
C1jVPLdbWX67pSHe3aG4nP+0iDB4LjnCct/N1aiZ/VcERa18qLRy+pnjzENHcADG4TCZwlN3/UGp
0aHC7btxrHOKh6CdW2ELqbF2HlBr1QnG0v/5xy7QOmYCDrPgepaFJh4FQOZnaDUjPu5WXFDrsoKj
5gq2BRYU3AdvYCfWb6EtnUZ4VgbuuQaLslognLY3Af619O6hZu/LODsYwGoheYNNH+5Tp9oCMN7v
2EBCPorQDaUGqVntPwJJOuv1uuBanK1j5Px4kdBzILUkAExgu+EKBjrdy9YVrgLH2LsBJT4MCZSb
5NvDnWUqF5pLV9C9P4YSPxlIkgLXeMvO5mHRzyoWzvKNfkobSEj1Q5ve/58Nkr5yuD+/gCMc09Yb
iPAMGSQQBqpAfpnwb7omL7DuvIq9Ew/X+BPblixhwc9Zh2MtIK6xwcQpDeNUotPy5priQ+TBaKpK
mB37dUVd3gtoy2dAyvB+1aCwuois1QFeVfXhRRwwom3b6mBFphh9VRomi/KAv8CPwSvcg2IQXB8X
dvkDDh7W38j67EdyKHdn+F2euXtLnewEyd0cc4wTKWYX0kmNrvCFpOlLtvM1OKXKWLf6nQ01Ohay
3cbKsWxLDboJYjGtFRcDLLl/ZllH0+7EjLe9On9GOqdk/NiXp57Etl7lKHmcUlvGB29VVQ6QVb+o
sISTiVKpFMjmlXnOA65vVtQ1SylN7zRHC6O/+ItkJxiZ8A0TlfbjvFuPlaRTWMGMjp0uPLHB8uKZ
qK13q7jcVqyrmjfgnVuHL2dCOgjR2Lg0ZYZo8UJO58RX20MNFV29m3mj1ATfRBUTlW0ELMa34yRG
w30PF4vrZFRHd8VotQysoWt+QnASRZuX5ntp3wsxb4MFqXh3ZdYUxVVHu3gykwmvoUhgqw0gLwXN
7p0B61RuD/elm5uY9m4bvj6ok7chQOWur2fUUDTxFMhbPozVp/wevHDuGOiqQy5zvUMegCx2nsyM
+pUvLEvJwSgmqRhv+iS22pKBKdWmR5ikmb2YPG+t+MUDy1PLR3Ctd/D7MGhCufP/UMpr5Vwqhukd
bHKi+OHLX08/TMxncfNIP+JPS3BQnrCm7VGR65hSiSX/8h2MqNXMvne6YPX0LnE7vpdKWVtrooVw
KHR2IZhlr7WpxWEB9J2ugUzOo9jtseX2aB5dkNhpwSoBnE7Mz+KUQWXDoouL2Ug82++3icN+zI2u
w5Qg61DqiCJCGKmnTqxviw8nNyXbnCKLEDaN+NZUUq4wlXsr1gvUPgKFPUn+CfgBT1WosbBkQZda
itjbTPGY0WBdaIp3eikXoPVluqFPSXaBgczP22auBvSuwhuR/H3MW6b2M8PZL3j4zLYXFnSIzPus
mq/2jtsOSWLXRbeNI4lW1gJG/sPPBSFjRjSJvO+YwGrklPSW0Pvskth4Adbk/rRlH9hm1jPHptU/
W9W4hvImrd1WUAIC9cNehHdeKbf3ftrgleY8Z/JndKqEUvQz4+wLFx6pTZNSheGWtpVd0giwSZcR
pzNYwofcrBSDhEl53udY1qC/4C3gKzoBBHHVW1H4jbjxYGP2l4VO/qgG03Zv80PkDsVLVupnJh9k
D5ff1qML0CdshEdeDUxAzbyjb9bSpbqRPCAOS2l0U1tACKuhz9ST/CfnnNdCq/zjoW39CdgL38iE
2CO5W0QdhbQNBhTr4Ut3epwmqu+fy9uzQ55hcglFQ6NO7wGM3kAoJThh3Po9dSakNgaw2oWzuHl+
smxdz5Peynh9qvcR1XZB6UYU+vKrilK+LNyoot/jQaDHRh+wtuh0oVxn50/ihEfql+O1k+2wbUFo
m84uHRUIOSYDGZmGpuuVLYHoKTMTLvi+StIqzU6U8yOlMUtcm/vl2qq8nvq8KIRhAR4JZ7nyCpLS
wMILDfN+0qD9xU52vnIsTFk23e6FhV2/OvNd95nb7FFnT0Dl+iMbYjs5KXl2dmJhxsCC5Uva4/am
xgFhidlyy3dsSM1mukK/dcFQ7tsLGMsSa8xH0dMep/rK/C4eSV1HxDoyCICPW4Gjthec4uOJOnXq
kHBej8cmx58ND0VpwsEG3hRh0HaQB/BF+dAvSlspFpQFKN8Qfu3xXrdMuKaE+5ca7WgW0ZvLDt4S
kFMrHyzybqbRhA+YhBZfi5whlzNwkY0O+iHGuROzZFqWMrlHxOxEctaLWzXJhNj/0nXHxBFYiQrI
QN/FO4NsoYhsTSG9drT/ERC/pqs4ifkh663/+/3aDuUqwi/F/zgJppsYhg2uneO2GSiWnEp8hotv
D9FFEsjzpkyec9VUX31FZ6HCBzNpPw3m6ofvJid5LqzKp4h04M52/u+PErKzCDF2MSjjij4oKMex
aE3heTi6V8ea2aXTboeZog43jLQQmqN0fPvit2Q2RykWQDlAci8PTvLFAmNg+HSA3CvrLSs17WoZ
WyNp5dMFILvdPK9Kf/kXaJ6bpUrlbSU3oMbSAhyGVcxBhOi9fvBeX4voK7IzSb/+yGdER1x3Y6v+
mauRy2cO2f5tPXjE44aHnBHrGhqEs4LXHzArTtJvgr+v6Hr6ZvtZEC9ar6L15DbxtbNbLPM7h4ye
4BaYVhADIErIp0bdOwzMIGuYafS8S8hovSKZMEvsvhNEdvYABH9hnPZKr8S/2sjzctkQ9BBZWXoj
oTdrGGlIt3GI9O1vwHZU48enmCEAI6dO0CadYYlMrE0yRUJgfNNaiY/YyYjsWPcxdWMzLE6cXKey
cB5QDkbm4k+0yYJa97nOvYd5bKt0DAHxF4kLoi1r0zbtsGdOSu2+zb/+ZgaIihSLo/0V2EDJcnqD
omnJ7io3wVzPeSIcGaUWvvovUvTn6gvDo/UVIuKCnf+WSGr7xeEi3awkmBRt4ZI02jQDtDS0W4aK
BrngZ9R524mnf7d/bBOr8LEzy3GZzAc6y/rIg1Ccu6Qr5YpX7IjwPgJwvEtXfSdBl59mVxPHwfBy
8C/SNsXNDYj5QO7tWY1vF27ITRelt8ucRoF8znXX8bsA5jkt4eobNPrmFNL/UKhO2Lnc/z0B6XjD
2lmff+VSQNnbvSRIhW4iKDWhF5wPuQwiA05UysLPWJ3jEnyTu57aCPmmS/nBoz9mTEfNVpRWITj2
yjO6pLXpFutLzztaNk2iRPs4Z8ixFZ4OHQmvAfCPsJq3GmTjA1pgmHoOpP/C/xvUPt0tvY5M+14A
9bFVY5fIEOJqiaWGGEIBbuNZUs0tM8rEP3qbX39BYWp6p9u5tXCeGIfXgskCCqCtu76UQ2IHWA4B
ME+fN6KPSiBxjbz4W6mCfq125fjGWVcZtEI66POPiPLs0PzO36NlNFzWKaGjQW2biwlt16sSxCp6
4lVD0nLGn20FsUT4zN2jdTP6/f6AyiHiL5sIImbyvmPDljoNBhPXc96Kcewz2TrP4NnQQsjcUYvF
tHXP8PBRAZsUdBOCjLYX8RwygiOKgWy4tsaf41HcqD0ipbf9lCxWBYMQca/qt21aEuNq28ylsE4l
ZY+RO5euxSejgOUI7U1x2QF4YnBF2+bpnObzpYNjTUWAwo/B6oUQiBQPZdlrDOc8P3vjWCQQv0fC
VqcsUCaXkmb/uSKtyK3o2+xBz3spUZ7C78xf7+VUBKBn9FRUft1ldAESwPFlTHXqR752kyng9dGP
7iI1oWWDWasYBxcZFMMvOSE02EiFiZwibNsxIelbpp8GC5OUYjDxFL+FkaLKVZJqmlf+9rn5IEWx
Wq04xER2J+3WVOY/jPLy4wFgkBb3faZmYRFAGyxkTxZw9dLUm6g7VOxmtR0itoy+diWk+9m8wtpJ
fSKNKZhAPiunPqicC2Ayx9pORdVzCA98nrCf1w0/nCfG9kAAcvhrwbIiQ9AVtWqnLa2bDQIJquJn
oUxYWwO9fNzzMlcV+ZzTRGl/8iMOzf68KDVoOrOAlfbCnYWUox7mPqLnfkBCxG/siB0LJ/mbGZFc
4TlJfMkPf4+91qLy88zfCJjdmN4SNbkI3jydjKJ9Q9u1pY0CRV13xlrzJwFtkIvFzIxjDItzw0Eb
8YL5locXS4hdtjvr+Ypg5nQCX1CqTbQM5MT/tIRlP0PvvBW4HxelwKAOrdG/ta8IOi9EV0g0TmnH
IkTjfaVas6SjE0cqeWg53I+Kaf3a6hzONRg8BjNej+l/T7ycNM4ptwGUALJuSUapWizTFgzRR2os
GnaJ6bl48+aYCSEch/ujDHGGt/L0Y6NTSN3yQDCJ7KLLU3jbiBFJ2z9uK0gQ1wVKFZ1lJNLH01M9
nvUCDokbTHGcn1d4D6bTmZVEkicbUynBd+j+Ae3XTRZler2cqcY6TpRYeZ0KGSNRIZ0XUKknLMj7
0G0SbYPfbLnesZD9XhecX3czWQWwveAczvdOu5FLghgz1mySZxxXkNMAx+9MCYTaCrQHeP+g2N41
o7Gt/GSw0ZXZr0coiNhS8dthR3YQ2qTh0jn+d47i0LNBFf6ocuFmxsY0Z+jrMxhQJhwWJBvKa/He
+hsfUNN7orKtp/IUm8FdrzsiLVyVC5JyTESN03BY3ENoBxkktguyDtnwZk35K/3XDAMNCS6jMfw0
vNuiDMZIa3QEONuqAoag3MK5nFIqJs8WGL6yDKzoSaMqgR13tdV1v7L5ECNk80uwXrOmOc2jZXgM
Rfqa1Hj91iY2IWnQsYvfGqT3cf3jp+zVVj7nOFe16XeFkCQVC9ont8EIN1mTdgq8MjYIVqIndGFH
WwVYkV7l3eqbxjmlWwgskYR0fxM1JRoM7iyIvG6zj40SdD5DffaNoNvJOJy4xRmm36Op3e11JO0C
ztQxIsx9MvNtNzBdFgzvW/cPbJ/vlw97Ay0WrHaggWUihpvArwnTB+fXhLtlD5ZSCxPCpW4fEgcJ
PTgJMWyQxFQUQU6bRC/QMSk38JAQJUlXZ3qrK7JX2ck73ro0vDbQnhsEN0814gfrD02ggMp2EPKA
WpnJ9n/8ckqAy8gV2/6FiddKOtH+0oeVBUBqeXdOX8m3GVZbztNiOUSOGY04fWcLpeBj+0wj21nu
/pY41aCxel4oJpzZyv6BMf79Ktp6pgXA17+6LC+y04Uh/qSCPJm88upL4p/3GtdHZ6mjBVqLOrL2
8ZnQymWN/rmXdzgL26vWFZqmPyMlHaXZrqV77zMuJ3U39nCP8x0moE9utGO2gsg14jbIssw6sPHN
L39rV151M3MSdU0UPmyDon6yUpNj8P5ElckxJHf4oqBIjm42D6f87K8+UHyTS4zBWpndG12lpL19
McECqX3PdpR3D+dv3MVrct4p0xG/durUZ0hJHyxcu7yUZI5h3NrLtaQh8ZTQcmiMRuSMEW5ARmGy
LoCQIQoJLld0GqWOMKaXbb+FGejDwTedNPa7ivpD+yppTUGL5dpCzHeoR7rROKbBX4ZtYnSyg8Jo
LQasidgmCKzZNrXwUfADcwuSFBSW4I81jMXnPWwacrKdXeai375BcsYsfeLek3bETvrKhvJsAtZG
h3aXp7bGP8QTCZ2YXDyzUyhPuqkEeHNMBgYqeW3MTwPEoCxqDMF+p8AEde6rPLFzQpQadLsVw3kD
M6mXlGAG5+IjSh3nzoijeDoAML03QfTquuEedi9LWC5pTqphNwW1IjWA0bsYFlbxvfIUxEovAY6I
r7XQ3Mds2R/KOXNLY0bR6tP8Hc38vKLhQe1L1cUtlpS4f0ctzHefIB8QWup8TYti9YHkpBSaO6o6
T5UNuyn3Hm7j2jBn0gWDcstQZ0gVGaJy9GPzSgnC/kILQltblQMbe5MRYg4ngYJzDOlJSh5G71S0
JAsfnEFZhXAK52FjSvz1zZ3asvE380r+6Cm6/NMLb0FxVU0CJoQUNfDhI7WX8XoHdCzlq9ONTFl0
lDQnIObbWLybI6a8F1VIGjxa/iKir8NoTqCtUfFfcL57nZ9qKrkjDoJBdLJGm6wxWs7fnt2fxRnT
7P4opt8IdQ0TukOSzuD7CV4xYUOAozCbEBM3AhBgUC02JAcWo/HYTTxueDGkRAiViuT8pieZFhDu
Cyq//PhGPby3kqNz8Y3QSQR8jdJp/KsB8eelzpBcKBpSArteehIdMD12eje4bo3nRRP+VYX6WjXL
QiLHJ8BRSAHRmROb/IL2vvbky7zYqc3+djvPHL9PTm8BDdoqB8Gi6OuGsszkCRsLSrDiuop31LTr
onGNXZqOnlEURFEkYVhUEFF1WuAZfP+2NV+1G/jdL893S0/jIpEH3qesjX4b9MEM9Swsd++BhMEu
3QA/GLm0I5qkoHAJlbn+IDtygqUzWot5OsqLQa29DlGWtTLo/B/YRklgla3TFznfkNiXJV+bfQ8u
9VzwgErRQ7g6OhUX462/G9iUCDBzSbYrAzK1oqnoSNMJBulB5ws/hlphE2Vkdbt8BAEyXMUXuFrg
XsGypGpLBumfuAIwWdGfimwDl6cifxS6f4Qm1GOZ2zMdJOsGH9BtVlnSLm6z27uFlBAC9Arz9WT4
rKiX9i/w8g8Soom31pSPnRfMPgV+eblxv4dvCf/IE1+EHxDkIiGAqxxJnOgME3WpOBzyDy4kVBN2
VhBwptDqzMCvTTK0kmhTKmDNlR3ue+5KLc1oyrpwxWXJ7Azcf/qlbDDb7VJ1+7w2g2U8uXIF9iBw
rV9rwxxVpHb17U91PhTe6rzFUpswNpejesF+GRYKFlahWi8R+aW0tARACW+5cxFvYO/0fh/SnRrF
C8MDMDv46SCEryfCP/ygx09FUOUYtb+Nfs6zP13GBBIgiAlsUheLcjRkVIt4DudUj7JvsDRr5foT
LdKDwb7XUnLH32adqgO+BH1P1pdwn0JnIu/Cc+ReLUKEHLzw964oH3sjWUalv+2ZAy2VZObmEn7Q
YtHUTsDB+e+0wFxb38k1Y/nZ88PhK7kmGshAbpWD7ujoFaf4JaFIxL/8BWsRFimoyBDzxTQDl8Ia
D/UV5q6y1bKhPfLlcIYRs67P584u5xHG/lqtZqoDWL8NS8IwdDbeFs6qibS+mEGtsgDJuOkJXMlT
6r3Z45SBCOgCyzY0T4idkT25RvMSudu8+XMa7WdFc/JqpHTuBSv6qd1lytrhFXGqnWyaw6htT1J4
y7QGz9idc7Oyqdn3iD4n0UJpZ9lcy/4E+gd7RuyLRbLod86JsHlR8yZ2397V0b8R3MRcVdld9ZCM
y0VcKg4EfyLS7iIcAPPgKgC10awsuk0wFY7yYtxu9jTPdZHyAcnQTCqAUGnBBN9BB1LUaAwuCtK1
6huEBenlmx6Ql68zn0Lmkrw/gOBC9JtvaJTmrkPnK9LpJMl4Mx5x51ESBkRS2FRgQzaJ3R7CfZlD
NVZ5Sxt7/nuVKW0TGFMEkxnFTBuIsd3kFtLzxUcW33v5hkXzsjZ9jtkj2aKkEotPAE0zZ6GFqjXM
mvPHAaM5SWh2okl+ODgiXNbAwBKa0X2InGGcc4TOCJjDdgjGaEhqbi8W1V4267BB2fpYPw7i+HAa
B7N3dO4ckG0UoNuNVWWzUf20xK1Af6sIT/LPv75Jufq0U016oeqTYEzxbWnlJM/6YS6BZATrxyPd
pk3vE2JD/JD+2a8rvKjmDlrg0YVbIvtfqJUZtzf0k8s9FlkJTNGtvnUTRLaKJu1MEbDTN/6Gw0G1
4SfLCmqX38iDj2F5+7tJyyTBxWBjYg7n+IMfs2nipc3RzsD+IYMy8pKkpZlFTyCqdP7XNpyteRIH
FVikpSe/802OINcN3+Hedrme9BvlcHJc/w4xnGxjdqEIQmZ3zZafK9OKzdaTlnMRTPIC2ivpTqae
T2+LQ1lWwmdc6bkE/bCBQb7DfL20rh+iseYoDlne/LDf1dDH+EGNr31StTCZmXkUd9FJoayZ9TXw
pMKcbABfSCHNjM+a+MTZJcsAkqo+bsV8+7YatcM1tEc9y9E9tHF4A+FQkVCYRxTAhunhb0A0T3lY
8T9Hz5yTxG0edVq+ZhdckL+U9PmwN13v1dCqN6ZmwvZ7jnlyA4fjL05xYrcJBngEPkhFusIYm9FW
QBhTlYYMd6NyPKem33gPyWKSQ4aW1ZEK6Y9uRbLsomWSAb4oUX2i9HJRVyvX1rcZbuph+d0g+XAu
dAk1ZQokiuel6VMbvOZ5qKG0OQ7nG+Rjw/Y5mPu6tez4LAQpEmI9TeUO/QS8maDPxJJggr+5XlvM
hSX6QUEy/wkYPyqCG3N1B4yJf+1qZg2kty8bHAaHL1yHi2eZQ8g1KED7Wd9gW/izuGYRyKuiWXOk
u9G7pblxreLfOaTEQX74cqOIUF9gzOWZgj4vOZN+wu/+guj+dU1lHJuG/2zZaluzPOfcDRS9vOD5
3O3s6amfr0EzhmFie8yrw4qWyDfOOg1T3oEO7skvkB0h7ibKvfUiGcwUEl347ZPSNl0DfHv5gdSM
JfjDE+C+SJCYVGZU9Qkh0UXvEV+NoMRWJR8qA+EBoj3ebxDeiTwALz1g6636pHKsK+vYHkCftKL/
yAquqWhHxS2DrzYX8dTk3pjteSR0wt9m2OU9uG+HUmF+ywbeTdgCO1yKtB6rFLJ/WcefD51mTNBK
WTij4sCq0hw5nTK0s4XVOTVk6qMwcGJmChtFw6KRQIGfKB8mNI6lzHTQQZVom4T4v1IxohEvzJu+
rEtG4yBPbFFnN96EQ11cNwzOpWDWKf5lI2dOW3S6NfV/epcK7G87DkwAAICNO0YBoKXCgVJYIWp5
dcEZ0btoD19oADZS+hX+wGaL1JzhHaA8ZD+xLQXIjokUEEbduKBMqojQZx7ICIZ0hY34QBm8ys4a
kFDxYunjSXQYIOzKOr1fddPfsYd+Os0B/rVhyBi+GQ9s6ds2n1VZmLeTV35wl/ZYNtkiG2eCA0S3
kphTJmBGeGg7BWFYg7dgev1cc9tws+xqq9buiJdF7J/JayZXPP4dGI0zuzcGUitXg0KquOtleUgA
UkabA7qvp0VQn5zbn6rNU1QaeKGjqIHpqHJbUhWJ/lKhnr0rBm1zO5vszbdqbGja02xxIrObnOwo
dh3O3JHOLuqZdLFoT+Q56B1RW/tWX/qT1kYLpeZhBWrnbl9mPTqv+BFKEtjkP+lPPwUXlV33tTOK
g1keVi4haKXYDDv2DxJms6ftDSnuxOdZBnB/lhzeR4vL17PO96t1t+yfeio63aU/yutbymAAnHGT
z388HG4rjpviznVy2oTeux1exV/xALCtIsLwXC0DVnE++F1vLrp0rAQrlZ2RpD5c5R1Z7PoOfjoR
a8loqAlisR7Q0Jm8laF3udyf4bXwvDEB75WE/XwTeHua+CGudl5lTtlAR6teNPyPoE0RACIxDTeQ
5rV2CjTXH/kYNKZdjd8j+4co269XFk/jd+ROE79EJz7lB9vn4M688c0425YdgjGFg6+ppF6VUmlE
GlD6NzX65iFqfEiRNoLY93Grr0GbUeLbh5MFIUBdcvO7d1v/Ps1Vj6pKifLPuYyn6wd/+v2h+vL/
KbQkUmm+u0HFOAWquomuGbnyGgdV4a7OvOZGJI61x0cl1wJYrd6uIWMpxfTIhR4RCpyumXbqBQ4C
ThzlQXaBXJjZ/3hyOMLf7H4gtYbaNAvJc91O8jI9WUGIxaj8JUK7npjzL8RuM4pBLThQd/1XA1Is
9m5tPy2hVJvtw1Pgc5CGNiHoAS0z0WBRBKvmVMvRSq1L9/CpmPBb3LKQgSe9BOwbPhmnd/OPvMaH
ayRpa6a0a+pa0vgR5K8wdyl8z9Si/DewBwNNx0aJuhmSjk0iSpM82UxMVagdiXZI1EtyPRxabOXq
A19gO7MQSnvD8udn9lIdyTlWc3hj9ELLbaH62ODwHR5WrZLEHBWgHVsEAB4PeVaqMr8HLjgW4FK+
5cGbhPROTPPeXZZosTdVXa2N6Zj8FRZ0Esjrv8AAPU/gbTPgDgHpMLMFA+g+7tM1Eg7DR4JbVDqg
q+XQuC9GQnWJ/GKym8/u0hcs5bUUa842s4Pl7efAGGA3dlpgFm56UegzFS7+Z1Gp4+ZDFKBigQ/a
U9GD9xlOhGqqbBdtzkc/tEbH1ugQZGLreIJ088RIblWvCpoLK1soXqyqZlZZdxRWdEoTvrCo/9/J
kebLXF6IL9VX/fbwBJ6DZsiR+du1soCLOlN8ZrCbmXJx+n7GCQSOpE42s08NYRjIpiSsG1TMi7ZQ
/JeVeQ/RjhUkxFNXa8688TEcu71HROEQKu2ZDi1bjZPM221M4QZFc6NfgaRxBbQ3HohBl9YsesL+
RT4xEXPBOLtk1xf4YZMWRilnZnNW+68LIXI4p7cKXuPICQV6e5zEF5thYAUyZVAQkeOqTYGWr0L1
n40JZSCdi6F44L2mUe7nV8PKAwN89dEKdnlzOkEbXZD9DnFonfO03pA7hqknCNz/Lvk2gnCO9v5f
M0Z3ZdyWG2lB2vlsYgP8Ks5mY89/nXf860bvYum9kelHAWELV5yv9+kJC6V2oE8zddDYoxaPApGl
OIDIx51hjrFYbeOUfcvkaTfQL6TaR832CBqwwI8KOHNfnJjCqyY6FpqxZzWdFliGg2YPNuscsz9f
FcnVLQ9Br7AmajusixaljYo6R6ajEqIXm9wk6v2p49pEkWIUWCp/LPayTsMZK+f/Pcg60lr/gBBt
/wcliG3UviOp0UzB3wrckXxZjJvBB2oXd58s1B/oSXaKsUG/vWawipf6gWZRvTxEl3I3HmFXc6pU
+wy/xKBq55LBDi7zd3byga/yCGv4POc1kDQKZWFv69DnfGRakZnCsQ4jllNtNVbVXix6fUh6hVZD
Qeisj4CQdCq1H29mnFwrPlEKG6TfRTAiuQ9O++pMaf1AH4HsUgI6qIh/gjwoaYILcu2OBb9YV6s1
wxwYcWiikQI0qbUQnyYMk9BoJIH3yE9WzKFf1hQmyTUJWUYGBdIXJzYnlOej+nG7m6183PrKfZFb
bOSS8USBUQJVmEGWMgOdJXao9wc/OEcz1v/4zMTJnlxU4EgpEzT7H5FLJt9FUnLsfqyOcUuNTwI9
WmzToeaFXYZI5/t0HwflpRG0pyNcoUmzeC/OnGQNwlvy4Jw9daafyu09kCXGeRrFLLktXd3z69aX
KxwT8adIyYrp9iBxX4UZ6Bg0xHo8x9c2VPH3MfvtfrwZiVbc6BHBsQ0/ZfHku9iNI+rbjQvOvB+y
adKR9Zbz8cOYxBXcPAQl2PYrAnCGo6mbBf9W3wqxVVJnqKDp6YTOwIwAqnTmgZJMFGttiiKyKqqk
3Ht6HliDFghjIq+Y4OHTnTWTWQuJutEcd2FBMSVz4wdUSnYhwbK1RlbG0yKH6s6jGzhF3krrryhY
0jM+FOw2on2+LrBSfamnwtIrupooNBKVd0ogWPgRD+5MPX70XRCOF7wX8WDN2F76xjkQ4vdm1lOJ
JKxxJbH01PuBOo44Md1CGxIcaQAen3EkEJ0Uh54HARupHIfzXnIBH4HDafhecZWjPM6kd7SPFusZ
cza2155+aXXuQ15GZ2tiI7vDj7RJ7bur6ULpFFnqCbRCfZ8+jOKRh8rKL2dRAguURfgbPBYHXAcg
5wnYrR4360daqWtN9S6rpDBFjvRnQNxzOYwF1abDCLdyNvKPqu1bS5aCgnTb0vtZGMaCgWBinKGr
5THCsMsT3OTV2Bd6Ap206innQabmRS/n1UHKpipDsrRZEnq/wcFSa88tDhIxncWXka171T3pyY7x
gfvUoUdveu8/aEiP6tL3Fy4WVGB6jfUMbd1zqWFE4gHyDLn1eJ5G0k8kDMiQ4k1OQrO95E6G/DMw
R/1CdPtLGLgjnQ5CCoyuU7FqUcQ8XB306QSrAcqEqc0FU0aRTpy3Ec4Vje+OEdeQvdGH/P03KGW7
QhESm02FPKwA6wyCr6zipvJwKEFZ5Mfvz5qSUuJy6zDDbGHDhs1LL3cOF2mWamjENP0ytdfnjcoi
xK5ljcxNCl8tXuZib70BwcycfgvneOeuyeHl7FHsW1ONXYwjleQrc/Z8ENxZ+V+XS0ik0fN9cYuO
Drk8lN0HM13uOfh9Ws4D0mtYiUWeWtd1NW2EGB3T5QDU0eP6Lq4Ite5NdzECpxBiBd6raDHEGSCI
1NrUhc2xgXmhmrA5a8t4Rp9qqIodEmLljFixYmLXwIutDPI0xfD5lgco0cvP3qro/jZri1qA+RG8
N4CLWX1ZP1749oj5EYXz6zLhOoIuojzqes9AF6vFTGX29AEH+5YzQK7y0OdmyTf9cBk88bIMhXdr
OC5YqE2PA94eAX39wfPrcM583ndZmrLrbCCfMKnTuzGl8BK5yKkPsmDYyJjuDj0ijKXqkBR8b24F
NNqw43FagZGRxNJk//GuR54dw3ZOMaV34zWdIGGp5qqU6fgRno2YZe0dUQDioGaZMzpO4zDTfA27
l9kjJWIu7T4//d9mbigUIZMs8Lvi80AUkLnIme5e0rgH8BFk6D6/t4uGlcOQjj1961OpKJWMHIH0
PKJZgdFicdvQwx6hen2WyCSYv0yInD57YxtFBKOHzlG8yutv0AeZGFbZPh6QKDJotfjUWS/8MNSW
ViyX4YUN2p4Gg334TJFu0XEXCnfIDU0UQnKT6mefl3aysU2FUHSAAuhJtq4L1eus/Pkkhz1lnK6D
VxoGF2YNbNptjBqZopZxc5AKe27II9Bg5jYFJfrLk38RJblhgEyHWGLMN02CHq+H1/+HJszWGzEE
hQb+BmepLMkFNSjLXTNLigsyerNn+Ds6mqHWhiqWDiQEoIy3nWxDk/BrfiiwRCU6g0J96jJ1bAoM
zxDRV+RtYQ4HOXgjUA0obbLrtYbiEJ4LhKbNUlXc+m2JMs8QS9+O0jw+HWJtXim87dsBHR5QMkqB
hJjzKpUjTc6tu3sNoZNrB1P5mMX+PJuGaOJEh0O0NYVk0qofY7fjcP0jIdObxrMKmwsutsxEKauI
Ed806ZSqrh5qkqJ/dd/xZvkq6LbkhgRF2u169Lhh0WZWxJSi6s5+1+c2fjySYbY6RXUGeVwVawVM
kwx3gFAIIHcP7Siu5LVVq4bFYt8lCGiNLugCPjLiJoefEBQE3LaSO5c/UMStaJ1zoxMBx1LHFVdI
95zm7TiH1TKdQZSLxecxtCyF6wdVgaivlSnjcpPXojQHBe9jtT1G+8z6XPgrm8LTHV6FaagGBNn+
FgvzZFRQuef2qCNtXaIh6f+LmKm0MfYRC7Sa3Kycj21yqIBLcM1jkJcnN8+kZQLGcqfaNH8QzWgj
ULwTIkB77q0vV1/DlSuJD7sjGTUEXR7h0VQIT1SgfsniSldQX1ok0JLNaRmf28V78lUn5dYHHu4W
UwOXfcV3tdk005J9ZJCiIj8sIq/vvATp+/vXbLOXVtAHdva8k45+1FAwNxLfKruheczmZNvWfzHq
jfafJ1xyOnJsOCLrarWHxlyzJU0Sx4ExJdoWijPfmpLz8MF/j9Yu12I+lg0sDQee4pYFhX/fIEVA
STbGSPl9a8tjw7bKcQpj4VWfF+2ydfQsfo+W0IPDcyGK3EPMy2nW53iLN/2EkR6DvVA+Epl96m0m
OgGbyHqCrfM5cq9YP5sqdfnEe7rx03c/afUlUkZo+llVwJK7nXpAfpzTYxCRchyg//Tdcb3MQiA5
ygfJ04lNgtfxd4cNywh/R4rQKjT6/5qK32ExlYrX1xo/1t5unncCZc/0wgLwDE0wiC/65zYCiHb/
aqgjn7Iv3/FPg39qlX1ggcBSSL3C97ZxRRiGJfhVR3iWLL8tbpw5NwRtP9NfG1FOvcZkdD2lsHQp
W3ZHGDfkt4cReahlUhQ5fRnwYK8y3xchvHNsuW/6SBsCIcqPoG+jxHKNB03W9bf9/7/TKn36U/R7
JD9rD/5zRKzm3mwN6qoVVjdOyekE+/2S6zNPp79bb6feLgOw/GkFBQ0mbb+DytQRg3M3h+4Uz9U3
BHe0GxiJF/chIyNbwlMWJF1W41FWy2baftZq4dco9m4sAyR70qXF4Gj5HzwPvE1DqQrKGGkkrFyW
jNIeOMzduSln+wy2XGbmasoQepW48fovi+4rclmBgosNVoZh5cXveOK+NJMGHUyvPNYWOy5is6HX
gaup9tDgpVQeME4QUiMOTMB467S/aHgt5G8Bo0C5xu0K491LL21hIKnkeai8UPWEPB3pC430NxLx
JU4pO/lquui1idfnOvCrCwvJGwEKj4g5/9c0OZEAUXTy1KhEkn8nzHZVhclHePPTVQHDltPCbikS
w7dWH+1ZqqNt6xfLBfuzERMfNafXTHtZE1HmT3PJ39UtzX45fOY6XbJUMxRtN3hn9csS0g3fRGKp
eBC/Ji0JnkkkwFkSm+oqBkLqSkwa0UAghrCeeFGMaT6pJEyJRNGv585esE67oBhIcxuTvNBFjJht
Town7YtBJxiiDAJeik75IQPV8uxMJnWkmFVWIi6H8+wpgVpe3Jp6Q4IOVGhVBP++uDKfoqYX74Tw
bMJ3spHx8DaRnIEzAsbP+FSUJu6kV0FH8NqRrmGOslHtf7Vpuqx9kBCY8UR+eTGXvJbw+W+o40iF
2xcs/D3jxgZlGKzp+3FNvuKRDAazA5PsIfAchtBwbIZdYkMPKia52u98MF/PeIHA0wdwW21VGf7s
mBOtbhNXigonHrplKrxEVPFiiyuvMLf4MPaFOrHGNS3JpmN1VBhZ37FiV6zUk7T4ewHrUnzBvNWF
0P7W+J5H/ot9NagSuj3yJdUOoZQRUI0t7TMF2RlxktRWKWjNawKwLC0prtwieMPWSW0pMmhayxvk
DDaql4kh6onIlluLJ1Skc8R4lzGjwkZwueO+GfQyHq07FILe/EL5P0S3OD9o6Brlx/I6EDu4EbTo
DDvn4i5FAOSRdZo0wTisdIl9+M4VLa88Hu4+aDow9V2pEZ5ujyl4Ux2ToY9wNl51/v6yt1HBFDTZ
9aXRyAQdzu/GOAd8lWOuIOOx/G5zwedOxYgGpsYEjyqXSQrW28rp5LwV+R6P0ZJ8qqYlUNijecum
5UGQGRZb/X2iOW0zH1lqD0uuUvN1z7jBV2Ml9vcne2+NmL/YchED/D4y2GxgPHftsySigAPWVg6r
x4rW796HzWwsFUjNnhMeHtqIKLJz0ePvt97jFtzn/npiJ9a2316CxDmrj0O7ww4KrmCYDVN86cYK
oUIP+E0t5znQG98KR0dXFLmTCA4kTMxPDG8qTprIen2ll3u5lHfmSGUpQ9wWeG+xiTWgeW4L+N5h
i5Bq0Xu3dgR8Un5SLbR1YIIYGuE9M0bqQQU6+ui0TpZZvDVI0UDX0MmPgMJDy8qG32HawNwNAae6
fu1CQKwyZpYiRqi4zRLvIs5iMkwIAYMNWXFMp7zxQ1YlbCXLeQvtBV7km54zVZpwyzX4TOzbTEHS
dA00/0aJyeAbepD+5J1Q8zGOkDm7agnQN8A3LM+nPowEKiViIK4kj6lzSnI6Sg+c2JnVhKNScPDA
rKXxfiY7jC/uq51MZuVJbgl7EGSmi1pgJW4PQ4R5S1wR/07DTMHhc+Jn8arrBtNdFydxyrvA40/L
S47QoiFQEf/lE70kWpFhOkWn8evKBrWox4dttZTqJYpq5NTIqOS2xzymdEoT9u3pkZE6Hq2snbAg
tBgBP/tm+FpARqQVITxYpamnlOjFPio11r6yZgNEuSk2J2SYv6FQLW93LSf3BhE/4KjLyHgjmB3x
VsYwEjUv06p48s/azHXnk7bgbyX1SHqxNtf+epz4lcaABlMdZvA4BStoWPOSXIQynScNlNBxNEJW
pnK1Td8CdB0goCC+63y1C13zCxtnB7h/S4beh8QCO/+jX3QuJZFkCfGI5ofVedPwvcpjbQZsR8Nz
Zv9QfJe56bQsBdJjBvg2BuKKS/DKs6BDwqgeFiG+tYKS3MCtf2PAQkOGH6IehWUSW5OMCB1q4PMm
6a2km1sagpH/PAKhglKsxgYOoOuvigQzD0VTWfd56nm6xKw2tZ0vVjwAubV66xndKdQU4xCVvwYz
djK6XmnmtWqPJN2R4MiJ7MS70moIG/KVcFSgnZFIucSw3jqoK7/fVt8ycEFm0ANNm4Jdh7bqYM3L
/sSNtIOrTyjpVgfIjBOCYC6ARy2KGuRLW6LzE8RSQx1uwk1G6eBhzyI5Hi+C85l7EfZ+4xPVcU5d
hszSUm+SaaHDpq1qLerSAySeQSotgBZQXfgyxwk3phX4BgWGPCk9KWyTqbySiE113/b9RJK3RcoO
gVd7tsmod6s1NRIE7eoU/Q0JnDLLbc3R5355Qv3IS0oNSLljNDY4PPjccI6e23zOWmZWnOGm2Gxd
4Kag5Ic9lCy/hknosGOUsHls9WW6zUC4XUnHp2QxHNQHpG4pk2eV9V/gsHdITARecN8wuvmx0HQ8
ZwkEpgEyCsTD5hCK6UB0CbBGXeHcDY8Bh0JykztZp6HHLeiyOOU0ltvx5dolQE/HeR0pMqMUI43B
w8tAbpdM7hsVaUaHq1tJSWfZvOJjWhj/pqHzYH56/JahDyR62/UyKDaN/GmC4BOHtjkBS6ilJJLU
lBRTT14xPHK3ckmK9elOgld+TyUOhDa4CUqhFqQJtAsfKkjWtiTco8tDM88rjL3zs8za3s2XXuij
eZW0DP04q1THGDVcF33stpl2l1pZG/LI+MEaRdWtSJoxAQL+GOIuM0ULAdob/1XvflsSpsVgtqDx
ocWOFvZ771yygI71OvkRUONmorKpQgTnhVi6Q9OWhaGTUwprpTSBRONswB18vCPf/aAC4uadfh+W
dfvG9e9lAkH2lTuJprgCr3E96esOnyG/WZebpj6H8Qdp700qpDPzl1PTwhthYSuZeaU5v9jPestj
1bfhB1BNbMcRcp135l+z+0UeXd6XjWSS8BzrsLejUf9d1LWY9b8cBzmlWKOQwb4HZfBBAjvI3KfE
PNUh48/t5yv4532O10IslHfn1x+EO+59uVPqJajPGUhRpRR+HqhDiK4I6aabhE2cMmdke0B09PQK
iA6iUOhSblzOh5iLnns7ld0OWKlnsd09zFXjeiFpXmyqftlbdpjMYNaYHZqknbq+q3lk/JNzNoHj
o9T7IDqGi/q3oYbfe+4U8vUCBHu5o1+ihLlTUA2KDwyt/ioYpdV7Z9pNUSQ+GXYiHxLPWZ97gc7G
YSHDQ9eYyoCcpkL6XjLq7NnReR+HbURkWF7XooiCd0tkTB0ZSaxMX5RawdWN7Ih7w8fVIMhVuoSm
4DK3NLGsO8IGtXqcqkDQdsflBY/uU2UtBF/svvunScrMYB45OmX0jDT4c433oOtYXMx9wtcQgrUG
MFwsyxs7SRQFxk0RWyRqC+mnYBEwlYGsFHgDE68QMZItDEmIzRh81z1ba+5HUXqpFImzjtB2l2ug
xQbBylfEsJPV/HpxDaoPy0y/F+tB+Dgv0wbkwklERYi7fusFIimQ+veRoewsEhrqunc4u/+ow8HQ
W0MkViySoCGmr/TR59rk7XPGzeqTkmDeV6hiUop0u/t2gkukRzBJ2mBYpGsNvJ1ffKHcP3LXVpoH
KcbDbv9tqUb78IpqUz6FR+M3WUBgMHDObAc13FC4WsOkAGp56N10ez4hFaGZZlhEVl3bNOGGFVeU
wHCTT5NKrkN/yR/zVV3Yitzojd5j7IQ4U81LsBL2LA+qduMnxlFyVKXL642v9Y+nCfw+VLb4HZ0H
ZxAB6H/k0BLUOU9uDbcYCay4uPWEF4kgJEhH+E1v0oNIk0AYxTSZFWCK/F8j6PGU3jaAJbJeMwGd
13vjtmv36Q44BrkWD6DTUkhyTZBuChru7JcbA7fnAp7Z9nVjIo+aS6HlK86OXFYU2UQix42ekK+s
sjLX1+3kfiWzxf9R0jtfYbY2ehiSNgmtyEoSkBagA2gnZCFgzsvabVtQqPWfUx3UqCHOUbKIznW/
cOGQ4oWwHgCK4+ey5DQMLrZSX65z93Yi4SjmO7eZEE982hNEzTiHY2usmeKUVMFOYVq3Dt3w/wua
324PEVoVNmTzUU2JzHbcwa+A7xTQNVFn9RO9N4URMpQAh1QwKyZ0i/N6pgoAQFrTzwqzvYyV3NLW
HcXKzmtZ4EkCmLYbf9Vk3gRDZ4w5m1+WKErlQtfEv+/l2qfIRC3212ZOE6aG3JH+Anl1cvs37DRp
YnyMthbb6EmQNBz0tsAG7Vt2kUhs941SFtIzdsqDgdQSTpjv4otR+ZpVaP6Y1NIOESTNoJ2s/B4L
aPbBg27g5cqsqLBH/7dXuUB8w3F9jkreYjMqaxTvKRu/XZzoqBgpdg3zSh+rlf1dUmt+FNgTmBxJ
1jpxkOV+p5M1JVHlue6IYjHnFQq3eTybpqYUJ562Yc85ik88MoIncYLli2PzzscmVdbxVaeMu62a
iOup4X0meDj+itcSvL3Tr6LWZkvr5iAIT21fdaCZaF+8qTQ3STlRhFF3WCAKzM5lCcno5Q2UV/KU
gjRSZtiGmLkJcejjR6dfVhCxwjn5l0f4D2jA/G1GF2bYWTJXhBqjYlDLIR1IBjPpat75pr/++2KA
uFda8CDfpX/rQSW+RQnCzlXycqPRi6F2FFoyRgQeiyp7oIgJQdbzSyGf7mWbIMQpkZxto+GaBhYB
yCEdYOhAdYokWnRqbHjFUO95WAU6peesLUaVJsydFUBbG2ER0f1aXw0ONgGyUdCtFw9nkWS2aPM8
IDCJEB0hVtGqUY+NTIA/maUAB/5QgeH1c4dvax8vay0jo+z+wICrINVoVxjPCQHecgpgL381ZD6Y
f6CESZn40fsVXRuaOrik7TS7zUvNS/bg7tYL5SpNDRshRtGTNarhvilEDgVZD+5nsx6VPyP0jQ02
xwpqwJlyU0Go6j+QGHDw2ld7aeIVa6XHA05mDQI3k16fisaQp/xilH3FlSiDcYKmyz0bG5N8tOfW
gnMEVpuMQoSgLDRMkTrN8IuX5rB+UhCEgKBjHKsP9qxRE+zTRBsGGHjrfhE4oUO3ww3BnSTqNp+Y
XVmfh2y8Bpd9UJLPtMLhWKBncsLiHwo/y1lMpwZN/vVkej37NV3LoQvJeLPCZFsV6jursToQQdlc
sDsOq1FLuu+58GCDvOxn27CFI14RTVr+sxLv1iLeQIDkAUCBe7+s0Ai80nCLxM3LwQ8ULv9h/XSY
OjpNrgvKmqnPCIeItrOlIlYsOP8DGntB2CBRvD1cBdR7RgV9aIzYCwG7lB95CWvN/TE9Bp9hJxNZ
wGktO2z4SCZGvsSYxgzFcKyZjt/Ef93rYSRis4kP2yciVb3b1PRIYs4RiEvk0G4lIE9Pkz0Ry0Ro
i/6OFY3UpJoQDzKfTzgMK+D0OxJJzGWGSO6+wW4Vz/vi1MLEdqMdJHIGWEMxGYJz4sZQ7fQEjBUZ
Qf9JgWtAmP+Yqh4BIRMk8C6U8EkAyJtfCh0fat9+m6GReDD+Au7eOdfr02ZkQyih6JePR4Vxh840
6Gfd7NAISOkSf0+ohCmG9ptSYERy2mpY0FVw4d8m7wekzhEfw+TlraB8XgLveIFdhQu+5uKGvWIK
EwA+w2/5yWQJexxv1+DpnZM1jHDNnmPuYIsoLFdkxmSQCTAksqxSUqdQSaT3MBuHTr8Gp9am6YGC
3uv1ofx8onTk5lrmMN3s7ionVX1BLKxkoJV8T7lReah8AaWN6bRRoSpf8zYVdJdR9KR4P6bK2DLa
MNV+Fr3L7PA0c+syazcwjxuxZ1jiAOmqgFyokj9iPI51SnUcXmao79WtS9BaWS9VQD532CD5QbAE
qx+O2eu3PpIcJSWdRNH07nUH6LMTULkHoU7F8qCnCsVMOmBOtF5ole1ogKLF+g/nGIhihQdgKt+z
apCwvKAJfobvtR+tqmb1+wZNRFmqJT/M7NO9XvTgC+OShefcCfowImW+Eo4Q4CTt0uD5UiBvd1BZ
29BNKVoPC3Gdm5eBB0DHLV/PPx66tK+ecx/Opff0Dgt2LTo0zGXnz7NFDccYTWoO97Rkww2xaOG9
eO6Y2zvaYTqbX7ZfYuJ3z1qsc1enxjT61Dv7N8D2lO3twnc+VYK1n30bqMgC/mMtXNIR/nb0ubVC
FihcInGEqee21+IAPwNFCtoPB8KhLK4VjJEM8p39w+t5dybx8kJS58v9RYWZv9z05J/soquOaOz2
F2E8JVLD4E6icf5piBK0KkcEMmhWX4UnvgE0rKa2x7w2fa8qHqaMjHRUIPmLB4i4/Af5Aqa45xl4
phhj+sbSFW+PNg3QwwSpFz+fUB+CU1dmB25kAjLQol17/M7ZNjOYPDrtymX7nDOrgWYk9NlahdgH
lY4Dh46v3RE12VBRiD5tQ/7ximmsp4LTv24BXiqArs8clcqhU0cEsiyDmpGM0AXrWcXapeX846R3
9DpQYl3NsFo/sw1ev1pMyUV6fr6r+7d/N54QkGXJLzHhkD9YkPT/OkVzNE/3yd9giC/ci5OQPkes
GbFITiCn/VNuTV8FD81mkF5gaImvioiqWkpXFHS2mVl5KlLfNbo7JjTypH53qYjeQjmLDNQODvL+
uVZn1etso5F3MH4O6+AnMdHEbkSSm0+r6rblolTrZ3Y44ukmMzks/5b0gUIkTJ2XshKTfLUc0zX7
5OVnPD5K4pxKIO+Z7oWs3k7D54+2uzbbQmq5v1O2ZIvuBK2wWxUpMeVQgvxouDV9ibS+4QXF9QXV
Yha7qO8YsY0Z6St0oQXcG2bf7bVCn22QyJOLBUyuYC9vTLPiJb6oi2iewjzRSRy9NB0CSzaU0sK7
bSWVjquEIxtRajHtftQdPHwTJnZc4LBOhXj2S+hez3CRQyfiqXlhqzLkjH4yMN0Z+P5LHkTBlWsF
hiYLD1J9vhWXtwbdX9ptAFU7u5+CeIP6yhIkEg6ZQd5rxfQEdkrCAduWIx+KdxREeFsUOtHqRHyn
5qfXbVeuDUsGvxDEqKW8cOm+FC9j7a+M8LNRpJXHhzCz3+7kjzSybKjzkxzFF5OsOEq9ileJpwte
yWUJdyavOnJFUn9t+9PoBxALasAVGTqk8xGOKNAIHvGwWJ2692LYexCvfmvn38xtJ/CCe6EdRzCn
WQGe4XOerPkuzsk6BK89qDin9Pp8A3IYk02iC1r9P5VWCFENpVWJ714AA+tYJo0WyI9zhlN97J4D
HJCHMOZC+5PbFcFrAyIApbiBxjYq2mOH5omod3MIMLtBF42X04oPR/WeTXhTuw2IUsxOmpfiOSlk
K85wR1pi1iEAcfB0oM3MABpeqZqTxb2s/psu2K7CRGto7wO5fW3PZ9e8rZmPmEjom00x0ICOmlv/
8G6I4RfbQ6acL6xPqsA0cE9cjI0iVnnZIA60LHd/KDFtkNdph9LChu9yG8cyQQK2ccUBrgp/Bo/f
8Z6W+Tm+gdTTYoke9UooZxSdjHesnqL42fuvKNc80Ee58wNr//IhxoijWqjW/5AGitWbVYV6Rdpl
1vMrJehrLCBEjNcjlzID8cgZlmGdorXq6u/55hO0VQkjbxv/P5uSDejKry+ZDwLHCS4N+Ng34TJd
TF00lmEXKRMH6vQzgaDE9+fioWAPEBG/YkwKNwvf0F3JsTO+H9PAdvwklS1/piguNi7wkGrLfbDr
hBvaHbEHKkFs6uCjTjiuBiqj4EyQ5ukDhEmiOJ3xUOxaIT5XVNxRpVdox2kF5DIM9WqKXhFzY++H
axY3nq7gU31rY6gV8Q7yLkN3NV94H7ZtHps3P9cTSQZT22oENSTMA6YIcD9o942QIvkq87tisEAT
HC6n8eHPj/6ONLOGpvVccZs/v+t3gHI/8ZOQd/+9cOQcMzXtpvC/iY9J6vm+dnm7C3bz6QSe78Xv
ejelcUgborqF/lx/9bqdvNHElVOH5xsw90iCKnRieiI+strWUDAwnsLFngKR+W9+BBu6lqL4U6Rk
ph+k1LcU7KxYAx8auP752t/x6Tezi0qqXPuAIT0Ng6hk24//NQx7uUGN3itJ3Z69GZlak5g6UGt1
/B0TWr/jMbATQgSJWb3nMqUlIhnQpTQAz4MXG/03bFXNObcHOKfK4trKo0jPXFYi5bT1lXVZrp2g
RgJFvyLOvEPh1IAJxx+v8UY6aqhinos8QJQ4QxdD1+dnlahQzAayfdow68UbFXcBqQmZfRaCVdfr
VvnbTw5iKmPaTGwX/yTtDn4bj89s1stO9L1Fb+3Q9FrZxT/f3h5sjxspn2gAJ/nyFWUWdS3d017T
ON/k9A+R0QirC2fBhFmIMkvETswQ3nYy06j+RpyqfF0vW7KpbPyfgN35w0ndrPcQ8acGtEdqWW/R
5LJN1/OOeMGLilhOqcn21yFRjaEqXLlB/plbxFISeDTrlohfbnde1dGR8u045Fk44AM1f6UAOWWf
p720WODSF/5GKbXcHy6Skt2oHDphVPAnJ5sXwipnEQKMOhueh+ESjXOIFelfasCWLZLUqz+ZGMr3
u7PURbMb0DFzthQMaTBiAhPN+FUm4rEU+GzwHgjdtGqUaKV/ioNinrSYfd8GSMemOII0xMVLCAq/
Ltx7T7SxXcqTFPNyqFXup7Hb9ftMK8DLrKYpyI4NoPR2MhFpGomQAFnuCa20YDfuGLWDfHJURB/B
7qAUiO/i78oUlhHC0lX27XsRXJa1byKQp/tpKRI2hDNaUcnaMrt2dIjVaJfVKxx5JD2A356eDx0S
96rfuZvnLq/VoAoZhCENXmfNbP5nS7rN+PxcUaCJ2YcaMtbWBMvDXjlMcm2Ao3GmnLMj0LkfTZa7
OsIc18R8ELvt+6yPXJJJURj4JmmvI6HB0KDBS8+0wZjIee0LXSR2LTlk3XTeGITSnW/OHYXeV4vB
c8Jz3Zwz0bYi0ao/ba5kFS4gLNCXbAnbuu23H9rVMVW9YwyaVl7bMCGnBRhBTGyo+2fmcAVUVaZW
9pFWTERTzHnaJbA9+gq+Fna8RFjxTgWOPJgHiGer0OSTMQneYIQvkjmWUrK6tOVOjGswJ7MSnKCD
YgIcoDvm3IJvzrz4KdkEomM+VsOYjFxFbowbJebt7ZNSk4FVvYB+JLQsrKlS53ePKkUwe/TDErqE
qtCvUwoGvL9D1pyPEYJLVJ9EQ2fg7Fa3shtUA8XDduFqyahm/tYI4taot3PVb3MHceuEz4gnSFu+
wPc72YHra0zzwjbKKiGZw4aGwMGl9ZfTne3sfUBgo9aCO8agV1pjlthqg7yVeEmMqsYj8sYEnuVO
m2D6Dt5ezbB3Xb49wismuhf6wOBQhJm8wIGQr80xthmvKIfedR8TfeojgSOQuNlEH9NglEisPyS3
+0cF69frJ6QfmIDjzBUwko//e9HRjH8UU9+sfEdJz5xkyVcjzc8WKO7Cg0YX5im07BSdUM8vZzXh
0a2sYEKVzLVWUclFbXk0WII/uhfGlKIudknQF6An0Q9DcrC6wAya+mSofnhNfjFEPCrs6aOo+qy6
9l+lW73AZ7IamNl4Sz4O/9Vh7t0v4KbRG8bpNY4Pudt3iS56lVgKfNUzgfUFBeNOk/0LTEZXiKlo
XY3bDQXSJdJsPr94pkpPXln3R5Uk+fcCvukf3g3vSUAeBBysZrxkAr/ZGKoNXlHYIYBqPqEX7A5x
iTJbpg6CfLGpGgbmMhnX0V2Jm4suIVbdF8ySecWX/2C3SFQ9LSiB4Id3Pwn8Vs9pKZG98hjYMCrb
f+vnL3EGD6PhNoF74vQ0y8CjXv17/hUR6BkWpK4k/8TS0WQ3tfjTTsrl892maJylptm7aPryU3d1
C0lnTTPlvavCxFq4n+CpPWbLIqFHjoJUS5KJveerHa2XvMP4Qx2dBPKsVr5xqEwfkUge3gIONz75
J5UK0CGJk2g5cqU9lBfOxwZ9QUCCxLwByeFX6JSTP5iBztgwuCPP0dA47E2RHjSmI5ISdDOTtx7Q
6YsA2qn0wenF7iHiH6EH20aqL31MsjXKnJJPfsfdVPfARPfbUwb3MHz0VQ1tOLK7FTSDYwO5Gp9i
XvZyQUYNMz57+2vJrpjEWkGFW/ai3m/jIrKYSbmKzVLslYKO3e1tAPUvZl3gAY/y+DjeINsFDKVw
H56Bf7Mp0mdw7B0JM1gFE0XbMJR7DTiVKHX9Wcs7v07aZZuzo30vmRns7kFHY0iOqVIQKmbtlhfK
iLMQeRB5/CTP5bENM457qFT3z/WR7nRV+KCKPTn+uigmWq9s2ul1vGZuQm7jaXBdlpy9vDULCft6
KtguqtGUGx8LEGusfva2oDkK1W1zfZPkWzIDxipG0jgywNsPXJodHYuJVVSrLu86BQSIhpiHeMbg
RmheRYvLwCo4l965blajXA3zgdfAEGYvFt67MmPoTKeugg6i9tpHZzIeHFEa2VN/5iviPyVbw+Uh
OB6YEe3bDTTTaC30xrWSIBWubMOa6E46qbUwzqaT9U72MY1LzmA9oyOpfnCl0x59T95Lg4hlm7BP
6+AKsNPyAVDKytiFzjTZmNiamtuUrKorz3DWape38X9FICgo0DVG8Fyvpz3tsMbNaszNsNw8EnGm
AkxpZDWe67sVeup4J4EaFHmW6bHcU0M701tIUB/b14Rht8XJdSuGfZ4t34oSBtyaTroE70nvY85d
BP23UGVWUyh6XuZIru9nKK8zSACpnP0ReKo+P0tI3LXkiiWlUFAqHnxCHFxsBBW48vAEwj8ethR3
H1rD0TXQnhmqzti8ygF4mt9/qKZzt3a0knOORdpWfEaB7y3vwo7R/6H671s/yetbbMszKlbQtfr8
Uzt+p8fdssKobJVvBaLqEpZuPv4mgs2YmoqjlAYcERzGLPKsba0jGH7iVeuppl2hVjOTYLRFldhf
YjQddXP4s7WWVV3ek0IMD03jmSKj5Fqp/V1s+2/uwuLP4Fcvwz69ehdri+zN/h63XAYvrT/8AHfY
vpqwyRBEE1dcWwc6/5VOXXILm5YoZWBgrD3S9ziZvxHxa00yhFfafnJdbIIH6SARshnlvr7eIjK4
ut7WUBvBaZPBl8B5lJaIgOxt6UtBlNViweuBo5CZp7rykDkQaHY0+tCEGVYbh6kyM78gydgSQBx9
HwyJ7f2lhb1Z6qVzIm8EECyP2JWuEE9iCylgqKshZLBDJg+nks62Q/UrBq9AmGgUIqHoOl7rCdBo
Urh72urIU0v7s6mVLZ0ORpBMsooDT4VjNZupBTLqttCfirHx+Y0Wf2RU3Na6AVhDQVt/tWQMa2is
oCjsbwwmjzpuFHFxL0bR3zBPpBjKK/OcbYebFIEh42z8HsZi8OeyO6H+nhEu5/4dKhj/vafhVrPG
QNukeQ8gWJJJjG0zF4NLhlFvvjrZw90hSTQjtCaIyNhjRED+oztdngLhAXplyE7yO+78a+8cFK8h
+hKj6Xs6JlZvvcIl4pfFZnyQ39JO4JbLLMwRjJcFa3Ol7Dl5v8nL4uTfs/4QM/XYDhLEkcSlfaVu
QXRBZRwjCIHwwUbiDwDmH4c3MmCBsT6/f3BK95Rt95uc4oNY7r/Sk6tfxBO4IQWOQGKicEMttVFY
frjcUwzZ8eiWmWDvyWo40gMgdjBmwAxcDH1GB4pfiLJaJscbbtXvYRgM1rhtg1wCUgaFYIFfs+6L
vhbX34xY12CJ1jWU0LxYHK8D2b1UsraEhH2g4dHDOPNurAe69ug0uisWyeTZZf2COA4Ug9QuCdv4
07nJBnYPkBC3PkaqMCXKAlcUgczhFV+Q6dRXSNsHXxl2FbR68NyRUCjROd6tYvb1b5VLV/zUnoEo
MUpstZjk/z+hzOc7t35DNQm6YjbU38MWIkY4rC5DlESJMvfGkndKkc5XBagNIesKfvKu86vRkA6+
TSroetSudBTj+gct6ukMUlJq1Zxed8cR4sfj7xC/tUyGzEezuE5cmYoLRfAKDvoSGBvFcHLDidb1
V1W0IWx1QwobvkHzyrTfNH5Vtl6KH9vGIp8mfBcaiDsmYJHqDTkY1f79l6md7onXWe99vLcDLkfN
zz2KZhLRg1Jzzgi/cL0m8UeSi0ERJJbQ4q//K10F1sMsBmNbSVAQLRNKiAFeDw4+0UsmmfQ7gwzV
aT+buVBITyZmztlqhrPBLXstAV5DbGnV+pSBmQUSVme081U5VBjGjv8ZVX8QElyY2LQGOXBCi0Uu
SmXpovT7ICKK2KYp2REKhNMRbHI6eTdDSlC+EHDTsP3cW7byXcZWnG3LdJoe5G0lRCK/e6Gzq6qp
Pqwjes1fxYceS7yfQi1sZvhdlotKyCwqilsYq4k38B41Uo7MzhB+vgEh7JLACv9xq5qJEIDUk2fx
GJ3ldYC1mAzsf4e3WWqOncXO+9cLX+Th0KWp9Jqq/YcdUezjga0YGfK/crHRQFuBh99SJpHZThUt
ZpqAhgLYRnn+JlgW/ryvuOmNlFNdGp0I0IpS3dDjYJb+RQvrOWwZA9aLUClYaJPGOxEbdtiuUsWg
xR8gxNo8YKEiLhQyeVmQp6ToXl1XjB4cxvFlWXu42249o/9CngzW2j2althkx65u4KOAJa7af+R0
CSNZR2LRhjQCp857ktXcRLpBVLSo19s8QxixRns2By4Qw3TczDkaArOUtvGWj+W9RpzDTwh8XldV
iXd2olyzOyZ1LZLhREgKfayAnxkRAjSwu/NS2Kkjzpgd/txhdg5IpbPK8BgvgbC+XjhcD1pSEZAk
yMpDP13tlwDWPD/EcOGXcpVnxWpkAqsZMtBNE67p4jNZ3B/ryWsRS7P+kabn5bM/yL6JPgpjX6ln
416eN+xVhGti9GkTb0fCk5H4T5i5sy8Yf0VVPANuuvZJCZuls6N7kn8YiVCgms8RNFcAWwvT0mxj
ME7QV75ZZ0R2Iy0JyEx9tcKu0ovQLZsXz7ejPPJFA9tjXY77QAhUcmtH4Mwduhpu9/zMklIgJZT5
VY01MMo+naouoIkPlF16vSoYXaIzFpvUXQgMWgflRKZP5GvdHtVlCZ5SGq0torPPxE17AVLhsL8a
Meua56de3ehhTxfyf/kFY03z0OXJBQCadu7NeUuLn4cTKH7IIbXyepOzMF/GxK8Hl+ggpp+oT7xA
8Jvk5VWhYU/vkdRHXpmBcfI6UwIjhtYVhIT2AJaYf7F83E+cMquDpFKpjun0Tn9BIQNvd2EJ7NCG
kemiJhI6f75AA4TiEcT1/v+C10c7wXycSD5mE3z6GQD/iX0Uo/je50v1S6uO2jzv0A+BJEXgUuzG
jIrFTv4wSmYRrH+/j5fEGz+edKLbs4J5I38TN2zI2eGdDEQInCkYWUMmBk8xahb310sQLFB7AzbJ
dRYyhXgxHWINoHNKNmLGiHwSQKNOSoeFUSeCl1gZhVDVbGa5sdE6DGH622HTmcCP33IgpFi8Lwvm
eIlamVIwm+mxRNXdPcC9/L2axFkCq0GAGpx7KWdbvyAt/XRxgzOCvurRqQ5UZ5hkBWBCNr2pOy8o
B52rCsNVFGPK6Ez3i0jCV526fal9LTViogBr7BBEKKSDEYBhpDLzezrtQPT14pJDBX4vcbKTUNos
gd0F1Gl0Jf788EapGzL69q+/2QWfWf11wVK5+HlBUS+7fHjjnq7uXYPtqd+A3k6omj/XhWKE4OrS
9EHEIArEdJk5y73cr/Zy6KGP+Sk5qupeuwUdIc5s1Lk6Q4eqr8EG/KBA1vQed4zR9likeS6Gf77w
b3qAlP7t1R3V5hvBxUuSUiJM6HcE8yhQOaqIk77RS7bSKBH7bIg5lWx9zo8SBcB7m2x5ZrukORZn
KQ5ZhmDFmAH6O1tFT19KGUOGBrVsIbCphWRM8/QJJTK538IwsUbNF1M9L8g0hu9dxG5U0doNYOgY
oXNJSd8gy5RyfbDSf7v2vex3z9unZtSh9dGORQAS7o6TdwZCmbZHHSLx/6kaC5QrgLDBCGO5FFlL
+aJhre9JawjJzeqkvQfY24wEfg0rwd/iQIR7ABAwC0C14cgB8j7E49NZpQLwf3h+nmJxlWsPf+Jz
fWj4HikYDbl/KDxgJPDpLW/+SC9LhyrOSRUqL7pm7NHIz7cBnFCgcjdwLRrIDFNpDRiMH6Feb2M4
U5W2cyXv498tu4q1aBHp3nQCUBj2LWDns+K2f6UlNJS65qZFtKG3gJ+Xkz8QHV24WID182yQtMCL
HmCm7BWuLRlw9rUZbaOKF9hTEJG5Ly3W+vAIH61UPvUd+rFkpEfXtve5gGXRcnh9U2SwW7G+nRHP
ZmBWCdgVVSoQe1BjgD9wUapU/gIzOApoQtnTnsKPkwVUuWbxWxZJAuihPqeNfy2G8+PfmZTVtySr
8CRDQJ1nWet+N3xQzf5nTMLOC227wOqbcW+GXf0CG6BDPcOY1fE+bvlUG/1P4xQbofstHr6SXlgQ
fLmrKxgfGVQbq+eDw2S+3ZM0n2To/jts96h+066mhWF6JEtUYxPR3B+nYwGXxoh12F5IxClfUq1X
D711v5N0ZncYDDLOWhmm9bqxwxNVOWjL8VTRnTppfOo3G0V6n5mtW3+BQaImvdN7ibn0LgoeFIas
l7+tvXarZFEz9jy8qsLsD0umeZi9QRX1ANj7xO4a9lTuXXNb1NcUN+ZBZKt7VpyIxMCHGBoHmFBd
LRv8crAD5LHaojIVK0XICJEFLBlqcoS35ie/WlnjHXAsGC3JZJ26h3KhNtI8FSYp9aycJg3jN8qb
2O0IV0NYkOx6PbjNm4G/aeM+K/S6F1DcYw8neaQF3mdQJR6a1Sw5r6kArK7gksBGjZBl/JFAb5Bm
JrAHVkBMxFRkPEv9FFsHqQVYaEk6OzT2LbAYthl/VqQxpbWwb6XU9LNzwzXYPqzWgq9DkMGGfnG2
EoF0NYBGE7NrK9ax5jaeL7Z60RY3WWW1Gh5Zw5GwRfaiF9seZaEWIbEFzfzGXIjmxw4MF9qb1J9H
NyXD85nioA4UMOPBoYyE/3zi1JqIOtzFyFa49dD23AtaeaX2ycP1rxrtwdKwHR5BUsk7QQt3zgHG
yDzqF7bof4zMgMnGEocwDg+5HewHe+mzylAskPAawE9yQLN0vgZqtBwT7OsXTP/T6BEc2kgoKLNR
pHev+CNKQcFni6iwleSbpCZgyHYeNS4HqjRJDGYVffR3eimjQNWumM521K0J2pZtO3RNanZXfXL2
rs4CmBg0wLJWGKxNnFtPuN3WWCGJSwN9NRQDIwGL4iRmso2LBsrdAnYVKDml/7VU+7/wnb7EtCVh
ppWsdQD3x+DWE6GBE5N35p9M3plmed9/5I7YA7FxKFugufq1wNGHm2WOXBaOOFcD/k1zgsFc58ts
DyCSJKAHsr9F1wmJvYneRLX0XK4LzbH/ctgUqnfmLAJP8o6YtwkzI1P8EW7nLkNSCKrHZQyD9jLl
WWES27eZUQ58HYKROti7WfPk70+Fq7lynZnNcnKJJj77sSGPwtkXQ+aEITgrgJbkTbTV9ZwdAvCt
S/ooz+HkVADcPjIGBNpKqzHLcGN+KhXqQI0mcPkgyP+fU2Xez1oc+OKkpvKcFiTsbHiTxYPawNIS
6YiqtS3+3MVfwDBHWHEBSH5vKXXYGwBSnNVuibazcYgpKCmlWaAZIoHdrVWYWDm50QkLK5bbp1cP
zm2FO/gQpB/Eey8mItrEMRwBNteAgLCDU+A5SJH8qpIVkuS57SddyFMTmy87tbSb+PGfTK2EIL4Y
yhtYJVmcTYpY0PZPKVa0qMTBexS/8YFgnZEWkWNYf7BBmKbXfANXQHLOYvhpg8u/fKHRac2VwyYx
9AsvRcPE0i3VoaSXLDBKL/srd4a7YhlhelzDrK0L/TWN8yimgBB3cRk8lgqoUzLR/B6HsswkOn40
7wG3ciguhQTfKooGGC/+HWVfShECrvCfxdCNZpjPlQe4dsk3FX0xhLCbz2Gt7UcToDLUQ8W9Wy17
Fsl4fVMHKf3OSp+0A0r2x39Jr5928Aogx62SLbEps+fuWEWPDUMaFiGCyJLG3vUJeJVmoMeHPyxM
hxV4/lghH8JNr8nFKUMF2WaqiH2k8gRS3kV5V4FGwon4Qlkp404TJMZEdnYdm6/FYngLfqA/GwL3
27JYDrYbmKHDq50VtqbuczAhQXH0G+Yyxc6v1n9+1vv1M6ezJGaIOIYuP1UlSCfvb5V31i0jOjar
RYr+V6mJd6sfvn/Jz+nn0iGKQlB8MtDz0gUbk/cEZAF5uR7FWTU5LN45myPlau0VL5fqlgO6JvM9
tYvZcaOrIB1YF9LiA4ti5KxM28vH2lc+ND+3h4T6uFlF+kT05B+CTreoeN1c0X1eE3CekybdRJq1
+g4MjdivWbQs+/1zUxQ4XF9/jAxXiBChiGYDzS9PfMDxiUHhK8+A9MrD5Fw11DnXFxOYe1o7lru+
anvXENFd9/WbAmz44jcPnxy5q5+LoRq/w/UCtH1PsDha0guEOlWApYsm5Z4eMPuLZ3VWgyqkwza7
waeBKzCT1wbMoWudP8JuNiWxsh9Jnb4oVVC2S8nMWRJy40ua3JFaVcz+DL0s2DF4fMW3TM7DsDzf
a4WOzGLTVFu5qZ3QdGYA4nbMakmVImjGIwwhEVX0Mvpz1pdR817MCqixA3rFBFkrXckqmAgzI0Kn
BZ9ne7oHShYOco+ZmlG5zisvbFFG1JmjoZrZP+YSwvWu7917EW5PgTu8BNFq+eKDSIW93hi+xXUv
ip8pDZYtUdaOGsXB221ltIxf9yErlZ3T2DZmrbbZMeZSHCAOObbAcSXWeR4Zxad/g0IMSuln9q+x
4kOwZVLrXQpCWFz2sq52MMT6l0bunESZ0UKWNW83mpkmPq1NqY/MulFWnbg+d7Xb9vkmc0mVNF7X
j1Zmni7lsj0P1p3k20sb9B0RbKGJ+X3revGklkcRo7mnqQWxAvGLMMh4416bB2kv5VWV9HErAqyu
XZ/IsWbKC7GBfnn60u+3yDJDbAhrj0qRuT2cKLvEMwu44WzsRyxC9syQKoANeEtNLFbRnhjTHYwg
qZazND78jR22MQDEzgmz/3utKQNzyfrN9/5why1VMzjjb6DuPjabJ70yXVG4dYNSdV1S6/NEj27Y
QjdX/O1jSxndb+R1eH6i7PBQvPdO9dvumtanatcb5EXk+Up/RM8JXRcCAinxCL/wE1ObzpbeVulE
0LDNVH0ys810OYUt10saZWyQdP4PZvsVGbdz6DrEgazVk7tI67n71N/0xLzsZhzVL9g78DgWiYto
R/ixej/6uPx3gZ35FJx07Rh3GC8IBnl6CyXOgVct9JAWL9eTGj0DUTJ4BaAB692BQo8qvujd2Hhl
z9/LIu12C9YdGJoCqa4YKcX01BZFQeS4uVAQc519OkK3K6RxezEQyIOU/HtncIeOAce9l+jx9zV+
Ik+3kaC6q5wwmxsVU+4NXG7aoje2o2ukVmmH2WNW/ChrMIZrXsWx70HvpzivuJiKDNep9+0gDMpI
GvDcuBW7xS6yXG0K7noprn78XRgkUeXoZGRFSSKiu5WVfHza+l2p1dsT2q1XC4sQPXnG+mGiCBT9
eo9LGhh9l1tbhT9XQjbaK4R/4nxYsk1T+9T8g50JNfyenUjYZNTxVZTL+VkSFPiRgGi6F308xCJB
futIuMXeV0Ehuh7pn9ceaZLG3BzG2/0/+83eb0q6eUuP6Ln8HXuAsMwnti9wzIi46zgHni+bv67C
pz4vadGgb66dSg4W52W19CuEKp4MKlTsK2iPJjAUOrFJR5pWTsLxUakICaDWjrP0jMOgaahtSu34
PkxrA+EUQlTqd5WerfUjcv7VcnwGxN5N7CSJQJ1Jh0WZ2Ea3RNckjgkw51Mg8omvSo7xbnu6Z0vV
HuhvEaq1q7l1GIpg40Aus9Ny3MGVfDiC5L1C7ZmKJnRiEVfavBh7MVaza+eaSHNObvzqadFmRav7
RWa9XMxSZZj4bsa5fWMP+UAecx0CSA3ixIQS6+falF3ZC00WvfahRodNcg/5ASqyN+oq+8jOiLwi
77GOUW50BAbwldrmfdooEaZt+uhlbk1Ocbj0kVtEmG/684xg3BS2L1Lc7OYJ2yhrdfTGZVtIcT2a
x22SQGEr5injBd3nm6T7wb8iHB0zqPuhav80LcLybBGwI0N0nGEZqmqgqX3dk9FbF5sQ5ckbp9f2
18SnuFyCenwEqh4uqNsQQrJnaVGMIci3nx+pJx1Xd5AuYk13cRPaE45B2v/re3lxG8Mu94bX/H7o
72MjFpdzSjp8lTy8Yn7AWZL+RIgeUmcyfzLqYGAfhwHbs0zBe64Ugx0QGt25Wapp0i0TzujBdXaW
uSo/WUgLgxsvl6Gr/1w17Y1Ap8kC78/URI+gwi/uXexsyN59iYqpX76sW7bkPABDHGXd4FkIc38d
/CuNPcZD8CYLzxjY/Rr5JycSz6ZRolsv92e+RMo5cNscLiL9xbOxqfn/8wgQIIJQCZMTlTCLYCk5
8xH8vbPm29wI3dACx38qdtLmsSvh2K4oDnaZ+LYSNhX+Y+bjpqlrFxy8FgWnTXRWWO2LBg8si2dC
4Q/2MuFZsJ9gIKcvDpBeiqhp74GfNDsgPdJUrmt2Ewcy2dQMVl4Qunt2e4pwGBDeYzl5HG850z6M
gtMavrrR6bvRYCgaxTKGKGgVLaGSCkOuKCZI0TBp41NzQaBzhoFHy5xSYoNYUQ5mvdawyAGWBttP
9yP/jK6X9hCRCuuZw+OUF5bVi9fQ5zhT8qgUMThiIJun+bjZeq8ni0D1yZy7TVc4ltlxP3AW7jLk
NkZ7RVUIhGhr0dGbhHW52fLBLWrTxVuwJCfsel7xffmAI50IpOKAjuaA5euqaUTuXm9tjKl6Hn82
Jee6fZRzotqyYJrQyv6i3IKdsMBNE/bgaVEvTkZQ/S2arPqw7JNfE3JFUFWbLcoPioLgvOhRTyVA
++lGkheEcNxh+ecSx7zm1r0JVRbwogC9XcCSDnKKl+t69mQq13SkRN0c3xQk5AY6ga/lK3Akn7w2
zt3v11T1WE+mZgHNKw8To0EOAgbqbWaFE9zdUflESm5LaoRmv2cwhAkwHiXNYnHssc104fpjlquZ
yB2xWfjyvrEhaoKtxo0kU3nyWAihByTzxsDUIBRCzm8Z0yETQlM9u8Zvgt6MxVYk+/pa+Lx50MD8
4lEizuhEcwEL0RNnk+JgMtaHu3q7BiLNRnKbYNqpZ2qWdJFOdiAMBRt057ENx2I/tblnSZAj+KTJ
gmU6TAkEpd7/yeAvQjJHpyKTaL6PwnPeTP+a3wixteBwp9p9/VBImJCpJkGcMGnpaDz1lMFI2Vsi
6gbDlpNnnJh/cWcGaMWTFijuhJR6JFGxp/sht42dkfk+FxoI+sg+wbltzgikfZSMcROUCBltCRFI
RIzhUGimYWGr4kohQ6C5nvUVJPuuEKAayRG4fIAZ4L7vmcpGzNQ06vJt+wihmxUNodbMrJ5fwV6g
pq+JGm1t5Vsm4Gg3Sct3bSSrjI7TM8ojqHuiihKU09GeuTDdyKnVWvTdQqUmH2WaaUMEeRhtMkkT
1hNsqU/2UM3G0lk8LMQzyC2UuvqPi8Xw84AKCMdlZPbqeQhFJL1EkVfvCm0DGfvSW1E1Qspt2sW+
b1Qubf+Uy7dpaLnvVkn0bPclpNq8B8QaPE10m2Mm2xKLpa0D0melpvrMKMUg/oZ6QXaknnan0oFB
yDXoZh+kQbzR0rh190kQ4bra3kFaKEsVI//RPwf0PuQKZz3qrijkGNGheJ23DsL9+wOuvZsrh8UT
kL0b83OG32DKJvnLiuuIF9z9VnWUct6o4kMPbcqQ7m/TGnohsoZfxM2RCawTXX4rVNtlXY0Xq/Id
jSH72Aiv8lJ0CfP7mVQCJTU+BLELQJckUMFNj6henYeUeUzWTzQgskfN4e2VryGUqTq67ZK0yZys
6mjdlaJJ7yKp1hQQeeW3eVFmolj4cYKToAW8JljWuIK5J/02A07JLCBLVm8eqzj0m7Q18dwda1+p
OnqzT6gnZPbVxKRyALH3L5gkQ3dT7FR8RyHj3tRkCSINhifRNtT/Hr4eAyL/PKGUr11mMsKga+/r
3idK6pIzuBpCEFoBkiKOjmJoqxuSFEjUj74AUMhMTzN1T2OW2oeeeP72tu/tVyBGrsFs15C6Wl9G
PYZT3UoJq+Ukh3oDfAAh0WPhM9owxRMY1C3GPHUSN9oLugiJT3VAiKXXoeHtl8Qzmpv03mRPcjz3
RkEuFQcRzTs6I6DgSmU7Lnp1M+rB4LKLnouzLO4cClZuoUrxGf0vMJpbIBK8p1D+gKZzSCBtdBSp
RxXSGQsCwfL+Nn0lhH54CeKcU1Qz/ewyMrX3qxAASRg5z3qH8GnE1V5aTsJQqsHOuZSt2R8Hsobr
PJpSZR4TyugAXyUlNtcFxBMD07cl5G1r+q8BY/PuXNV1/3J6f3V30/msgd0C8iJXIProf1REwMiX
pFWv5ftG96/yr1Ld24WULNtcdj3CnpSwEGiQx/SyV2uaVN7zPaLt6fl4LSgzaQ4YzyT3tdPn0TV2
5m7XvfMMatfWEzsE7vV+EkcUb+Ch9ogKqEBYeyoxtLVVxJqboys/b4AlWdRHESJA5MavA0hx8h/i
/DneY9eExXikK6kC/RskAm1qLbomrSgmiAQ5GzmxdVX6qzuE0R4VrNzJPxs7QAjF9LUvDyJMAdzI
GiDE6v0Tbo8ZyvW3Xy5ZuxDZB0erKP2ukY9Q0bqwUcmNCB324ax1eKj35Qr8ONq1gJ0F9bch3dLC
Xq4kLKB/dJZU5dbnP00+E1rgRVUf06Uk5mpFe9+pkmQb04eaPMpowo6WwQaGpkFokO3fNk54/hcI
XyEJKHmU2mxtBJOS9faBqg+MTYzRCEPcNIdBgpDW2UB7IoGHO/pmkbcxm1nG55/WLxP6Zhouv4mi
/QCtHNQk/2k0d+uPHugr9YNpR12W1EaKWT4S5CV3V2kMAR9KxO1h/OLBetwQev2nYEChBGguQNoz
Vr7oHK0QU9Zs1gzUTBcmCtT0m4yDduyVof8Ejo6PYc2jzhzz8otngB3VvOPr8l1hDQaQjJVwaBsV
SbiVMCMy7wizqkMZI8gcp1WUAPMNtpazop9Ql97NAQ+QsshG/CVAMhOGhOLCsoDnSLpAz2dvc3Q5
GNOC9deOr6A6jjnowAYpilCj1K1RrjbS3zjtHSho8SjUYC5YVnUIEX5hLOwXkLMWfVIeFgptKIPx
WA9IeuZ26kY2jBKUEHWqjzTQ11mQBjIXAWQPx3+IwPAuavOuYgrZBrFBcNfp121q+e4A9UTdFNwX
i6Vd2gHVTECMIfvjZtGiOljZ5nQJl0cmokh06gWkbggH5iys7Dd+T+lz11EKorxK8TbsVDPdVZSw
etOgb/mOHx90J6AAIWcNkQV/GY8Rpp4pejIVP2e6Bey9ANap+wE90dAtxGrtOzp5ugrC65CN1pzf
hxmlf1LvVluPlyVkX3GsXpZQ9NJaifhAYSrfopRAzcwG/jYegeByKZlvmU0VBR5L+hTlFxE/modO
1JrUFxiEzUZQPtTQQ8omqQ0J27rcqOd2TdDR0VDGTFl9EgS4hb4PbjGq3AN6fJNTzlAt9zQ7V2kG
fBUSHSCSDNFDZdmSQo+Vq+b0vsuLpwnllX6naMG+vhwombuQgEspO/wwpTBMStng0hucuapICKV2
szjs9Y3dodud9b05nZzDy+2cwDgSQ5cPI6VFdnKhB0RuxEbF2cVWH4Ojch11Uh5ddxGD16cpRNBW
RUvK9u+Nq9OoXZexFjJ2OhC5p7cdIYTimyqQtEwY2j6aAWqXhXB/c8FN4zhMxwyMos/PY3zisgir
h7uaJuM6CCdUzHFcLYkKujcmarVn0S5xRd3221oxkADDRFlBXrYMutxHso/8wZNYPTy2PFoDIgYu
KRpvhRsxPzcvEEpJ6tdvotdIb7ohmoqubT/Kc30PtEdnsM591OiDJFLbP7A+D2jOr7vkNrPDf1Nz
hSTxAhzyaka9OL5nezteuQtryszAWqwDs0ZQEE68fGgqy9XJd9YWzRJIFCxkWdz465BqgJtBtRe/
73UeE+rs5gpSUl4vtCUAwGUnAKloNILRX1IpHKjX9CukVQA0sKgU6Fvbiej6iSu549xtu//bkrp+
ef/fNcGa6SuI+kw4TMqTFOziaqfSAlk3TshLMja8r4Ie55ntcwNXYVR3hCUgo86Fue6tHSQSydAS
MiDCwvjUbU+PZI+8FQtg4W0clgxFAEcG9V9ZvpkEk1GC1zor85EPhy/Cgu11Bwqn9lr8QQs+raVN
DPaksxD+i8ZOE64QtZ+sI6oqozy/tWxfKSJ5p9ElZiUcUAXAl/qJWktKzUos+6LC7z7l9CbaFl8n
AYUc6hCFCbuH6SEBk/3/kvd4QqWarUmMH1MkCJIJk8fjp0w6UuzYX81II9m/57viy7/VGtkfO5wd
iw/wE+XgHioQgEX0zyO204ljhfou8z+JS721eMRIlzB5dg7QozGvd2mwiPHklTDSrbH4i3YQOcDn
0ipMisQJhQMmYZ8vRtIsHF0gUatUstgfMrJ6XscAkod/bQSCr8XOJXZZabXIBjo/IJL+Ok72GWxF
SAP/aMDn++OZVShlX1eQbtv+p4OZfMO/XKeqr/4m/dT3XKaa9AJ8D2dgdDSwKzX74vtVeadCz85N
Zh0wijzTYQS3wA8aoIRMxqfadCd8UCEkuh04w2d0yVqocuKMVxyNLAcxIXAE3ChQOLg7J6ptKfC9
SA/xdjSPgU9qXpCWTGEC5b7zm3DisVBhXzlQgiAx/n20cz4o1irl4kaBllHgW0IvUmdVfn5Pt2V7
sR5hDWot8AtSxLf2SGVm1xq8XiIp/NK9o4ml2oRNSZjhCFJ1JAYIR5lxZwBsDaLF0n7HUh8ikPhT
rK/FXkmNeHLHV3s0Idv5fzbF2USX9qLjn/AeUPJyV2tNuYemXRb5JeZIu7uDeVWIf3TOEqaktSoc
nuCiREp7pZ3tbNpaWWgVWpBDajDQVySVvGclb+cGNhcWcSZ4Sj9tKVgisfXsZHkeAZW76mcVoTgD
p8H3EjmXTuZ3ugu40nrr66dqmY/cWt4HD7wH5+qb3/FyfFW93QPvbAHzGaXuuIms9ph0Jq9KaKWX
/6n4kL7Y8yVBUHh11SwQFBLhjVV+53qWoXmxTof60zrafOik9omSGGKUhNsrxhpvywpHlnKrQyRF
RWMN0vZkZ+7HK0kNirJ1rzYmq1VnCAVArIgD6uPUaRtRcjObTJAacSFe0ke3mKjCFfTH8mIzCdx/
tgWlMxNi55gnh0Idp71gnS7RqeA18gjuBaJMn+smYLM3VGGyFRtMm6AGyyOY2IkPeq6fQApMSw7b
51G7x5Jo2c+UW6284w2/IPCHnGMMrOW2TwF57TPYzhanm/3Ki7FlZH6FHFk8CysAviEcRWjVJuye
A33fsZbCz6HRDupzkEVstDo3Wh/L1UPEeL9PSqrzpXRUoz2YEGikKFKAUkf29nKK2cguwySffhcj
0trbGouQswzNxyQdy4eBJRbUUSkfeIOjTtyXOaWHqDk95vorCLnUoNz8mYmh3GfwEHpMKLxCeJaM
8wD7Vl7ugkH55g9FAnfA0oBboAYvk8WxYJjvZZ7Q1xj8cSv6jGGYhgm5fPxi7fkRqYjcw+oTVTjN
SpkKopZ0fqYr6xIa90P6p6wGewO628LxYESejNtrlVRqM3qDLTi5XzbLkKR29ByQ25QUHYexFmOC
TUeu0LKoG3Ogiv/b2jySwhPJTWgloMroTPahIldKXQkwSs9bh6eNe52WoWuMepUIJDDJU4GtPunI
IzCs1Kx84lhx0DnfE/l4mQTvuxnVl64DFS2hABoH9Z7IVva9vhFHBYSNb502qQBBysnQmvnnsTjM
jHudATdKMxhDJLu7wU9f+A9APzZkmm0QB8tkrTKTV9VFGtEn2G6KoTKiDYnNv1j7Sh+QNk5OTJS5
6gQp/NE9s4jrm6yuaAGXypiWWegTgWvyovrvRspQYjMhjI8ba2rMxtwbccTB/sBotpZcz6jX6UK5
azLsy4dLwxs8vqKdw85O2dBM7sjRgZ6wpDkf+ZsCDGsQ/NXa4TiaPQBgElJzojj5hLIJmqXAUdo4
sJ/o9SU+RbY9k4u0stbsmI49YIsl8aAAPxqR1Nqd/oNeVdnBwoimkdjXLkAdYMeZ+fEwCSPu/BrJ
F2mMuN3pphyalHO//1aj4oOXLUjoqLs8721wUZaRGVAEaWUnOo56uDWhfLZfLlZIrBk7YkajA4qB
3qxZGoTuMMfxrOVf6QW6woo/G9UcKFBA6MUw9IKSS8wQYOmOm3V0P/TflgX9XR2DiL+RHHxDXYQk
x/3NIjuIdROS1xO+SYbtMCiYD0k347Ga1Z0LRKViFkVkls3+njr1a9tsiorVGwbQ7nhV2iL+E5C2
0lkR5oRnW0hzTIWEilDbxcOfWEIJ7MJyD8ohVN4uSehRQefBCPPyLSDnX82S904mO3HOqzrT03Th
biRTqdKTioZyZ1IMdoJeY5EbNZ5zPDTDIooyVKccT4D7xHrZGwZ/EQ46z/yAheezDshirZcGVD80
pS+5d4gi+Ehl1I23GYpu1ltLnO/wQxMoXHLFhSsG3GATzAUbMLqp9kqjJXRCO0c4LqC1HbYoUatb
zs1MPwJ96Cx3LJXQWc7V8idaRpIKpeiAUSZVKYYSXdQYiCmgUsjo3L8nInrSYlfiEsQSonKoScfR
byJP17rutFd49kceJvtN0JpvPcVuAV8DlOMtm4Zr3TOVOPxnKl19n7jLHYHE5ESOY4vGxCeyMWWw
bLJ//nzG3AS0tP8/U+jO6bKZnJOcDZ4VVuCosb/FqrIcfebmxpsm5TohHnoVNwYqUBosL9WaFGvz
DgExeQlqFVbMjOwRrIk4ygyS9IzGtJ76vcsTqW0EuffVFyGb9/ioCm+b8YOoA2ZakdL4hQt2eUB5
Ltn2j0Eg3E9u/JvT/sDCptu/LgwrmZN8mjdakJHnhNjTj+M+uc+HRWWP2NpDVbgyHrizPvRwWdC1
YfLb+eBXiDUkebBi2vuCbto8pvALb86HnBILvBp6blfSUHf57XSE7DLewKjet1uP56VSaPsM0eEg
jYRMZvXAS5vEwghiXESE5XMWHPoG3lM2ElMaDE0KotkHPZcDVxVOQokHzNE2LgeTZ0+0OP4XO1th
MhipXiM5YAJN4wrjOLHxPEn0UKubB5GV5cFzl+S4SuQ2SEtei+26fGM6bUSzv2ytYg7q746UAk2h
smy4WwKqanS/kTTV8BWaE4DRKC9P3HYdjdiqj/98AWjeh/U125K0C2UjHUeGWqCwOVlW3C5njBg/
ybA6txjz5mwmu74GO2EGmVdTMqYNIJhPLl0qCDTkYsCwpRlWLBTZpqSJROXn20jpFQF875wG3Ek2
b8vczcmvHYgg5GbkcdasHRVSsXMIxkN207yBYJT2Xz9EvkjK38hjF59Wf8Zt7y1YuYYSgU8SYC8o
QXMuW0bEF2G6qlMo+bjaSD+EU4zMIOVh8uvkNZ3ncRwhsmSktmIFae/HowHN1vzXQQ/ocqi4MrVv
dxV/gW5Rds5kzJb4HNmBH0kk6TDf7LYIyoaZTD0/ihrLTkajztK3Pv1yuH/gTUCR50KS4q92ya5s
iM/6Y01oFuAeHMbvr/otdEoiz3QoX/LTiZWcWe6x2YtxSGoqPt47690RCzd+QqqeRLR8mNCks3nB
KeBRDIed5HjzRumGDnrQuvTNYrFtaqdz72El/JqhUJD7JdQpFBKjut+2GaxuzRX/aZrAa18C1R6r
9GBq4ESFtnaPZcs7OEdMgae4jFqwCJFtE0Ozbs4YLH3YOQlJl34U55QR9uXVpd4tCKcxqbdDdSF4
GK+LMNyp4QNrIPuFDHjBApA2M0OGj23qZ2LQWijUi0gvsJqncTqsnKmIuNqJhbtJxLPwpYfRpMC8
gg+0WrSqyfkkevoGBwvym7E7EB9f1kinIvcBISL2MBtO5vFAn19loRm1wUWI0mdWgV5G+RUWO0VQ
uapU5QFXpPDFWST6rJuBsEnlLrjmCvuSemtLshj0w24TduS8cgm/JPUtQNG2Piyljqm4ZYJDQILN
ROIdVvTCLpM1ah7n1XcD+UXGUPM92ZUvFo1Sdj/6GT/qTn51bHHC/BqislOS7eaOR0EoThV3gV9N
mkl2x6hfYfllwCAfWezmWfNIfVgr1qdeX6B8Q5CnA9M6u/p9u3pwVCCgyYGHPLZ2tUg0e30IITQF
dhWN+dXoRtQbFiL4yJSNqeIx3ru3IG5mHH1ERJtp+WGHYV5Xg64LsMznB9sjWqbVbt/ZrwSqYlWM
uMPPbVtRpb48nsfXx8n8q2EsYgCu2GbM9a7BkuVClcnr0o5DYuhrher+YZSCMyduiRVEMKdq9+1e
XdEgyr2aczTk7P4Cg7lJv6ZLUkVZlwSCHMEEfKdIDYJpFRxv+HxuNpqrz4UGEIiLNA0tGopMv2jF
hPk2nYY4Q2737OjHysFSJN3MPUb3g5zKmB8N4CJyyobCYoUZQFjRsJk2ccbyFXIC4xd7Q3EvhRh6
BXpjjYH634h+aXwet/l5/dPUYFv/B8uU2SCzmNGsHeSfjnrFOuA3TGqx4gDw4K/jolcFh16Qn/r3
ptNEnXroiWa7J2aD7J4bm0jfo3QD08XAcTKJTfld8QjP6uAFuQIn7Ya/aAadkJpSX6wBN9JjfJ+W
jpeSWGTwaEm58VIUNp44lACH9rZ3Bo+XqJk/833Nz8yHr3eEbHBbqgWtdQxqL+YOER1kcvoLGpmg
RBdAZDsFwKPP1vghHnv7L8S4Ri+aGy1/I+RopqfSJr+BTmGxutv2vk3EyHiN9n5B13ZX/13AyDyw
Kfp4XOc1Slu8gw0wtBHeoIdGhERAKoqv4M9jJ5ZZpkosZzpsO1nsFwLZ8orQrwtYOmtVcUNjDyjm
4iL70lCxattihs1BUPxUat2lY4f/JLh2acLO0Ki/SjfXAeJOHITZjVciJhCQmWS+Q0kaC9gZ+MWF
VgDPwX+ybilnQI3+G3QIzbLUddfY+5Qlx+XApwlXhsNjPgBZgLy0reooH3JvKAM6eMUc4ID8roqu
bx/kZ/iXA0Uv8F3f9D6iEDTVGHucoWGcoxPKeV+HVlYhMTW4pqcTjYXhK5ONk41x269eWPOFOh9n
u8bYKhjIY4CF3bOivSaeviO6MRKkFu0X48C59W+m2UKhZVSKk4wrt2cWNyXKS3+QOwLvKSbbxqRa
/ykAbyuhs9EUqOLyRw3WpgJs9PLA5l8igqhYrUWG4pG7uvJy8w79nnSmQokprMhR/HsjFx6wUTu7
Ud2J958LpX82RTGQM/0Fc2KZyKmJ8nPUikgDK9b1LZlKbUjQOmvxRfMa9Y9bSVOFifbcVigWDlpM
E24zj+P06DszunyKw2bPSDSmTXqzpuUn9athmh75wzcUYOK5y2mXWlC1vf3CWCFDjXcXfV/5ZPO9
vGkgge+r1wKl9EuvGKsm1sZgxqj0zffGPLPuN4HeW+9yqkAo7T7Wt1duG/gQfDNW3fQwq9UGSkYF
k62EDz1J85KA5biCFEfk63NhX9pIwi419sV/SPiW00cROTkEXsDDomVFSnzRg2ZWXjVXMG5HwsYx
dPKZp7YR5ruGCBLZYmynUZZC37+dVhR7Uz7dViLrY78L3hrPNDKCPN5U/9GWQAxP8XMBQJZ+kGHP
PlXcJKe8ljBRl5fLipmno4b1b4BOwks3HMkkKG48gKQGAuHeFdPCti8HTz2cZFGwMfqRLyYDvN9W
0Hz4hLblImCvVZhtPDFYcNskhpc5d58Eh6sVNZuERwKBoV4JDN0+EuzSYTevszLzfvAXQLuWtywU
oBtbaUuC2EBXm62gRHt2EJQbe+SF07DrMppUKNvmTl/mYKp0G18xLJTA+IYYbR3dPuPOErYWT8hb
cv1GyGHkjHOpDbx8Q0LHn0pCUGcitNtWSR7m/0dTJNcfH1NFQrH7fjPP4m34PeCJLdr9Zdli7091
05rrVDY0awr5Cdw7AIlUDBOcEmEa9uGX0eQ8GBKuaxHyIQhbZEGZ+H7JNel5T4aRTcoWgeiVfF6n
vT1gT/zlCu/kFP1R7YfpM4ToV96IZd+dtZMFLqUIhok6HZMMUZhtIygk6BYiCLB2Mu4T7Hn+1Unx
7YNDL2C4ivMqoaYeHxy2VWzRfTmiFGyo7tel9ezm4ZNlWkrqNuNee2UPqgYYDn1tmkU5FwLamnBW
sOQIk8w6n4XcC6PffNeNSEGpIXrx/5iSHu6ACwR2Z51T8ydtCSorpGjX1HpPpUJbez1fnJO4Gu6+
fkZpvo7Stk7GjkPaPquPLMvbXyiTE6bw680++TCWk76ScWpCAfNU8BlYqjN9FoLemYGeVfVVzw5G
oodN1+QEz5I/k33IUO1B6s8EjeAyIndkNxT12UuCq4my01PfdlVZmNDygYEaBDN9tmPIRhiTY9rM
7HVZRJuEF3EVsYjm5m1VcK4+jp8yBAurZdAy27hYnjDs8FF47mkl2G1kI+zl4spF0mU/KG3gYseS
UHZnmeO3m01OBnHjq/3grUuB/608GOFlKUSrXbDuTpq9whjRySOGONf5asEt5moZrom2we173NFs
ddI5/6V8JEqTu1ZcORPjuH8NyrM786Q2OUcW3M/mazSHwGn5fO6/e6/MZ/Q7PbavjpJj/NWpqoBx
964bPDy0rTIedIO5QIKiiuNimbQ0+KyHxuUrkCjzEctS+YXxNjrH6Iz9ZZO3zGYBE2zjSWyou0Mh
4FEOrkVs7wFrJXJ6kWjFhupdNQSvwvwjGUrW8H8YgHIRrgdO0LjxcF5GovcQ7MqACZqG0OUbjfe/
VRJOq8KZdOaqY3++Ep5qiFPvNmJ9lS9ycGBbFdWQCU8PGQlPTNSzJ5hSWz1LZ4b+Vs0zqCU01hlp
XKy2Zp7imH2ZvGUgN+3iFdJtR8BslUqy4KdW4QxRRzg/h7Wb31Zb89jXOj7r/wzW3BgFbDyhuvIN
N9AJgokcMdqnAzRhIGs281IrO6boQHcaPxmF+GTuBF0NJZqrRReH7VZ8+03Qq8t8zpX7FcisXkwY
y6ydYlL7weWfgFERGmuTs2kEY22QI5XlJPavMX2WTe3vA68qhErEOG0tEV/ImJ+p2ze/oSJHVE7h
ZKG0qXAgpKQnRL4V9grYCXlQJmPaX1N3C7mgzS3nk+KQqjq3uTjrdzbsI2PPEOlkSWk/N4no6fzB
R8OXUJMLYZ+kCDM19aCiisvNNzWLaX1sIlHW5YD7qnJGnvysgpRG/oe/49rfhwe8UApzP5Mm/vZ7
ia8SAkLFzeYKLc/Vq0uZ9CAgFVnQ+P+ex0W91KcHKcvhnW/fq99ti6kmwqRXratCscTZ2K97/qXH
kasuLqqbw0S1/IqmyM2qtOrVHqft9LT/RF4pVHdlqX4hzB8WmJjDpXODsObqBKjA+nLHy16TF2Ap
keDtEtUF0ODQqMeY3k7obK5ey/12CxxnFXy0cmEGKPg8dzb2w/k0nnISeKyH1HNwsk2hWTFFAh7B
hXKY42rW5T5w2RxA4ywXzHor3QjH0rO0HlRPyF0GTX86hOvJ99H5ke3d+rQWC3sGcZdjdqWjlT9H
+MLsH5WgHte/OO5ZRbFe0IdrCjwL0fhDbQARFTR5paPpUC4mGCvUFi0UWzD671pY1n5vtEeGBWXx
Mul2stlDlnHq5G0abewS9WT42y0lTLKevs9Q2wI4F15VLnyzXHRYUg222rPBDtIsO8kXiTT0mELk
O8zia6AKmX4hH4hcovSUbrZRV3mxaEz/P3wHWsQVXpqyMFioCKUZ+TJ6RQBVgaU39F8MIKYXtvGe
nrwLPRlwAgJDP3zkC0Jh3v8ra7vkfYvDwdvcJZrhW5DPvfVkjKTgjc3+aU+rMyphv2mJwMkB13Za
7FBNfL1Gvh7yqV+h6YiXz5CFNMtBYwcHaUq7H5hk8Bq7L2dUhFmY3m/ivEl4Iq0jcd10tPedozb8
FzY64B/3qcw+f3aDddYWjPM2Qus4N/cBL3M66exepClkDzj6+Ty6gQmNZSVYWTZKw22X4OVoR5HC
Fd9SyGQ1qjFrze4zSZE2QmxPZFRG2iCrDrGMTKH4NUbcLQz8JZLtx1hDBjf0QLw77noah/H/1vqC
Y1lFpTsJ74g0J/k1sNzBxuAT1mRMYcGYBbEUpVv9g/YbfDO0ZSQ8SAUTB7watZmruiIZAXBgseHL
ZV6HB11IJCrEPZcInduqzdhn8hMAXFoxFZ1VKqSY3xvm/fiNrOYJaYnadDwTDAwXF+tH6jtIdD5Q
ucxRxEHoeyTEoziAzlgzs1GF02P4qAG7xWofCl1ArBCkAxl/Gtjbc95uf+5+TOr57cr8RZpTi9A6
UHeEqdw+cSBl2LXqTVX3nyVYKcQ2vJBrVaT1fiH7b4aNNpRneQ+pyEF3J0OaajqFLJPjjQwZuxCa
1loV0FbzyG3g0V9mRdROxaUB9PeFyOsu42x03EQkqCM/XB5AyoV9qXF9gqlUgG+OPcfUdW+yQo3i
QBAubnqNIbSEtIeQQJswRVYnuEdk57OHY/io6mhZx0wpMH43jnu9jCuvucE1xfJTKEHmd4gbL/ub
4WopwNc/xAcQY5m/7w0VPVPoa+r3I7g5GEiKtNitwMnxPgxvj9HGDoC3QH5OUd7zqVfQo/39FWnM
h3EGafgZDzp8DRaxEDPInJaCiZng+pUSLpynWo+zRzXM44WkgG/JYvRSjxgtWXRLGcDmd435vmko
cej/51KgjAddAAPteHzaRtH2gBxNj+rrxd1FwEHdqL3rpVvUKwuYAcDPd/va/85qGzNFdbBRAL/F
KDlxbEEfHC48x5BfVk4OSYULs5HfXOw+zyD2mAwBA5KbW5fSh9Qa9J9ZOY00IuacrHsmoJeoUmzU
+0RmiRLe6bjILVOHPmfXKPV67LhY6vVqdFIecc2GDGyaeoHVQjej0DQfFLulNl/boQjhoj7+vCFk
WLOaA4fWVToZd/dOKoQg6D79E3TbkQvyrIvjqIdRu03FYjo3xvTj5MHjiLgBg8ewUo1ZcRVoEEgd
Nyda2KrfzuOUBPxuko2+uLNg7DYgtCPdyfePBPsA2YaSZDnNz4Xd0kDaLHUJOMTWvKJbbTVJlZ9f
SdkrATHAShqDnxeWUwCbGxjWdrB1Ds0xrQBBX9F5MrSQ7TJxI9h66LV2JDhnPCT00H7BxBoSu5XG
XFQg3CSW+OVn+0KpN1zYi56qI9ZBzsh9w4wYkCvIguG2WzhOtxW2RlJh94epwedg78pvagqbq/sj
i+3fxzOmzaniiFiKelu4w2ot8XW5JjfEvZQDmdl0YmcGa9z4O29GO65/BFqJDBhUJHWttJO1miEW
3MyXB5ZUKnhLyPRvcLgADMb/b0ZjjhNCKgQCm6H+T9TWNNyTUi88H4YKtqZjxsA5EZyWpVOBf1MW
tKEoX+s3muBKgaWZAJb0MXLv5Td+K+X7dWT7Enk/3doHU9zVHeMr5yZ65YSGJ/qB36e/OR5NQH2T
4s+RxZQj5Zv/L5HSosEMBkQPxSjomSv5U1AY9NuzLqg7ZC1mO86nLmPIwOmB0bUJBXvawpF7gY6i
Lhj7C6rLpje4EYsg/XwaVPFRPuezL8ct2yq0iZls8J3m1tNQdsjxUfVracgs54IQMREuApn376fA
LsLKS9pVkqWFohTl1wJku9uPn0HOBMx6kgFwPzf8a8RiSSt5PjBgt+yrBjLSAXRMjI1MyUY/Xnj6
/WvWlroF4rZw0lTmLJ6Mv2yl5oYUmVFDHG5WCoDh6W45ZcL39Iko2ulomNz4MBbgPBLNsXi8L90u
5Vd6PbblP2NFlQp+IkBElKVecaWQ/JG55T0Sjz9k/vs2AiimdX76j9udBwlLxdtOE1B2hOvtsgCp
5JAY2g3ylJQc865/sV/4nSUbOrRSZKEXABdspNZ6KRNIIHHmqyEfmSuYq7Ye/0CGeriTJoR1+WYg
YfS351nThsAak58tHK+S4RN8OBKgXJ/fbTXc6RgnEs6ETSFsWYMBXlRSGEwdixMILWeWgSQXLpzo
tLE6VXAzZVPnx/2JsoZEa5ClGI60SSVO0cUxIUiEI+vZMmi7hmDssZq7L+YmCYRoFYyijLpoCNS0
C7fGWU7i0nIKlazHovfaJdagDhEyVBMhrPbIWjYTOn+WUSP18o6mJpnu4HsQOQUoYUVu7dmcf1vd
mhChCAiDBPz+I+a2G83ZjGksVLyLQR1pU9L5KqzCdQHD1AWQrCV6y4h+yVVsu2cxMOVy12goU7EJ
DFD+ENWfYg4Zw66nQ74YH0cvrNDX3iEOySlEsaG3yXy0UrrgLd5A3NXl0ALPQVCwJvgLPwpoeGij
k9g8eHPI2k/ZTjwyY1Y2TevjcYk6AUO5yc+4B8+GPXx2Yk9Tpkvw1IOgQTbtDy9rSR0B9NfWq7MY
exuc5T6G5kQMr2YNXWn3N5tsaxJu5hed1ztzOUhowiC8SpMrkXwxALJSxc6kTLEJwWSS0PFbR1Bb
HxmdI/29hTPj1eKWlC3NGnpm8xT3vEUlbQhHsKlrtGnDvsE/17WdNH9u1ymBeKZP1s8/fOZ9lXLG
b34pexacgpp3k5nbereFMNh36SpMWY/D2N2F5RJfgz/95/6ZVyazaxyf1Wnr05lMC/ykfvoWFmX8
rhqkn7Yrv/bRXfeP3GzBaZUWoWCHLDRpK9epyRIhgTlkbq0mB29A9LW0DPQy1kKLX6u+Fp8thxd9
HOTsmwlIRPdE8aibsXh5s59eVOsspHE4i9NgwERMBRxp8owaGZkLhnU4kVJykPMRoHiqa/E/wtEd
YY9QVz5O5CVKipX/utDp8fSaI7qesRjqewVHnmh9o5BKouyb02oTePsbpVAzpcQsQ+A8bN4PfXb/
j3sgh0FT7rZuZLgBBZm2tF3a+IrTcIeSmoPOZECu9bKj9uUulsaXHqMqlTQGPil2YpGR1mMLqV8k
DMkl/uv2PhOX/macCndag7S0Z6cXU1zkD2rQLW9X+WPZfV8NZSnU0MwW90PGTZqg0zEy80brkVsw
UNsprDADqVUbDhGiuUSRlFakZQMxiCPCEnhHT3iQuqHeIU1F7AJ+AJkHGbU/QMxed0bgN3vuHmeV
3vKx+zFHKmhanM24YzF7/lkdi5ycpjBjQuJOlOVQAzrtkTWYP2h7j0R/Lwrit7gATo+szNvZYgHq
U+Po0TlMNkVSm/KrrS4DohWRd6YoG4VEC96KyN/Gt5CQwhXqC6vQqCghRfzrdwHv/5i8zu6Shjsj
HEPpi5/Dss40PWic8xDnHT83iRKvzQibKljvHGUyLFtXmXTRb9ewN6UUDk10D6HnEqzMAt6KeRzp
Gygdu7lFNZcCu6rg91Ds68ZT40WJi/qiSy1UYWhZIEXZqoRXg6zgHNcY5pa6jvAdAzFA583zqBWh
rG+3Npc0Eri0a6+cW+pHD/Lm4q2tbYnXtFHGFo9bxS2qFOiO4Q9cuiQi3Aj4iaS2dL+tyv2ec/CD
qcn23qcmvcd6DsSIoj0TUSxxQaQmEgOWMd0HVLrJ7XiKKT4YU32Rn9Xr4pvWfZ7Wof5j1WILFRo4
el2HFNxKi5MyNL3ameXsvJ8DAldF90v1cjQmP2xPlKLPqQO/QtHH8jasrrt4VF0YfjJT/WvE05zh
5DLAb1iq928/2pzont4MkChi9zuaLm4cPkHNQ4Y6JKL/dim5n4gfxYyw7v9WaQpcPUmdCuntAhz9
pn7GfNmKubqPjIvcK7ZvzwIikzvgCV46DJbSmKjFd1VfZbsI3E4w2Gh88rr2rn6ELwOcGZZs1b6m
yDsMP5exoeK5pErf1GdS2jK3Ri0Z8BdYX6ulktYZO8hjlN6TNpvN2ZFmlYsDfwQ8Lkh1LGSQeAYk
MBs5yagiOdWuRaoRV/zHJVPM2BuuyqRkGl7rO0/ZokEocozW5qtbvCFoUj4Hyn7XqCRTKVyiSZA+
HAqoMBf4QVI+x+FwGe4WwJ4nWr/7IItnOP46jn580FOpotja6AcR1T45PZAlQB5ojHyWbzUpIbbQ
Q5xXVE8aChLtG53qfo16zIuEoFP9qrDZFwPheUkZyFW0gbvVTTBj8RiNPCdv3wBWdvGpOo9mVmkt
6z5m1029EbZGki0uZ4q7WGWdln8SCBjtm/Z40iV+0kSIVcLj6GdlkvSNe0j2i/2pTsPn9u9jHqxG
XFj7wosXo2+O1wu6VVgoGcKQvHiDv6F5B/MAYibrIvEVyTp/oMO0HpvRQp3ZTkcccyjtYWXVTmuf
pRFsPIzdwrgIPJjkTihPrSZtuMNYz76nrnrLumvg1UXzQNkFTg2uvc4uR5RdgX5qNBsegJmlhw1a
rGhb8Ho5q5XgRmL34evHfty21Cs3+cqWWPydLy7b8ntvt9bjY/s02d6uR/HXesVplXaCgqxDjibv
Tkg5Oh1SrkrrgmrOmAeG3BgtZBbfU+NLjyfBAKL+q/fv1cezK65DWy5pRnr2hyAzvhlQYMG84W4Q
Ul1ge0Wqq2Jj4nT263HU1HA8k1U2SJy8kWFSPSFyPE3dZZ01I/NLSebeuhMvHDu3d3Zm/MwUVTR6
RUlZKb1QjGdmtAhp2D51JHrQmlENlCVRxtKzSnasC7MK1IvbytqWiAlJ6mmrO1vlL2tFPHlXPWAj
oIFsHmqP6BI234Ob15xKgbxWj/JR2NZcV0ZYEizyNYnyfD8+oVj5KoDPwVPdOOb0II6W5cznUt+8
ZtWovSnBM8NtDLBGHsI+rLnH9ww1jsSpoeVrjYUuqCi7IieE+Bg+bFfOMQrJNvyGzBI7KsO1+dEF
1F37HlINe33Caa6GC8QvVt/CZeBi1HA4+NuGNEP4SUpc8WVZHiQ7nAAGz8oJzXGd4d59voPn6cc7
VrGQ7ynq3Qs15CXCog/vvhBjjH3MT0SKZPsAFDCzVXOlaFWRVOApwFU625UdDp3EJfMjPFetLE6g
sXGLqvaSpTIqiKpt67TYMd64plIpA7oMj84XqBa8A0atXX0e9a4iptzFyg+Q+/Avm7CuQHza2RQW
FT+dn4K3bBBLLy5g4xgEmhhEADCho1P/Cq71YOsCnlwxp3gwaDSMGNP6e5rnPIOPEJ+5tWIEQLOp
Q2Ahueo/CZFeLB0SkBcPKhyB07Migt/1W1jeHr83hZhElIMcAXfn64htrxOy7+fu8mo6zCMNIBzR
+Rc1JyVrQdeXyFZOtAq5CrGnwbjsVuIJSIZH7wmrkFhbG/m/+wb3dBl+4n4YRx59NzHHjat7jGZp
ec+LfudqtnOk0//p24bzydzONF+6eGWhToHYLgdnpW0Ce3bByxW9Aebq847LX4fNKHMWDZbJtLwQ
+uIc+/Rv2Eifln6UTosFFYhFBXJ/gJlWFrEBBoh2sgu/ZIe3DdCqBvxkryJn7x3AFpndKBXkGt9v
+ZRxDw9lzj5mHxbV+jVl69OFowCyR6GnGrIGX5vFDXb0O345Hni2gR21sHSUWSHvSUPN2zUlhtZs
EaMGz183Qvju3umcI3jIjqK0ClVVcB+O2jLZanSPZ+TijXnzEgUMNTvhrVDOaCrbCI5LMRKeKCY0
v6B0CcbJqXo0W4Rq+HsD7+jYehgL6fOhdJoqUXk0EMRslYBOlVKrTUL8+iworUlZ+8yAyam10NH5
mx/ERbCsBNKvGNXuAf0/DkZEZZqRe0lvnMkD3H1AahueQit5/wCQlc1ViuKkp/0gSSACmY8NXDlj
ha/eFV622Pzbv+nccm58Ou8TD/s3nE3eDSnaMA5b60OxggNrmXYEsDV1A0N9ZPYMx2VOkuNTdNLu
XwB6J80hH1i3Pc1tbRq/MUDi0XP4z8qn5JSRQlVOGbq/22vhw1fltWDtgzDNUr2BLmw29zDXRNGW
pnyUydAt1/ZSAliYkyouQyCZGI7WSrFuxlGapxSyuQ4oLFPSGu0IY+RTmHbjRZHIdn+31qQ7O+UN
JYhEx2t1cnO3fbHE21z3Vvgg0/dHxG43qCd4WgRdxKrIajcQjAmJUeXUA4Z/U0oXFi+6DLR0xayu
8shkn5OQ2vfgqJmE6ad5grHpNu+BRoYFYBmEBOMZu3FRpxiO8Ffq0AyY88L0caONjYPr3J8Dlgez
entpg1iidnTgPscgGnJm0JQ+AZPAFzRtuOFpuJSj5gbWRaRcyqDeCv3EHVhBQKObV9VkjplmsJMa
DgIZAodSXerW2yQkhAnocXnM43SNjJmBn3LJF9capE4+ZI0QvrhEFLXIGzYeC9iCY4J23UPTehGn
qD9utZLmw95PcZELGbFP3ih6oRu3eD6NmLxdp1DaAYt+/Qk9GG0C5gTfS7VJIln5X3j5JY8JzxJJ
OOV7osnS3X9AXyzbi4MlH7DvTqn28CkJWMZtksl0J6A6XoQYH346TytSvQcWaNUwexngJwxOpk1B
aSM9H9x1ZZSThbmw6LKrbWouCf2rhNP3sh3NULnOw+cMTvtQdFc4abGN+31LOS8wNVLwn2XmUBvG
3sEVuj4pvFzqyaQqUFpXwoBRO1BQ6zXKY91tsQ1gWzKYgD6VXGzCYuMgr9a6hT5zGucvXg9euvv1
3acfLbp0T+r+nwN2npcj5FYfUvVYaXE3MY8l3AqW4Gd+X3Lvw5Axb7c5NbaRKh32T5nxMOaSd2eL
9aT3ZrzEHVeU7pu3lljzRP+opFedJ/kRSHQ0BEwTyNgVEr0IuxXKi+c3HG/EONv2XFQzqn8yvwGd
C/Na5nL0QuyRJCToFqQlNSfWTd3/NPd7wLvIK6tWTIKc0yTKX9IunJ5rlL+ltDgIXuiEM436DXAc
3ulyUYFmU+btySU1ToKaFSgOPgi0Ig+AoNMjtX0n2N3sHCtxXE2jQuDb8NwiUn6+J7muzO3uv/It
mwRQ1Uvp+ltZ0X0QjElNjZToQBg2IM8fMhtTMwAC4Tv2EnZFqI/3zqiNTqh6uXJdFa7Dux+8D2tm
WwYi7MF7hbnDTM94W6V4v2vYjGVG1hgmamrMMhOtffxXnCY72erG8WDfmQi4exwH7AJWocjX6/Zo
xnMacGq4DiGh9V41swFEZ7QurSVelzm0VrdN5Ww5BwjDdR9to7I2wJ0gaTwvkcFcux2Ywp5UfIZR
GmYEOC8RIawlT8kQEAgGjzdkjwaJS1p/S2ds5k6g9JupieIa/WRgVQ8FRm3c0yjjJoS/TsckR7pn
ynADIOyb8o64bKJLQEK7wvgVtZfQrC7hT/kloVV/bxKyMzqUND/kdJnuKru3/RT+PWZ8PuUFAhSI
TPdgCxtV9uTT6J93xAvO5gl4gcqheH6eQncBQkjwHnjtQkxiU8YKodlvVEOQhkhfwH4OQtCriWyT
z58JCu6MtXG1ai6GX9d4nMNj6cl7nu81DWQf3JPbdnUVCBQfCI8J9RLuHpSzPMAltVN6c/up8qAn
E+c86agvwNObRR4N0gLV7OQ82XM9yvNB5w2ssrYvCuTZhMu1c1wa9+6fnRduSLCWdE9o7hsipOFQ
nXoo8jEjPZoxYbV6cRPDg6ZHb8z3ULWHpqy72W8LydzP6cranxTmRCXYKE9/grqot3oc2YWMylUE
41Lr9SWY+SdfK9jAYNaecmwlDrKo2i+aPO56mLznW4zXhjgBoR/lI+dtO0zdCZU30++iGT9/SzE4
za73kFcOCS+VGen0/TuSHBgDlVWdaCihnURuU/hKiYCMxMuVm83mfE5fLvvEFNf2jr4yVv75jIvB
xlhpTRzHxApHVSFPJzZM4GMY1QXuEI0dgyQgPI/uS8VcFW6OTfsKYmkV4aUwIpCUm37pN4evgD31
tWqPvqgQ0KWu60pcXOZxrtKOGaoLS+KwfxmaP2aw0+Oiby8ydIkQscNEnHJF6oE7VjtPHOtiFkkP
52+l11obcfvr7YgS/myhrvNstxBG2e9m6oDXAXLG9iWvBFhO336LHO3tYF0SeFvb6JUbiBs6OQ+k
N6XI47tPUZFVN2n8ETw86pMoz/KLK94lgK0PWloHhE6C4Qj9VNvn3icARSlvchrSaID7uLVn1chL
64TFaRIt6XIS3TBkmYNaHk0Lh1hadd/L33XD13yjNkDZOYXw5kq33E566mUdxiX4sRuxPgF1yZ2B
esYP877z1kRmt7lqC17QLU8146aY2zaH/EVosTT5OQBbaSW/vMvHNhqtRRCwRXmIpObHgPGB8gFb
u5R6S7PwO7NczHicocaK5FXX1NkYAvrNwyxilEodBpgMBw5HY1v5KQdzfl1H/h0WE2WjLEtaoHcL
6tMVFZ2hrEok+hd4M7mQJHAfWIC+/xC1/gswHXtXy3TXRtgLVxVk6k7HZL1hgkXnp35I9BlM85n6
n/49vx86fbKUAd/k7EpGHfmF2I61nLI8Up+6EN8a1hXiGEdchkK+Si1aUx9AfZZ35a/Fqu7B1cch
fcOlsiICFf94BG6XSgVSswvOjcjS8XgTHwQcSfQTj5g2oaX3dLobcGQIPSQQvGrT/dlDe/LpqIAW
XUNv3biSAsZtE/RxgwsKquZ2uMf1attAgpHxXmrBghj8KLAjZgj3UFRwHplvT6uEru2drGiWnVYU
JopBwmUZ8JwV6S/9vL0L634Lepl+ixdlwXL2qkg+mGbrbIDjuV1QdA2oA5d+75tgeVa1LeAieI0R
hGTtgxoehEB8dcjQL9qByyd+ODrSBO/lFPfn+dhi39NVeichbBrCkdMrLeWPJpm+r6PjwTNhBcFN
FUqB+9jJsDymYsPsWsWj/Tk3cZ7SbDL/q7vuNYBSe0z/uZ9UIpk0Ebwz44VRh7HqiuViyR7zRiMG
oCkIl1IWR24d+57I4V5r3m8vieMP20R7P7Tkt5AX4deaujX4jc3WOZiLeecsFgBDWuedBbme/nqY
IBvSA8UmHllEOb8jRnwN2Zn8nZZRzObeIObBFTW3iFwPtLXsIx9TZgXBHmGO7q3v8g/+NeA25g4h
r+c8m4cKKOl8bACbDnOjJfeSJ1fN7CyLnBMm9FONfZDpdKGcQkRhnRNBJWUOeqfixYVs6v3UKCAN
G/fZkSZjEKtYuBYk/gR1ANWOyH8EqIqQ/Sry7uUQaIurGIuHfkp5hCQjOJ45XEGHQPa8uPFfFQyV
N2GMgc2LP+AMJE/U45BU/rZXkpWjlrxSlzUUrjrHLfJRwVcvaKHik7V9PzzZsN5Xj3aLbgQTmu/j
eF5SDBDBYqgJw2M2u/naktdUqgRHMz+fiBKt3OBWVorZGtjIC+c76+3nWvuTLHtvtymlX3DGnnD6
07qoD7WKfUHqcKcUl1Qb2DOqDRxJPRqYc0k9M+ltvEI7t3WS/UyTd27Pw4g3yz3Z4op/zAz29lxt
cQlJQwgFvE7Uda62eHv2G95nVBnpNFuWfGQECa26r9BVoxqP+18IHRlHyV8KLRrCVJJ/gTBA59MI
Xjyf7+1PiwtsAKJUb8lfJkDDIgVWmRYxVf3r33zlMJMsbglzgvj2etqn2D5yhJf0dA7lH8WmZxk/
SjXQwAk+Vxjvjlxc4b/6oK4wktU7xT+IS0yTWN2+PIj1Qjp+XKMWgji5FFWDdkgzWyDss4rJ1RQb
Eq8oUjgkj9dD6zTFoY8bYerKWqHilZgUz472ii0ixtZL/D5TZVrytHZB5vchcRMoyW5ib3oSgOQA
6VCB/63ZHeQvkkRLoLHOD+iBX+GzFzm99lZKqP7WB+FKfgB21wGg6j6YhhIjoKRQ193eeQ5dW+Yy
k3MR1oOfrj4NRRfTLWH1BtLncLzFiZzBWZP2W/xRDuXXanNYT2xRoc/VI+UAStrAHOSI+m7Eb8QY
uY952cGQXRIJJhMTpaYh3EDIPSsi1iGkas8CykD7BCz/hitU63BD3OmhfWSv58BlDjODx356u9Qj
bh4fCbW7fXllVv4TjOaat488WKD2cNkocaOhMHdKWJnOPPtW0oUZBz7xiQHhKuCG19K4sPcSkywM
9YYn6mwpd1TRUhcQPJn0MhDT/4FepujVaibZieeR/0TzHRDFslKlFCMKaIy9zOPjSG+Aqr5QLgaY
0P7DFMj3/O/372IUbzGGgOO8HU3ojE6onqajNV0uWPAsLmiLoLRSZD0eVGhc52eLPC04S/3xW2R9
+Ma4h8Ev8ZvWOFF8Estks/Ym3NI/J1tUfPde+Eia/BICwetKvjiQ/vn2xzG9WqnFpTLGMOWDyz7c
Rny2CgkeaKd63E7f3fEC7KN8acydg8pwqB0XigbnR+WPdbD/rAZ4QoDFraZVrTboY6jmwcuD4d/0
qUrtlEZF0RflnB7odT6ISqyqxzRdCvvRZi6K/yZ9sMJV3s+6+D+l91Y9YUJb/3VugbQVIwGu9hXe
ustxiVlfPuEl7l4I+Tkp/BGuUgrE9EXuu+p0HMUSNPse/3d+eTpYHZrgTypLiIhRprOfh2b7y5t4
C57/xVKvpI/hEqe0e+DmhcSwh9RIZKA2MrjXPA8HvXIVFdsq54X/YhLU89nJseqrGpGRGtTEHqiK
GEgECPDX1UbzRjNYZBhPYWzNz8LsWlCGGyKHaQn7pwiEAh3lS+CPKhiQJPc4vf0r1/J36U6OaBIx
yEjgweC73/osnHpYVK/WZo/kiw5VJIpSywnERK+PS9BYF5UsDoDcJbGSAr9yIWNVt1423vKcX5aj
KpuE7maa4wWPQfTDuZzKqrAoQWNUzTwJVGA9jjAWlwdyeg+RYM9LcadWyahNGyucI01OFr4yEFQm
NDGXuqDgq9i9At6CTcaBdiwHbf027ZmgiLYMNm1PbxXwKvrIoDt8iI6z4CeO/HfwRXMw6vhbQaqG
bMUDIIfJ427/p+yYz/OKY75R9JC3n6u2LrSW2DYvcz6Sfna7lJjve8Oo1L/tvuc7mhe2Y3sfFwi/
CfhPQQqZCcsWq5nlhvFqz2sivpEltvmaeR58AbivVRzSoBJtl0QjCvWaR2lwHuoUXNAaxQTGBUEo
ww0UNUJuKHNQHEEyAUemCcxiU+KC1W6YCHj/XZi7PWmZnuwLdu8ZWnueQqoPH0qqsAZzPQTfmsJh
dTc+nZkSC/hMxXbgUB59q2hRNBg3tf2LkEli6QWJioTu4SjPXD1X24bev3BIAl2Vt5YtXcPt5ZsS
VNCNrXENDZaT1SbVUt/uo+tLMiuex61C1jiIAcbi9H21BZjtle1fTmWIOPbTQ4eIZ4esHRFl31Vu
gQ9sh2rBn9TVYeIshUmnQ0rYsz5YOtGMPH/G8aA2UW0FPJ7LE68Sgkb5sWYtk5VLUCF5cmZ82Ytn
2U5hc1+YPvQSkvi5Kh3cFFP9VrgmrDyxRQ8tRsG/LsNb0frtGR4rs1ipo6rpT1jbhBwOoB4T4G3b
NbUA8YTUZ1YXB+OvSSeTzapfwKzo0Aa0wtInPF3jslRy060L/gQNSRd5tqjDC5Ix6jvncjb4t46J
k7HsYbS7/bnkmk0IFV9oXnrlLAk7SXaWpnctgMI826sXMmCU/pMRtasyWTggVLnzZzYkmc7edg/w
TFiwlEmVaNjHtJEoxerTOpzrew471xAcicoCgUDcnsaU0LDsZptVEMZMgxKtiqrp3bARnJd5qfqs
VR7urh6dwcAwkbNCtNFF6eq5T4OLwYrvqPqukGF6hgm0ctsUE9ROGD0IvND99FhAbcOxbUIYnyso
O+zSxYjrj3DyRr0blI1KyKS41Kg0l3nht8/5SluRE+dj2VLiH0pvpEpt18GQaFZ+RZiANcUmleE0
OSFVG9l6UPnLwnZrMFL/jlRxmKZQMgdOiqGKXHfQSyXhj9ZS7LaGlS+mN8jC4iy9ePfxdJJSAPOh
l3sdxBAO3UH5h/bCFIwVmMMKjGlZRH5Bl2DC5cBqtZ4flrsVccWER1XbLNSof5CtmJu67ZRN2zI5
PTvBH98WXw090znfUyDv/XsiPt8NX3Jq+8VkiOdETW03KpcVO0A5ehSoBQOVC/oPTkjb1PmYUz14
z885HAktu305KFjnSR16ql1ctYDTAHq6kt2AEyw9Fdsi5Z0Yb1O9La+xp3ZUTPX+Ed5cFaOU0qqg
bt/f3IpEbesAtd+Kx/TB+jx330V+roj0rny77OKWwhl2z0+Qski7KrcXGAXSckrKjVHu5aVba59g
GeH/fi5Q1M9JUVsaRcB3JJ8kadENCKWEN47xzPONdGd5DVuQ2NXPJzk0o3tMZjdjX/EWOxKXbTMm
deo2yb+crDGAvg8yQlQOoT6tgO63nyIfnzoD/m+n5lJhcloafBqNZprQ65m5tx8sYfzMtIv7qNCF
JabtFWDst5c8aC6lFhkX4zJ1/HDBMSQgjTZSsfkh9Y137R0DnhuTupiG4WRbKyniFbriCxpkCqkj
h+QP3gNJtht2rBifBX5DkIejo/x9ee8gcYzOmWVnb75QMOi34DE7JbfbQz2GF81OQR1VbpVKFD5F
y0eMlIhPkR31uJflDCbofiD30Z+4mhaJ/+Xx1vJmHk2Z2Ba5shH+TsHMQpAPufL1m2F82uqVlGo5
P8eDDETdcLT4a6blZRb3/CTSdD9u64y74/vadaug3XsvHIcWD/8ebE4pdmX3koE67hg9b09eNLig
PoRq2/jjcppFmNxlq1vBIjv4vpovbez7/hzrZrteoTanKQejl3FUrsTaBPyXOYJ1nK7XpvcHY9ns
urtt7tBhljZDomakRGK/lHZKqH1wTRzz6ONl60NRIZ8sbMydBJLJ1nZ6MmGk4zzemC99sPsggHZ6
JIjClyHQFz8lk+bgTW9e4q0KxsVGF7vg44MIKlX4SAGXgi90QNXtFflZc38aCBcvZDKdTSVqJkNv
uhO8XMeDJ18IheSZLWFlXk+X9Lm1wURBtLBpeqpEWAeMiFor+2MQ5NDVlZpKhMV0Ts+VGHeBKjxV
n64cdvHONI1yy2/50eYmyoKf3GPA31JZ2DEM27rR7l7AKrbT5KEaGbSBJwV1+BNMkNpo6Nf50mOj
kSJhJDxLtdZQKoyNPIkHcBqfLcOcq+IwxG2S+bKe4qb51NZKvGrEf2pQzNknwmdvfGaDeP/fLphF
zBzuD4PnnQRSQHVTUqwsKMlvCHH+VGc8EwO33viT4rEZ9o+1meGmqfq5L2FvLStL/wNuUkW5sAaE
ngWZfBa3C+8noDe/eCu04JgM8i1ngcvMrjtiICHiU0WvfMPm9FKQsEn8A0jKMMMkVpnp9kKA/I+X
DD4yXwiqZWKxZOUhodoTx2IZ04+si9J25eFb3wfflJDDl0rY+vt7HTicBgKIaLFS1AqE2oYV70Vb
8LLO/q5kOfDa16NFU+0HdnI8C14jezZ8/GlrssQ7Hrrbf2QjgDqCmxcRU3qjAj6rCBSIrP6tuZkB
VFmDwMslnbo94ELsEeuWD2ZV04VAjV8Nwx4l9J45v33ncO/kJBYxASU5mYCVRjMxsp1rLGzhqvy9
ZfoAuLqQo8AI3aqhYHxP5mgMtq98scD657H0F8Djc3DEWb9eucoRFfBO4cL2yC3HIvK27+RfZz/F
gx57Y/9eVWsC+SK2QbSMd7e3pxt3QOyCrrv0yO2Otl5eLy117DfEg7N0Twvzjs5gUrFQmh2B4/s7
N6Soeo4ghGHruJtndvv/KfHl2C/b2HeoIQSNJx59q64A1UuKAoltuHO7uxRngptLWDxomNNplAMk
NhEfRJR2+81LyN0nfCqTxoj5MU9Dg5ic872YQUH8WR2QxYp1hesmexoB4aHEg/F/4tCamymhGOyy
csOJJ46dF3OcIV2y/8QV5+FxPMrfu3fQw1n9RuaJoNc94ANnNIzYqn8GFE2sZnrHGGKUtSKfVFeL
d0mNdM8tEmpmj+HUv8Jq5b8XyHvXIOZvG135n5ZuS7rtwrrVjkA/l1/tq1adrI3X5I1xNW/PnNXF
+qzc3Fvg+AiVN5j18kqGl9PVOlTTMdUK9pwVwnbnN4RFMgdfQdjsYVMBWkPa5tlOVZ51XqZ1pvSQ
390kWGcpZR3qaSm255YPF4FnPiiuvU7EiUtAx7/AXgnVb+iCgaE0vy/2om68Ya2iMrctmYxaEsb1
3NfPhgNsMPcoUzKQsq4daMR2s8nFWuULV/zswSg7qPE1guHcs+5bB3NIse/iT7L3TaHBmnV3aC6c
s8wWPmc1BN3CFpp4amlM5TzE+y60nfvdP5jfMFwn8v3yMucvPwGt+8VEnuwITxgCXRZsDj9/7096
QDjL4wpms/VKwQXJ9VhEeNaP+d88INN7J2IVmH/P/3o3+GirY7zVPE129+p3/KYOAZu8Z3ZgBfPc
HWqEWoiTrN5qI91d7DAugNwqlkmtxcGUWdF8lq82uPslH8OCBlJlLmgOLPnPImfb7gZsG/VNT5dM
vwWKo2cTY7hUqSLCnco3Qj8FSfUH2HZMsNGq6u5IcuFmiq3bPaL2VEV4MHuz72STRuc0Lu+BNEtg
zGqwiOGskyvdo+3ipYqSVRHZY+7zksJrXHl0d7GGWHAvZrvw2leVfR8Aojo9Wf82O9rhjIjqQxeQ
s0XcQGMG/b7C/Zc4YhGAnQJKft+LCbj1hH3NWcY/6UYUUIY/s2qcDq/mmyXHEjHAOAM967bJSEdf
7+S7DI53y1zc5WKTYIUG2/TMmZsdMeVhwPXy3aCKbgbiZq2c26RIjX/bzdIkrLoilWHg24C/O81U
j/j6r6pS+OL9o2Q7d4alUv8shQLNYzmLUaTTsKIbM8W3VMLJ6Fv7sIq4PeZNpO5jezUGwqkTcpVP
2+tpCFKEuLGySFtahMOtNVoeJMvTVBw+DktscwJ2K5mL8UHe/i1WgwoKk5kBbu9RIbYZ/5tH7Iig
+PFr+Qf3eKLNmVlso8VSX8BgaexKLnfRzKfCzg1l6oMk1W9WTCm9TxbVq/MOcJKXC0DmP8BPSL3z
geQueVktReGhZ4XZ10sNc8V4blMjNWGNcBtTQTwpHnH0DQHD3XVgnY7s9kgLfQg5GCLGtg1jcpJ8
SiVJ42h+Kw7BtQ+RM6Si6yrH4wfKF15cI6WXHbGQ6BCDuYvB8wERqym9J4y5GLI0gsBV2KirU+IV
7ZlKllg6Uli0BL5dPJnmZSqyxrIG8EwnQbRyj9RZPhPi0WCam+0nX4d9HVD1JuNH20f7dAQLeblM
uO6dB5a5cwZdi5G571OTvwao0vsofOGxCbIojC1k27lqtj2nMF3xz57mkBUbAyQmFvtH8xDpV74J
4aZo6f7ZWH/tDs9zSE5rGxGjJzmSo43950/7CroBP6vV38bH5IBfXpqEVz1qvOQ9Srp/K2zQ7HgZ
iy/cqph0iyPqnW9wgvK+fE6etGZhtwdcxplzZp+vjXAlIz4R4+oYlMLB5beZ8iZKw+xtNXwbNFd/
kbURruy0OiL64yBwRWkS5cwKlFBn78oE5biAFN4nCTJDuONHHrs0NxfIvXcAbYg4UbsBzbIvognK
SDJX3yOXiFPGdkyTb6PmwfU0LVC46FvFNwKHv1S/ppVh98RFKcNZ/cnKelKqlxSwuCXnCFbsnKaG
cPrtYzNeaeHG6W6qfDvs2Of8BywTrvChbDmlfr5VMIG1hIQCkdEqO12jEzEpw7rnioiwgCdBpu7w
weWH4zaMGsvLwL6mConAsD2gh0tWXIBoMXZ6OBAtu/hOgxal4e+Vj+GoU3vfSbP/8+rru2uV00C9
XSYjIZl7x251uLL+9/slvX7fVFeRBEu5CI4TJ4n8opFlJrwQrOc2yhXH348W3h9gjgOFP+5uy1NX
WODxuExXhFD0HspSDF+Jimz6gHFAzFafYTdagXnpuhLxpQKtzl3+a0lAltX3gQOyEhdOA6QbCmnD
1RweeWNPn/E1mzgBgaaxPaDpjp8VbfYcn/C33Tq2wCxo/ENYik0ITUuxYdpgcb3jugyZ6UyxXJZj
Ze4A1o+GhmmHhaM+oPuOw/8xk02O82NwpqszV2ploqchGChV0N71B5zt8uuGzJdp8dZLDwpaJErM
/SuwRPI0mi0F0+uWXlBnr4qpGprM0J4CQSukRXYlTlIuiTW+RHGEDAvaO26X3WCi2/4Cgf/f57oU
NrIkYqw4atF/jaljCniRSHe+6a6jI4Ft2mcyhhUw880gjPPrtx4kXBOJgcEgAqgkh10Mov5whV04
QHdbyjKkfZ/kstr8Rciw1CEVj1y72tkLko0ZO3Dogiwsp/HkJJvnlq+7meDzds2/W1uu5DvixvYM
EJiCWQF1Uy2CiKp7Yl4HWWcZSfNPxVZ2lAnDTqr7qduiXtsfez2pm3kGxiZt7gVOBk6OrWJwSktn
iUvc0xaQiJUax6h+Wd6ezM3Lojz9IFiZ02KDN1OFLW5qi9pw7cQw1PitsTM5MOy7PWoUo4i+Py0c
3Ey3KGvLyUf2qbc9NYsjl+E10XxWzu1nI6x/+ZQdHK24nfCoQuf+leC1jWpWZ+4LbSgnpjXjG2XX
8o5IVlWtNw/z9cQo/vdr7QN17hTzzG4OzO3e3VmTGphfi54waBiWNkOHwwIfc7UWfF31qtZKfnO4
3ex3Z3tpxp9Mf7DjKYEAxLDjGvKbQJTi2IvYHqCrk51GDZy/yE1CMfATDsljgzhKER7dYnD+r002
FWM7m6R+OkWn5l+SivSKGjMEntbWKPnlbUipWddZIu0qt/ClN1GJyp1q7EK8dAubiUDxNLDKg0BO
j1MfKkBHQHYEnAvxAslu3fTmhbgZJLUqZ2SvKP6k7qJCImO32IgkPKmrlc1F/O7Kj78/JE6iPNjz
VVBHrnj96S8EDDcLg/jQL+Tu6qKsvTC4IFKT3J5P4TSS73AH2bpbXISL4Q3xyw/3/YTfiKN2Xm7a
vlbWn8leHpo5j/nwr7Q8VQoPLYf0d5VBg9y9Sfx1Bz3f9uq/rf93nk5T1w5PRpYHq1DCgQg4BXy7
PmEJ7m7CWn5jEEhDzarl/hUZ9j6T7EDPa93jz+ur8xq72r/4x2T1Gh4RmXjVCq6hPCFDVZHGCmwA
4LYQxC+yJk42/oRnzkInAADMJy3bGOkknU7IrqbT4L42UeGOAJ7EkHWUB03utfulTsrcBNxAb/mb
QNseDpbewsbgqXz1HjiPVhzuws0r/K47TBvlodHZxAAm9LvHTadx4+9VVfGCD2jEo9+cwkDB6MQd
3PbUWpujZc1gwMq2wWPD3Om53xU4uBPW05lDAX8ci/bmD9gXNzTGHTbErHn6rvLx4FnT2Zs4ezLz
81O6+7Qwekin5ocO6guk4ItR/jIyG36sJrCsqNvDdRfO5BlwfEzOgEYP0u7ACC+WapK1gcYImzwh
an+kPVR71mJU68rPtX/BUL3y65wLgTay3f643RWR8+UAL39PVyF7vIFRaIs117yZhnE4fb/p3hCi
0tq2bL9MOTt1Z1Twr9g5rVtK0pKy+7kVgpPOAwwV0t6PSjQ/E0kkKazILkH6vhU+Y8Z/9FQ8+e2q
u8EyORQ3KA7TfkUhsRxLOEzL54bjPuXPbM/OLnasp5hgY6BgRGNiNV0uX0lzmS6YZOs3ply7TqBP
ZhZYXrJ+j+KzH0kDe/3HZAHDS0f6PO8G7hQMAA5WQcJQ4vVFNltA5VEVE85dHvSbo7qi9PUE+Sy/
p2C7ME8Bow3m37Dd53W/aTffkOFKjDvDWqmxLyDBYd0WmDjFIoC27cTAY45uNLs0mjVxmFnjhoqM
7VhWcyhYmAVyFPszGvCEPjKftsNiLHMPlXPqJIlJCLHHKVCVXuCjMi/u+yqur2AuJUQmFab21Kd8
BmmWHzPrv3gCfMtbj97nymAI6kvbez03GXhVRq5+hhl126SeumHFvTMLVbDK4ChR5bbFm5ZdN3Lg
SNkJI1x1RxOjRz9zsH4CvT42ZIC3TSy8DWiTDq2Bp1ikmHUkMVlG3lKfIJitbJR08bijCiul0yJJ
dakelFGJEntua+knaobm5ZJdiiP/609KJxvbsgPBpAdlp33r136CCcpaXEEx0/bvHgfPL42OrWpk
a9s2RHFWzkxD2m085ocoWbW57wPDdCUy6d9VWp1tXKhx/7TsH/VcHnEzh57WxRlux4tCbKx+IOJl
rTt9l8Av84UY8fiGxvBSm6mOT/RAqvhQbqYFjEhyE+R6soXUNApa8G2GonvNMrZyBQPK4V00XqR3
jynKqc3Qke5TRyzJ5DwjNSCgOPB3f18OxhInbsLZWNq6SdAtHGyNa4DM8EafldME1z+cZxAnXWUD
6KA7kraLftktezsIXPR+4oudaOA4xM4cJdvnmuYwQ2MfeOO2RTcheGwn9yt4q3Fci1DYKnL6FFVM
vh8DmUW6HXYAhwJc/f0eo6Z74kGqIunma5qkXuO/NQ2JM/HUU0PX4R7LM6k8eH2rDMbnRCMk2cU5
v7vAG4AbotwF/AIbxxW8kA20wYseBwkuGINoJaCr9p8Gwyut7TrZDXYbojDtZHY9WcxJm6N6oC2e
6JmczAm7sHDqIkRHCUh/PG72C0ojHUHk3CGuIupY8fZ+jynSvZAyF8NO+upOIQluUBp/MczAxSq6
4KIfGhFWCZc5FUwOvSI6rYYeZZow4d7DGNrUukG5qiKNPzBly4YH66Ut7wrK7moSd9xTM6aLTHF9
+JHCktvmo9CrKM4DMGgg2wse9LoA8gnEV8ZdPku9h2r31rzYNoRADHvAhnWNXpeXwsXRCrRtSDdX
Ept4nbWnT2Ec02cvCRVivsvqHQe0IoS75mrs5/B78Wy7LPeMg+I+g+E3YN3BDSzHP1yMoIeVfFT9
I0mZcnsIKIokNZprhravBqFC7LY4c0QfVt/j9sJfFFvHMD38f0owgKY+xOXnk0W6R0t/VJEU32nF
BxxrLVt4etQD/86DCUtflfQc8UJ0Vej0bClu8v6HDhp3wM1rdOks4oawWdVDZgMQ6LO0WRXA/JLj
GTIT1+t5uCrX096owLl5D2SUTLyDUiltV1Rfsp8MTonSJ4qfKl32dyc4XQoKDETEl2y+64xP4cwj
LMR6Njzj+pkZGKrqQO9LmnZYyUoRzb++pEjOvShnsZ9VP+HGvljia+fKTOcPMG8wpuG37ULAHVUh
/fnNAMPaN7BajOFJbQUUIjE/v3cmByZaccg9qpr2oNf1Do6DkkxAWzm72ElQQDJzV01M+ZY7LCOC
TkcaFT7NeaaM7fIvaawjIqBtOC6GqM/UZ0iwHNwOTAo5vOF/CPX1/WznlhsppPVJNFIb2DnKKDzi
u13B8PT2OEo2YMH4ZOREoFMZsQ61/fBi40/b8tYLMoNisomGMAhBUGQEEOsp4fvMgY/wGPAi8SUZ
zguPFqlYhrOQjFCNnZqgMp/gjlnJJNjvLGRfTBzFOsMGQnt+6miaVryczC98k7FjnAEtNGLn2VDF
lwEIfo7otZ+MaAR9lkkkiCwn1JfPcRK22Ea5rJ4BCfHiwLBCYvl7/c2RbpeWAj0+XDYJnuf+CnAh
yRaixVdADm6iNWQtsknQ5CAd/tNjSadWSskgxVUpOpYlqRK0kOIUXutZeTbjan7R4jyRmNjDJKrI
qyU/o0ozKD3r9QYlEAaaHJtrSEP3BkvLZWUibAeCDa1qI6A/YQeLA8pDnpS4ntAht/PA+zJ0L1c2
GwDf3bUo7pJZIU8E8NHG8cjW9UWumeND1WbMvJtKuA8wlQ9UsEgMpBlXYwZlEPzaNx7dGkXU4DDZ
KRWkH9Jqd8mBV+mQAvBynHcDrXJJzjlxwqr6rG81epSlHuJ6ohlwZZJZ9DTWJd5je9WywYij8QSL
IX82X5SU9LOZnlLus3fYCoTxaNm80xsEeAqaBjWiscKL5lvXlSikU5TsosTPYBXUVl1cjHr/t0mm
96zTu5N80Lgbk055j0lvBm4RpvNazQTxlnp6kESJZZaIk3syF1HLQCqXz4OqNRDtvVybEqtr4gUb
Db8J8CVbshpDhHsAKiBEJkqBm3rFQ+DXP8XkrHhM2Nx8X5S26e4KTgOxIaglyp5Lhhz/jYE/XGYz
eq3UeWkUVwYsXFOqoemmn/59lG/WARkT7EBtKwdqmKeQ4U09mdfFC87dxvQ4zr2+mi85QyOpkC1/
NzKY/t3wY58d4oL/yc9dk73bdh4tnePIY031DP9v4F4R2gnjc8UxFZj+tLwtZ4BTwQLqa7ciikWO
FJ8DMgn8CwuTXJmM0F8j6kR27hUy3qyHMhevM/vHWF66iGke8mrrOuknk8Ts21iygPPV2+RhNkEv
rFzGfu9+e1lbwnxo83NVf0cg8y/PRepnaIyqHiLoHG1vk0CpwHRHtpfHro1Qt3biDcdffA1Hkyq3
F1jpVQf7Wy+62Mc325t0XOIuMbdUODkGC/X5NmsqkXtU30qRzi6hjjjfdEUEqCDJLute9B1ECPVK
qh9r5lB7Xwh/gp8CVQNvrB9cMaZxr/Lu06mIxAscI357DFCJ7ioMtTYjwT91YgwZQvx95ePYFFkK
d4+lDqwu9acA6ozGch2YeeQukgTP4kAosohlg4RoYO4jpw9wa/CWxeHzaVpQFmT1WgWAMgSDWsNP
FDNpWRzyFRtnC/kxA1p05KYLhm1sPMcazH4ZN+1yDVWngR8VST8fReHEz7sX7w33f16XmzJdpyES
SL0rwtkl8ObCWnL/LDhCy3Yxosr/moVlGwztLyILashooyYomkt3Qnm/WrkRe7XSo/iHfUnmwOtU
dpDtY+hfD93psOxZlDMgv4/p91Yxc/ryRaAisrPvPYTDgCfpXqWNrexcTjEIQl9SjEBmQ8uFkU92
P0Mwf/v08rBGHoHUfdo863TG8INqQoQ+9ZB+NP9Zx4CCHFG+0rKjHkkLntHZ0+tXBMJsP1uTqgnK
dCm+y4SAu6TKGIHSHB9AdYaNE54MRsdrIUhevDKLL6Vev/6J1AiOcZC900fRg9JMJtzU8Miscpk6
t6F7VGRMvE2CrcCBpCvwyG4/r9wmsXoBs6YDvt+qpg+R/dukXywfRudxQhRRlxt9B3RY7SAnk/20
rjMaM4Cejnp0ImHGCwo6Y1e1i+WqJLwuWc6C3XrY7gkLmExN5Zitn4wyKESa4VIamWFZehpz6nsT
cIO492BGf7KUlzq729uaWeNl7W8ruKvbBsQDIbOSMg8DzCpUim6THUsDMT60drQs0JWp2uOw1Kh8
ycg/hR0Jd/Lsyrju/ID6g7dLinwm6V9w6uY2PHn6pEJPVL+oxKK7AFIQh1Qb4d2axL316gyuFyCh
fJf0zbZCoqRZOj5EgOlLA4A95UPE5MMARQqWzrR5gLfPgE/E1FsE17f8xaUe3tkhBoKs7kvlNQWM
qRl5Yf1yv/zBF2WH76f/5sVxoyVTM/458Kam5Fc/MJHUXCW1yf6ZqlnPjWX8/SijemjIz3ea4XS/
X2phdnSqrJt2KmkF+cOWnkCMshfA43YpRCjLG2p63+0GZSxh2m4F1v98DBByC+XV2P2ZoG4Jcp+P
vbkLu70e82MW27ejZCPRO2FS0INwBNS64QK7lpL+pMXiPb2VVprk+r3qN/LOZJX+Cf+SM6Ji6hyU
gbNn549VZRT2NtuzMP0eQMMrOckXEzQ0zBk0J9PJm5JKsHoP13UuXGYuQcCEuvpUt7Yn7k9TbpgC
ZqcHvwGB9n4FeWSWQBpNLcxO9APhpKjNJI+6aL1D379i66Tm4VAFv4ViyKK/bDGbnlPsyY6BYjJK
NwVyWuZzoYysPxoUuGmmAx1/s9Qmt5VVLACoN4um4MiCdA4blVkESu6LtE5VTjxCZ/9i1OHuKEui
I29Yc7TRBsoRjon+LTAyOFJOCU8o8YFHrdAfzZnNISovu9fiLO9OZ7zrOF8SfqN4bnIM7BlOdoZu
Xwo8QRY2JZIIcQGdr5bln/faqbWVc+SqhLGyQrgrtcu5HJJ3fmgWbW2YvsmhP6il5j67xqFpItvu
c5PwBiL32zyJEhiFump8ua4epqFl1x+1FjhH3D8PudOYQ47aKajBl2R27SFMXnBgpnYjJTylEtZF
T6FAlsE4lm31uVeOtJ+nYH8/TFIm28wQIQSkGAmOH7HDzBuGQkhRKIq6P/wavDVDdh1aadHrlObK
FdgywwkMrTFzdxNHWbW/TqqRLcKC/zX4N8toqx+hdTyj+riUb/9fjcGX/BGoDTdH5BNU6cfUw+Uz
Oew6toERjCJw5WalCQJSExqPA6xad4SQ9HGbh3d/nePK9Gj5uiVOA+NQTqXa7jvJRNzs9qtUDV9f
sGNtOJF3w4bDG6WMT21bH9wKt4LDtz8CqspFQynUxhCg0ozaYFNQgQZquncyv8Tf/5Otj+cb3IKN
5CVUPtSFLDaKKOggAi3iDJTtIerT7RFk/OhRTa+gldO5yVWSb8bDIelnFiFxO9nSta3Hl8hzp3yD
7zp9fvuTXX18HwXNvlsadPW1RJPZRrWWDoqdWrkc4QJT4ZAylfV8b7bu1lvfTgIqfAHQqajrNkbE
X3C33J02uwTTp4gPHA6s0wTX+lcAIt5w6PjuZiGnIgAqzyXD7/C55hZKAZir2nPax8f7CDhhm5zD
fIFV9zJ++cki5Gd+eeGIMY0UI62V+gUIJzzVnjM9slBcHlzHy1XARXVpDRich2rJD5lvxuVg70/c
Me9nitUPevt2q8SMq3lg+hG3Ie2AuGe/dSqQXQ9DWqWZprEJ19tYttnosaKdxDw5w+YKDL8ypEJF
G/BohhdkW22IZsD/26gDaJ61dOF1CXomZAF4tuUdoh8/upFTvVyYDHusPZReHryxP7D3+N5QQOc7
Vq+xM7FbsdHYENgmGStVzZkYVylOnz8KYQ4vA0prfPOInrF1vyrPBL1nbbnyqjTa9n+GLgvrfmtv
h7+CWDTNqfGAKLKdoKnpCiTyNTeEfyNchrlqnOcRKyKGCfcqDg0KDuo5iwWmsqNyeL486cvU7XGp
58eLCsjK046FWkMVzH04LHngVNPrVM7Gbj0vgp/uAyZ5ImJksgVmASfJ17OGLvdAdCXmcIB3nWWe
p3/JjgRoEUWEDT1G4PwnvCnEe897gKhJIUpSnrHzNrKAQ/pSADemk8BUcjVNWXSLxpymMe2bfoUT
tYtgNifc5FRBoNHHGhigIT+zdsJx1pKMhk+2H4ZxTPkGZo4tollsYt4sEVcHrEz1cK5Vs15iqJTa
MWUfNU8xTOjNAgnAKzkoXXxQdSNnSD3lIeHKoRTYE1kKYZGXlkoXJ0bV341bBCW/IIiA5GDjwUaT
eG90LjAW8NtXzH0eJX8QHVQG3+bv4w7bd2GRQaWc3x7Cz8JhgneysbL56lzClxx9Q8qUOFQ4iLAd
PgI8MplVg02PkShruEsOI3IcaS5PXZDiEti8kX6bcy1jDePSrnC6BQsGVf/6wn6OyCJmwnCjQ4aI
/zHiofmUsYDjbHvVcif5SKOj9SvRq9ACRryBv/+Rh4gyfmfHjVDGBNjTzeTlW0i+uAjY2yHTBCfw
3AEn/x/MBk4+S6glUpM6/ZDOradn6nlI5ILeuw4Cunjg3r1qqDViUktTNiXPtUmoiZtnhNHCevM9
+R4MsjjVF5c1LBD/pu6ZlJWhtCKCpW894MFvVUcAuaW7mGBqbV1LLGDDtHoaO6OJXnPThhn4H6MZ
h3EMbKGu5y+zbAIvZ8MT1V/iowLqO3MBOYG6db9QHGwibaQ6lAy4EVAXWE/rIFvedARLw/yVb++/
kl3bWuVd+GccU2e7uaJ/zgg+lbym5MbA9+FbJmRGoCLZEsufPkE2rVQPbRb7L+vlxxapRxNWPcVD
AwOxcjKie8fl48nrLvw30O1wxx9+Qh5uxZZO3//bLZwptWyw2qa1mg6LO+9Oaq+QLwb98mF71o0W
GGW3jSwu6wlaxQYW3Xuk+v43RnU4fM3ec+bfEl0vxzT3iv/wbTjztQUwCk3ISa8GfyA3ATp3e7PH
cwrvdfSAAv3PYApbQjKwU+nm3Gk8gNmxudYLMHplEXnZ8nq4hSihuzkS8mPEoO/YEc9TRF4cJl0f
GiYGLTHKHTxSsGDv4qXn9kmCs14DTdKFDWbh7FF3ITFNzoBeeMJ15qFapnhDr0ZepNY+QgI+KHh6
P3pP99wED1qgu7rGzeY1L2THmSEgwZha5TYrOdQLq+kmfwiJToTJy1bZP0kIu9+ehKVWnI5lew7f
swcc7qcINzs1Ofo1syZpXlDxJDRs8slElviHLIQu2SQAq/OgachCTXTOtP97JBl1IIcqPCYzwuX3
gn6P8ju1s5OSSKr6gWM9wyCU5j/HzDvj+pFEhJ608hpmAKHHCt4vbk7a2obHHG88UJy+qju+4NWT
IrCVN1HkU4/27cFnaZW+D8bux2b9D8DpvnLydaB1GvvcCnbnQxhjRrpe2vRuc/lHc4TxCQB5+oSh
vvh7yhiHzgIutwFKfFeQ+TUJZ6bSzeQwdQYPgtQM/0IkYIQfavWj+6ohCbEv1wCe3u1So8kp4K44
ubBqB1F+zGEaPLFMKiPT4buQTXeFOqUM4UdRQnuB2i9U41ckxIGceyFOObb8zEEFGsmt3LEo2G+r
LmUxWcnvDsxu+MGaTh327Ubb4hzz/9eLlNEFlNrvv6xo9m3H0MohOSybfY5YHfRPHDcWAKz69ZJJ
F8MSSp/rDt3XYtKkHApiAiLyVKzHFqNPoXrldTKEjXp22HFUxgmXEY95WGu0wrzqCoz93ROR8H4b
W0XEnoIVIZvlEjhGiUB29UFeBE5llsE+G8Kcw56mVEpAX2KocE6FZUh6q9Tb2U1+x2Vd4UGruEZG
5mQzGmmDIe/geKVJtAPwZiBg8SUnI7xAt0qe4XBMJjsSmRTFUXlaT4TGRZYWe2xk0jGbUV9UxXJQ
XFg4dHeQijxVLD6V/dUZBDPoLUxIP7e3bzOsUad6PBqSqP/XH/wLwUNS0msFmdIkOQb71zDQ2yC9
twgkyOV3XtN4cf8biq7m3UnJ1GEkCGsk8To8OozlU1sytfOMparqRQLFfmsNlzr5owd486VnhLZ5
qGyw6MICJg9JRuzww2SG64S17rTSP7Ffn5mpIQRG8xbMHOZAXs54X21YUYzkr4d0RYqk2pFz/Qsl
9bjdRoNquPZT4lJKQxZ6TZkxER01e1r0F0FuEg4LNFD7Iot1sOCSzXQqFumStzlJswsO0C8SGJ7o
ThI2UNnnideRENfcAu9UOzEJ9HvSK+o2JnjMZT2u8qA5enk5o0aa+niRakxRYbNOoFh0HXGmyuh9
/u+pi6wYBU9hzkac5jMCEzzE+G7/TD7UVfjbKKicge4ZyV17FHS6iK+aw+Z9C1QUTGWLpGAPJ097
GjhL7iV1QlHxdzNEQg6BiaLQtAtp9n4SjIiTlnHesJTF1mnztHo+uzBFD10iz9OReDlkR9NqSSgk
M++MZaPMCiQyQVAxNCwY85FB2tmVNp2HZ56o5lRn78nFv1JdaVTt0nkukBrujnBgXAhLS4lvF8eT
4BVR/UerLrSEDm4c4N1n6FXJSIjUWT7LfNuRLI9scMR7IioZl7rOXRy+BU9s3bXL4TTddvbfJCJ6
LD4XP+L8KPuAFWFUPx+MsqDZBJ+56vZCV2dGvSl26fuW7drKBqG6QArpJXbh49BJjjfUlXn8+Hyl
fgl4oXXfwYpnFoADcFDhaQK92lVrzpIhQXj1L3MN53Jwl4bTjcvP/df3ROg5vu0fs7uyUrdKZkay
fg2neSxCQEo8zBdyf9Ev0+7pMxEto6gFOTHlQPvab2aw6bLvHjsarzKGaWnlWX89BTMdse7Ayy5s
SVB5OLx7pn1Dnln2iqpNk4FjH79D6KarfoyMAqYhQ7/x9am21Hna6Tra16+x7z0je8eCerVlgMUR
aFZwvhTh+MBUqj9b7C29m5h4zAeY59unKRxZkVBN76XJkq3NtYucqhNH37GqYABRR1nIHY04PeIg
24JjUXpMO9NDkzIR3zGf+YpCt0j0XAQ4TggcTq9NUWg0vf16WhmYZ7MbP3hzBTT74/Mg/XBV51Z0
vTcciQ0mG4Z4BQUl3dwQQZ7Scrzu4OwSnKoqhPK8yecV46vjsO0OBWTvNoqm7603JmlSupbYIjJS
KNtm2auROS7om0ItAHqWK4FTs9ogordGW8Fm4f/zzv6B1Ko7EudTxywDtSh7veLbiiM+dbzi4bi2
L7BOd7KPLYXjvGNs9byNQq6xrLdtClIEOaw9FSOy+vwIb9deHAoFqT7NVlYNumR7mQX2j1dOlRLG
eIqufaQB73al4EnLiLql5texbmwab6DdNM6nKpfwYz3m16WBEJzxisG+5F4jz+cXFV6gzG0GGqNm
1T84m6EZP6zE4cmrBz3F9QBimgfpppCvnSQgnYckukyhw9bKr5EFQOfTNIGTpw7RBjgjZt0wEneg
q24MjWNI2uh6fUtaWR8qSjtuSeB62fU1G5TXM2VwvTov7ThCH0X7taFo+PzzjzYtIh17t92oR0g2
iqTe/j8Z7AfLuEm/YDkvSFgNWIS2LoSdbbEtafb0cDIK8A23oy9QwYbIrSFo4Gh2aJ9dXxQOiyJl
6ctnrnwwGFiTkUNhfL81qqULlTPv6zXT4dyRifY56WzATGgXfIdjAH9ZvYb/35oEQ12nR4CXYjSI
QI8+qviyXeDgCjaxQvJuLJQqDcPLED2tlfFjcguyj9Cc0zQp4jbz81yHmTx8tPzNbL8l+IpHCjpT
n2xKsjoL9FcCdFbvJWvJ6YyK5MlPBpNRlXYV3+GzY/x0CjMskbBCizCi1aiRDxwfA6qaPPQxO9xX
9YdpUNrUQWlMSy0xV53MSCZzK5S68LqSNYCwVVBYdqFtUgPLEYWg75VgNppf2B+VQbT4r3TXm+E8
N8XfzRAg7MkCs2OwqFnBAIxOZloIYDok9fE6eY8gP/OLWgGl5Pu68+3ebaXZb470MgHiAG/3wyNK
6/XdB6Z7vy8pcVTci9pAfgFX3GoSO4DWhai1Tp/eQS9nY+Gw+aLk37gDudbE0HE2wXRqSiUcqP9q
jsu5Ab+h0fL27s8aZQrFmi3TWc3ZjR6+BMf2BhO/ECI/NGoukPBKol2Yxe2pWsz12bVJVP5knZV6
XfOOyxwWfcT1iolQEAj9vXVhbCFkCK4clJNh6BybGFzykfl+LVJ9GYRqvzUDEYbQ4mXQrzMBuuHS
YufWo+dD8jhbjrboPNpmPWGWG7E9GGwbKIh3ZSatqYSWK4UlqSYDG1Oqq6FF8kOAu9CLSb6jKgpf
mOoQrv/VCi2avUfZP+CSuda1TZ58jIYpPsGLnwcT11oOTcc7aT2wBeZerZ1pcf7qQ8glDNB+ATQL
l6abMmMNQ4Z8ZRfWmGT8WIoe/eGAgNJos9steni4njcVmUgkEC5IS6X6iOlfcPOJndce0jXkN2g3
AQuCcohbiiGjegvGoN5Lb/skRyez0Xklem/e4aR84oLLnHFNqjii/jLZSC5ue4Mukit9ZWknh98H
mzMFfBsQGYidrDL7K9v5COTVRapoUPWuKBi5anGtVbFK18g9ZAkR4DGQdithA8qwWWNHSKlaQSaP
K6pw+p5RD9Te4DYahGUgTyBudMfIdh1JAkUJ1miYA8zGLzKXiZhXVXpomlQWSSanp+sMclCMf9X6
zRqPbKZbwoysLPVXDFZxFb4PZgbyJEVbJFCALc5jqhC5f0PKyt7Yc3QVFxYeQTwSVUjKT1IydrSj
MPNIDLe+wCbpM4olhjv8FxZwxXq3Wb9SQB/rAvYREfdUK1l7rYoAG6qDEV3asWQqucYriB1YcrFw
gKRUxNpW1MaRvvwhpdsmNpg3JLaMmr/upvhM3SAZkDOBqYa+qcY2xoh4EuDahHGwmEMLFoQYEvqP
lxGVcJwa2MQ8YIXgTGdI7pjv4g4BrJSKdZYoliwA+zaj+UULjSyS8l5ODDrUTFB3WQRU0VD9Q1r1
sJQKuoqGwWgkXUnSYdImKKoRPeVD2Sd2KnLPqYKY9gmxs9SYFqvhxw4Q67hWrUo2gsZqJwqT4jdD
5U8vmdQVsP7HCHq8Jb5XuwM9RmSNs7/WnQ5YZDX+O/a81ThbcZXRkrKVGclu7EXNSZ+xXLfv2qc+
Vi4bF8HOvNfmEyEJXrmVTGFDZoW4WKrUbF5UGFAw7/K5xq9uUoBX1Xsajn2qO4V7yuyHFt/8TOy5
7/+aXPQoN04/3fhCu4Ej5onRWbyxJ5fyKDIdcBcJXHMtcWvf4mH/Kgm17A6M7Lvs+B/nGOlTFoJ9
2FJ2i4bBPse8VlaYV3stCslGD4PmCbpXJDzMxKPdSRDvK33R7UeJjr33Knffqs7y1OuSzknvp3Op
QXbuh2MsI6OZtVo0OAnZFn3UM5rCf3EjGKcuXJdzwB1DEENYjU9Wt1lMAZkJ4ZorqSpLxGf+UMOn
EWeagAefmcYBiDj+d1g+/w32KqG3etzhvr6us3RX+WSNZBKyqYf1LmY/wFkAYCuR1kRk5qw6zt9u
x46rh1+u9yvk3JL37FhMlpixU2QAg41UU4VIQleLLkxqzt4NxWCOvd7rkAAY4+NsO1sgVFpBkDuw
Um1+9EhE7RpPV0swW1YUxEBiUaC0RH/2irdv1lVsurZ5RQ+goXb638g8vJtK6gLfWMogLVraCVxf
1o7VNHf1Zb+VTFeWlJRE0wZrw96FGkCH2GxBzQvHH9bgASXhm0TS/NRNconvSyr4bC0qVc/UIuSU
2A0B31mLMRnKDVEJiDMLMFnzTISxqtBHb2YtoNteXkxzWuHnwZw2To1edCIdpo+EStTYQNR9osRq
sDPFUTe8yxq5kl1OWrgf1NlTAfqYECrdu9kjSuE0COrLCavGyssc6Io+g64sRHHef7bidHdCYj9Z
P3qknEfRQOUa5v4ockPLtHsSQU6mGD1oQBjvqYSzS4I4QVYIU+6m4bnXiayPd2EtXwDytNCcwND5
KxnzkXBvaLFd4Mdzd96edZiEKyCrl71xg5qlnbIZHCEYxZj0GNK/UVZF+xgEuUzcTK59VNRELx2v
0sVHWbWjDDgUVFutMDYrybA7QdiMkixmwpv7T75bZDLQvqKnJp3mSSeZirSea74FXIeogyVqc2Ho
OlF8m8UkIZTy5eqLQ046YtBOxYxYi7FKyDIYSoiGC3QrMXj9/C2XyQVyHPUNLkcqTvjWiOXYBK0Y
8Ziv70a9bopsP+f1lXZjPG0N2E1AeSiwlxAIubKMs2eMJczKNcqkb7Len6ROEKaPyrH87vZ3+rWg
Q0GRZ5hyeRMVycZMxjcWll+9FS0KykyPvIlMxcXNb757ln3Ud6rlDlwSvZD07ezW2Nw8mGa/Yr/w
1uz4BNmGyWQf+Wm37eHaifpVCFSpZFxl2m7K/lOCnabZDsrU5AflvuTJ9QVG14ZK5Y4sJKRuWy/E
nEOyt5OoEbVS9XyXgpTY1vZUHVUrXvOPEpqRwe6KN1S8GoiXKD79glmo9knpWJwiLPakvj+ywDPo
6sL4jG//B19wA4cBPDVVpwg/zed6/uhKPAHJK3VFZ9rwgSD6MaZ7TZ8w8zFnsQtztVhwdt3Hh3fc
vpkvtgp0pv7wCRYCIPX5WyhS8Q2gWd5W4tUDIFr7edB+8ikjGmVFBMM1HSSWm4EJJ0r/mmdsHwdw
j7xBiovlRrF+lB4nhUeoY2JJkd+RtH8ES00GBaG7h0YHgWdxh6BTrPuVdrrl8Uo15MwjjPq29DAg
CnWhfiYKQBDuJbJECKlBOjSbPW2sHJwyQRb9po6reMZy7SCJkv8mBB1enLeAq8Ffzc2oQwWeEXdi
yR91j5La/NYR2y0ee7tSiDUBb7nBCPVe1qk7UMQ8GbW4DgmtUiedxfb71eGrzpkKRoz8CeK/067y
JtIYc1x0Lbfnur05veQkprHzpvg10LS+YP+R7VOfUPYSsALcTfYSLgZ6M7fR28us4IyZT+bPzCnP
Go0kz7u6I9dQun04LkWg2ZJ0lZmkVXUtC1qeQP/mUXnlq9Q3h0EswK5xuk74JuG+Ts5pWihNfaZS
/NNlSov7aSc1vJzHZex+PTXnjkVVMlkd9dBMNmt0sisYiIYOxU87p/FWE3kuvXgfu7l/QxKfb+Pm
g5+b21lEerVPVFyVIn0QlHwYPNncKAcBZtJRHk8RNaUtFhL0ZMrt5Kc+egYmzfbROrVubfTrSH4L
i2KI0BkV8nwFN2kaO1TzXHwUu3uDRJ376hDYA9Emtmk19rcyDkSRB5u5i0haeJgVW/28a1SaORZj
f3UCbRwS7ZIOWcZlNsYttgizKruDjr9IVAfC7p6mrKGBxw2oVhLYR41sDxMEKwkVjl68RM4zirDu
qbcxFMODiGrk+wUtgyPtkCBXDgc826ebelmXUD1aH5kBUwD2eIKv61+j8kL6t2Zd3Vu54QNyU+CI
ILRJ40t6Np5z9Y7MHjL8YlO6L/R1j9Je/ud894nPgVu0MhRVjb6OGJTPLGni7vWUq9SS8QmvBsja
Y7d8m00Ml2PURTRJyyhnX/YLoPZAifWnznBZY6/uTKXrUXljA/LRccGxm4m8KAvtZ/KkanDNMXaK
8EJUNRGuqtRY373jlkuP7ERk0IFhkt2jK22ueYdPcI7bu1byo4AeS9SfRa68Jhbculef3ZF81r5j
YJPDxhG1sD8tLLtoTQ0GzvaKm//upSnm/9ipynq8fD2FUYewsdz2mqOEVu/8TFNCuWvKz1qOXCzo
+h0VIcm+vsHBZvU3A3EUI8pyiRxGcdbBIQZtsV4TAe6d1LB2kwe2ahW80bGpB1tZPWmBIcwloG2c
AgZTGaJnQWxa9cgPz7wLga6M3+wThv3k+rgmVOEISNgwXZnuc12ZM1ViiPXGqBJ3tZY6urr9YA4R
G5Kad0FFM8WzzuBt+l9RrrQskDGxAzV0Df9EpQaafvg4/dHqqxg58rktMiD/xHHrWUT0htZO7ACP
KAX8x7FZAo1sjKYdp7D90bh+jVPUQr+zyh0PFU2k1eYRzFiFnok6ceCzguOepvPeuSGtQPMOqCUI
v5OoXm6cNGDjyoDDfRvP9AhW/iOwEfvPzGmRR1xrfLSHBSIuYvtYH1jWwCThXEJI+9axJPA33fRj
QZgD224OH+LIsS3N7Mk9Wf9ih+/4dYCLloAY3lnfWW8G6WYc+ATv94aMBAPztKHbsqPzPLH7hZM1
tjlrDNEmMtuh6g7jHCgADMnDfmNjghL/P3p43NMGcVATcRFD5VEHRxBYZvZDD2Kj0UcSd2su9iBP
zhZ6zgopZnXvhi+M5xDblqCgyurgBqOLt0d0ZApY5tUXrml8I7d1oC5bsz038Jh4+l1AnhbaI6zD
6OA/4XEGDPbHLz+lxUt5HG1sstQudpHTFC7nWcIAHpE9BaVIi/avD0UZEMZqS/ikDZ9gm+Cae3AT
R78lTuafBuROdxlY4Dy/kVcNCMgxzM/swN13UDatA4o7ibEcXgXIC7EyF/eTDRWHJeJCd6iKWWSo
KVGUklQA5ILKDCYkww2J587jVbEBVNDSN/GVW1HnX2el7e/1W8fldrCos1tkeD4eCLim+YLD+Y9r
Rzh+b6J4jWM+ru1JY3uPV9OBYlgSiWSFlGSBLQ6sH4nY3C+AIp2xN318NqgNV/vUWSph0KkAezaF
BWRQZD1s/S2QLqPWgGgxcvPkLK0L9rBaurUA4vhC8sFUMLkMOmpXf8MrM7Hxj3TbboaJ6NenQyzQ
QaVQCsRGFxaLVdW3yVzJ6kDpjzrbZqIFfPWlk34NSPomx3F3gaCEhmED5aVmnwP7/Usl7wi1/mS3
PJYiJl+IjHYjmI2sGPZFkRs2GT1BaZf5Kzy+NWJltAJYT2G7TSFJXedCc2vafUBIp7w56TfCCXUQ
fLGiv4BNG/a7Lm5FmLpkdFXpmw9yh4S5GIj5K2v/xeX41RB21Ufq6s7QZVUHSVHyFG0EL+DL7Yk6
7o1LhhnGXBVZMDVb0pUo/LNQ1wl+T+DgXP7o8SBhRsMDaz/0NQYp6+pNbJA8CIxuEda1xI7xVHPT
sS/D6+X9VpTtuOT7gq6MAZJPU14vrMlMdM29WbXddBFB2HYp6oSv7Wmovrjb0yg1Ujn6qKA/ggUr
e/JZb+38BUprePO+vWxRuuuJa9zoL9iQF7mdz3MhBlZyYg5q+E6o7E7H+YfZwPzNcZJKaUGBiFjV
tEmmKbdsj77XxXeGkwco4D7HmTdUhnALIwI3aTkujJguW6TBItmePIcM4zLUVOj1NLHCnMbKY1HJ
QnfyZycpNk/52We1cCsGYaPpW9HCJLXHXg256p/p1Krs3tzlWBjqLxVciRd5NqwXUqqUM73JvYi1
G/4CrA117VuBQKG0mJYRE5jAdpmOCMi8ZjcmOPOXiZXdQZw38U0ckg8197u/s/SGRCMLzrW3AH/9
mWDITkS6nDH+Yfn8oWzDnWtXrtpFWiJaCYYxVrFiaoUA35H8T14vHr8MN/XEB1tW3IrT9azB0eIO
DcEwpmUUzvVHmcLBI5YQ2mMNyTsYT83pUj6JAETIv+UHKrCbRBA4YlyBJ2JoPIcHnpeuW/002kjy
/ZOuaQmbluixAT6BE9c7OszcRdgtz8jgHvy18utyeCr5zdOUtAjjQZewMGiwQlEc2jfgacW+/W66
Z3bNpbkxPncylPFjvVBwFPOqDJhLb4eJ0z7WDRpUpsswlY1horcX2Jw4S9AAW8ypJOdBwxBRvotZ
fbajppnVqkyvwnCazddcfQMW1a6crIebMHc6FxsgDyKVHwj13cweLVE1G0jB0586dn5j6aI33jeo
6vR2Fx635ziH9iMwNPC2bNUH8bCgMAWDxz8uHX5PCy4F7ZfKCUD4iyeSJnJJn0dybNS5ZF9dizrJ
qHDz5XzjCha5Re6DovzY+4wVuKNyVuqAd39L5ctV0dP9ow/ACGmoZVM6otOMJye+urcZz/Qa/6nU
x4b/8ciD1sukgl7/jHYc8sIO+DFr2j2ybSf6/d2/jdjrTDpYDGLfKw6N4GDJGVDYHNoDX1eh3OwX
xUrUCkpof2UIY/yD8TWQfeCDNkRXqOP5XCd6qFVaMFs0bJVdC1CDsA46Q3aGytegr44+6M1/dOGn
RuT15Rr1LS0ztH/HsTmmTwEDHSbteEUjJ+n/PbEvgHgQjF/B+TB8fQDRGFH7YSoDq3FthOBM5EAj
D0PNpJhLJDTYqIba/j63IRaNIYRu5ReGiJJAO9DhuHwHGoIN+Bs+KTeDpvNSRH3W6TJ71u288rpA
GUb4g1WZg5RDOd/doVGGefimbVKU0+3eCVoqDVR9GQTw0fCgnnx1fpnQAYH4vFkNPpebhR6GjE7Y
ehXLnRKyGlUwvYPEi+msXkRQc2RZa6fbQ3xnVaAwvS5FdQadN4Ddj5Md2bMgciBVSdothzzTkEja
xg8l5StTNfozvwQ7UZpV98HiKiWPl9t9gQ8luN95r9mGT/g6VhvVQ1K8c3A7bndvGG7swIYA+pId
I0eo0omc+V85DmzFjdY9JJCjzKNtUcSG4/zzv+SdsIxH5xFh/SPXzKBkK2lScdISuYjqnpt/J58L
zGDF+bfgqQ/U3rz+UcxXNDsvLlEtxMzijOi7LYBQ6zQQ/elcbrPSVm9SK0nNv0wRsxLFBsKptTKM
9DvdFxPXM/nkNP3nX3a52m8SA7ZnGZ3Mua7gS2itcur/ZMYBULkNX2BAiUSHloVOa7x0JHXO4iab
L81EoI4RSG0WpYzxi+3L9WOUISfm7oP0hcJgGJkFUHnX47x+AQQT7T72OJPd3pyC67fLc+Z630PX
FE51KbNZLK4uQRveaNFS6u9w8NOWLDij8LeKSdYsrBEuTAX6fEBhzZXMrGw4NcX0/h8oaRcUB2VG
MYoyn9uBTXPJ8dB10Pl8BsyYnd0x0wUg7IaAw3CzupNv70UC8U4SLsHS7HoqELVjznqds2xDR2Eu
N8Jej+iG3Sk9zpmyxuDYCQ6o59qKXLB3R7jwcQPqpuTxaQIfTnU6FpVxc7KqJQoKYPTyx7RICnST
SleACOz2VdmxyS+or3lNBQJ4MIL2a9FFv9oPgAWBIbl8UbzPybj0VanaQNJxnqZVhTcWmHn/Xqby
PHwk5Zqw5NputJrKukC7lLFzvIIJiOEFF5AYxiEk6a7DxP3eZEhFfAuF6y9A+IR+U/eQf80spd5O
XInQfgo+QnbAhy0IXFEx206ExjFarqCWZPtqGhr8NzFRF5sARYcNXDofOtMPuXE3G4Y65K//Z3ui
oNxOU6YqFzlzA1hLpBR6Q2utzaurZJdRitQ8lApmbRa71hCxFxe1r6B+Z6WB1zG4q0a+TrhV8GFC
Uvc9x/jGrWcJ+S1gruJFY9G3lPh1ZtqFJ/uJGVdT+WO7kr4vAVta87O/+/IB7mFG5qJUwat9ydr5
jh/NlCijnaR2LmtmocDrTdiG8FlAoneIB6UuWd03GOnDyr3m1b/MG0DU5C2liBTN7j9Csh+pY3N9
AIle3Vxx8Brzi0cW/jwxPcFOIKHd9rZe+hR88W34LjMTXj2wo5SPI8OZoxQ2/tXJAYBZiw6e1/Dt
CEUwKVYynirU8ZkI5Bqq4UPfdLulMjeXYEyLy2Y8hv5ewT0L2BrYOT0YzFdAheXkbO1YRQW7541C
/trQ6JgE1upRv8iJHeO3kwWq98Wl8HXOg2Zp9Jc8a3Xsc2KiJR0OfsdYY/RB0B2UHGwE20NcMAeu
kux4JoZzv/UNG0dYH/aC+B6ecVL5LeFHJQVh++hVTdid9Zrf1J/7tzaeIquV4hCa9Ht8Brb4y1QC
0lrrfUFyyduw7G/T7cx6FwcJVuzN1jJP4HuznNqcBFnaaP6rqAFZD+zCJ4znK9nWWfR7el+/2Gxi
nkQMR0jy5VBp1OvHwVDyqrW8iT3M4hjxjSol8KhVQxuUGdFwemie2hXP+eanHDWkpjtGasFnLkEN
FnpDFC5UesyTvVj21hqNBIYDQCxnjT0r/HkXBopKwUtg0aT/MREQEzChk+Yu42Db3R1aBZ7vX0Nu
e4amlDW3wu9sKFSmxxdLgtQwBwU5ny3dRJdGS7ggfau/1SNbAV8AcrgRMmS5EjFN+FCqQuHv08kP
cwxPDlno5KW/y6vjE2UZVi5At9VT7//Oz4G5+zZKl415+HYG2iStQcudQc7CDg7ZeXZh7ygWWn4W
UJLTMcoXXHlEPwafNz0jzqc17qYTcFTUo3ruMR3Pt20WPK6N0JUt5TRQjYOoPIX6nHeBDAXbMZBk
lR2kpFNX1KTbYUtqBBeCXnD0Q/AQ4O/21ZbuiICmyoR6bzDmRvFw8adE62Khg6+myBQ8tCVC8X/A
4HSy9PWcoRY1L1su3w0fcTQgXz6TFXYiBdJsy95iWwnOI6K3Iar3euyPBeVCjpeLW/34j3K9dsUG
ZLTXH9zJiPbleGJErkVTcB4u9jV30k8DUewq5yhbjq0OOTGVLTPo9O2DEq9T/DhVdfnAB8FtVU65
ZQBvfmaabPQMmNWExycnTQr4/BKzjgbCutZywtW+9AHqdzXasxdB3mQFksMikV1x1WX5WJkwt6et
9swdIOz89eQEA4CrpjzSM/DZrNaQVheZpXxMfEh32WpaPLZZI+ddWIs/nS94OopH2kYP07aSOyC9
x6F5G7RQwCf7pSry9Xx4APkclQU6tsgJXTfgSr0UnefhV91OIG+EISVAGX4ye50aiMztiGs+8a9V
sGitk8sCBrGCYpt2P7hysPcVTDyYl4VRWLWZTo6/+nEL8D42BiiPqq2DH0mi8uTAAH+zMGVwABxH
mmfnKOdESiFHFihLoHlTpi1buPtWgmLH0UrYLBHgeEy4Io4omlqrzU9/T+IFwc/7vmAtjdXYwTRR
clbWTOk0W8GObQrbR+PT+XbUJBjQfdyncwDB6ZqCUQtwhXw50Q12Q2O1klilgINFaCaK5jmgFK7s
XnASV5T1u+Be28CJ+E2+XERWHvwVV0vDPiacsA5ko3mAiYMCXGTgW5eiHRWIyZdrkNbiAF12FZSK
jmf4iG1AjeaQcnmq7iO5P/nrHYwuftU1yTiCp+pDm65wbXntCWtwCxGBAetYcPQh84a4B1VmtTs1
vnxNwK6KqzM3NXW/GzfwxoKDwRBGwK+1c5WXeph0wb8QYmH/JG/VxjXq6LdKt16hq0t0aZPJdGsi
fTLesHE5W/hfgdSxWHkYU2w8S/49JZOhYuNwjYL55P05msWDRdSOiZZMrdeoAjmi05dYUzxEMImK
W/WucJqbWrLwXfkf7wC89+050B8dgU4SpBrrI3ziF1nvhV5KlH8UzbIT9GvqtrfpfODggPwTiERB
1cXchwNmH5TaiL+q6/kgBOqL4E1Spv5ltP9DtvtXV9VZIoUxMDulVCOvd0RKUI4nRbreTaXy4v22
iIA6AaNQNKqvgIXNlEeytGTTUK8nRHbd+q2TZ2N7mKONTOJda1JNRBPc35Xq7a0aZBOMBAVQB/P3
0p3oknCv+wIp65OkB9cUBvDLA0KnjV/D8Ux+gskM4tAilV8vW7U6UPt5a4XCHPrTPmHoWMhsJuvL
dnZSr6jfs8lmLL4AEVYgbs7cxT4057Fcl8iqAjKYupnUIhhDi6894ootIzD5HN9uZ7b3uCTLqvpl
yC9eHuBB2O5/LtDkryKi0fMdJnHQizYhtjytE9xvJys9ZDgx75ZKTTwWsxBCwTsRn2nEvctnTsIO
meHRghgv0FVQMK0XRWGXe2Y3jveK0+pLAaIX8AoULF2tvlBgAm18ulTXgJMly8wv9PVw/z5l50Lr
oq1LCh3g8DAcmZO9zcv8i1PefEUW4wpL7UM9ihTXMZ9Gd/n8Q0WvIJ3UT5mTosCD3dkmdls03YL1
CT3xztVSaxf2bKyXX7i7BFESNYHRZPvtS4s6Vr0MdBrli7sQ3b5ugjiMgZXLLfiwLYUdFx8EoPmd
WzsAdqXgItVTCACUROrdIoKGjMFjA9gvX0Ybi8/v7Kt8gTLY48XReLFkMbnUQJdpQs6iyXnP2G1v
gnsAqT19f+La9XNe0Hp81ZbHB1aL1Azbujxa6fAaZ44PSQmPwxnFrJJZLrbdIRNNlm2eqwN1f0J7
+YnnjhPm5pfUES7qbEMhYenVLRmOHfHwxkCpcvOKpxwJNkv4GQ54Dp+8THEs3lBauG2k1wiG8iqx
CyaBapY9MzD6CLN7izlW91jfmbdiNJSm6rtREffAtgOzCfszq/VBDmu04/MLG3eE8bqb679XSyxX
NPTPU7ty1VzEbC6yKvvVgmPkiqm6DC8fFjlU004KCAycPua2+ne7vkXbySA0GSwAVjJdUY/gmmmo
mBa1GRIxORd2OkYSQt+aFhtxLXFkeaG68rUwvR7C7HFMhSY4bSPadmtdl5KO9kZDkj/dqhlX5D70
JIAbhok60xjXmUyYZmiooZCMEgGMQO3a4T9Yc3PWV9DNHHNhb4Awe9ePfmUTKTzhwfGmGBm3r6VP
YOHO5GQIzon1MjIP3cnXlSBZZd1VYrthal3PYRPRZX6EIpK8PpuhJLh6YGOBgeNGOd9qkrnVvNGD
h4B3YEyrMbtPW4O0Axegr1dejBG6DVhkGvEkhszQoW2qPRj4dJrcttnQwVGeNey9Brie0IoOphbQ
Z2Htpzqs1FUIpYMqHOD3KFoYWzEkUQArBKC6ttNMYTVnN+okIVgV4Vi3PSnyrXwAQfOa5GnUdEcA
ichLl4R4iTXOT95MY9Q+jPh2TOl9fHeWUvm0tnRmoV6WDg1GENfwsC4DP2mUc1rDKvqMuIt5NvYr
MqPiDCJ40JRNRcKyfmd+O9oZoppFPA++vFl0o+QUISUZFrIOt1eK5daX8vAKn+Tcno5VWxF3pVuA
1d5jjUzRFZQftCc8E94vEB0Hmd/g9XAH3KTk5ML8BAKJdkqapC4q0hHoEIhzV3TKZZNVG0bIdrL8
QveWj0SAqAZf5WuDJ1NGfx06eZAxDwIyzed9PMYq4q5eKxBPQGDfdi3tynA4sQ1+6u5Ie0qe+QVR
jjPzrI/qPaQcxxrTo6bUlRQHY26EPFNjF4f2/oHKQlwNkWi7BFx2lNFT84UBsqZ/1CCWWGTIy/xN
QiMCTFyEEruW71sTcZwU0VNwSA1hMAARSEewanSRQi5cNkXT6Zq0XxF/6nFJ2EbkpvVI61GwwUxL
VqYh1iFRpTnbVLxIZM4ukBdqLB9rVTvEjk/B4qLInLJYd8/eV+7PYVCUoCXxrtLQLOnVITZAAsfj
EuKB1P0+zttH7/m/W3pHk52piRmK4hmBv7UiDBliWwSKppqKbs94p3Mq8xMXAkQlphotb+M+v2MZ
/Q8YRHmuIhAmihWdIa+/DZ397JwoPxgZX9U19s07iOJCIl6Co+by8n+grkbfsrjW0Za0Lwb1Zj6y
Zd0I1Z6fNP1/BPzmuIk4Q9GGDs6+gpNTyiXWaJwH0/JcsTTGDLOQhFS7fDYmlRJxN+i4QX5xXkc5
5Q4P2o2yXEj7rvENElYc4+PyRHiFG8TTkxCLAvJehTLwm9YnOm4ClxF4RPhB4ogXGaClIVNN1//S
Oev2CkAItwIsQxZ36aG9EEGc3d20T43dAlmfClMJWWE905ZpFGHWjc/BSIdWjv/SNCEfhDkwa6ZC
WuOEGKb27U0lDkt5awLPdJ6E8/sdRG+xOJAebtM/xv66RB4Z1GRgI4akFUnStDuGpmsN6/yLCY9w
FZBrKypxmTfkZgYOG352iahwZowR4Vo6A3M4nPxQQymGEc7R1heVDRSTgtcgpcN+W4iAsrJSmSvh
LjP6ZenqP7LlkASp4qXXNp7okHQFiO2+cMHJcc7SL0JSeyhwhzcD+d8qODA5qa3zTVU4Cs0M4jVk
zzb9QAI9cOQX2f/ynGLF29CS5Qr2LIweA4P0zBpMvNUkzRtNz5kqBOieH80iV9h5Uppih/9Jnhu8
QKw0pLYm9srXQOMPPJx/rLNM5z+HL9Obw/I42Ggg4W48Wl3eKao5doAKUzJIOx7/pGbEV5Mzk054
a6qo/nHEehrNMz59nwV3h+taOSj9237JhRqFcSXs+Ycm7hofVnG3u28MfBk7F5wTAiOwwMh2lR3n
9uTcHNySEA/lA9f6K0qoAQcXBFc9W939JdKY8dX5ZGK+dtkOWuvZFat5BYP41gbyKKzUqhr5RclI
pcE+jRB9sdRcc6aBM3JEosDn2W8XZ68lQYY9FPI7Ff0QHz5W6cLbxNnkEtX2mjp82cJA751xTYtc
GKVYbWXVPYBcq0Pw1UsBSnDbvWleNz1rSEANPz+nt0GwyYTXSbkYJIKyttctrcAHhC3CY3eZDWqX
oIgKOIN0GWCdJa46QpU9tx6kxBFOgfui8VBD02vhX3NyNBnuBywucglAB4qEzI2J8PqF2Z7BCv+1
qP1aJKk8KTgh52oxn1FUb25J9iV5+/5g+vE0n4c1uyxCCKagSNKz0Z+5b7Qk6uHnFFYi4tribhiM
P9cFML3NPHlTAHovXpiBhqRDJiSv+ukZSjlyCWAO99lNRHFBVzs6+7S8hBIlKwLCNrP94yQenAjr
vwqOeNMZZtcZsBIp+aPY9FZLw9oDyqHNPilQyR8ZCDsg9VppDuyXMT0wqIpESD12tPPKqhiwxtw6
nN4bS12UQp6bVlG7w16BgdOsUFQlLJQpWGlZXdo7p+/VzhupEtVgjo7V6VHiT4X5liuKW3ESk576
NtO0do85hcF+r0KATAFjizIwq1tearjHj9gqSKiaHh8DLKbhQJKYWrKKT+byehRje9ch+vJBpoaS
7CZqwY613e81zYWIefMUzLz5wVjN0WVbYhnqfSJ66MAqtQEyy4mAtJWBBH7PhhEiOZU/PxAu/2sw
SCq9rMma5apkfgzANE8+fd5g1f5j+FWhWNh/hwwwxquemFkuGxWfJy7aFrZ49y/EdSQ6bG1VZc8q
GsisiyMyi4jItqa8tccJS/YBDWopTIhvAAG/NdbntCrXA5/jSxQtrrzjwQB78lljBNE8l0BvQaQP
QlpL9ZQN6ZKakoE5wb2Y6ngsTEYuoA9lCPE8wg++t4DLVoNueKikfWzZ7jOWAuLhTYfAGprdalou
j0cYmjj3tbZpFPAoNCcnUMFc0v72G3p7Ko1dP1QK8VfaqU4VXWSzim27uJv4EV3bZPlcP45cKx87
2fpaa99O9mgSibd7yuWbZupkB4B+5OHdxhSQAga4AyttECCDw96dpp165VtWQ+JhhdSQvA3OVCxX
drilEIkiTWNx+6NFfNr2Y7BD+73kO0qIN4WwSTDMs5f6appy5josc+K74letvtCO9XITSYta0fy9
UMoRqRebk6EcAlyoLu0ioKpDL3uzggp7Z/n01C+KF/Wu+NbVzEGwOO3agx53usaxdTRxX7bqYwoU
CFmuodJKZuRxqOz5yy/mXBVRrJyZs/ogIxss9zfQ02Bol5Wz5Tis7xJKciOlHd1/L3nE1YIVzjta
oRojdykQjJO3uYxfM6XD8UYowNZ8NuWml55AdMXPKRdHDdzdATLH2T4QqGzp4xvusFVtNKgIQ5gX
CzHOpGZj9tbPZ7Ih6y/J4XEKbLZ9oXhab1Y+jA3oRpJUeOAhl9Xbf24qeJpbDBHpYLNc7g3mjP+G
WGuqtmrLginxWnC1v41sqgYPmR/Z4rE5FTmpzZGSIrufxrc6bHB7LbrTAx3TbdOtdAzdkLfdcYdI
WTCjydlsllPwB9eBvUWIPNdn2n61WAqdrkIIbF8t/9+0v/jvzVLvkbTl+nUC453MHebELZrqePOS
A3cW5ZIMbarRqoAwAUXs+hk/MsBAC8oiRp5DrmfCilJjeQaqgzoRZRmYuQmJXiAGhKANOJV3cVUX
aK9xNaKD6ATeUva1GLhLqoFkNNb343LgNEj08KYMgikObCGlePZkTH8u7PRFEDD38izfzBZ+qHjW
2OkhOnzlQRgjYG73j/thOcee4HSq5CCfyJmOu7GqOs7VXPxJ/3Ecig+ia2qfWnr449BDODAz3kVQ
U4ohB4SLUqmkDArp7PVTtDPzWxwDbWitQS91GE0H+JvyJgpwcJi00WKDReHqjiR7rZlBt4FPUoKe
psOrVZkegkqEevyZos/1sP/V6o4jK53E5wrP70s7cWZxsgDzxQnRdsdQBD8/QB/kN7AE+7HUUsLl
hDSrLBufWkSOeP29l64ciJQE74ms7OG4WyFqFn9niubPN15yQynbNpGIDMLvI97ae/1g2MMHs+Wi
/dK6TxxAef/ip0C8+IErrQYTrOy8dsTglMNgSD7qYUFmce57rqHbmtSKPcynyYuo+mGLancz84IX
XssEXmblsHQJMnVJlSCBAMp6//1pPx0XtwDkWQ34RWOXjQaLLNhDEJPQyvpmySR4Mc2Ou5+Ecnst
yP9oPJJppM2PowS7WslAht3SSFwzX8hyi+5z0E7wRFb6a/gHNyuq4+Z/GcNl3RJSP9ttPq4rIEtv
nh2hshnMtAoDpxwzVJItISHIzhfBSATmJZuKr+wECSvLgG/8G4Uly7nJK4wm1l8G9bYg6cZhl14r
D7VB92p5wnjWOzFPUA1vp4xurxKW+Bh7lAfJFSRc1smhfh85Tk0ktDJx9a7bLSFEYqz7wPYQdUgV
yBy2BIasTvW8Py6s2tZPNllpBg3poL8GqfdCSRBKyThFue4pBijtpzFLNFo17dV6nE/tILyzpMmB
v6+BQJynjFgjVFn7Qtbh+pdQHv6Wq8R3u283a+f1qGbI3sp33b8r7Lk0XCrT9fG7HPP5Bcf4+Est
hMjGANS7lieCvkKi62932LP0RcwTdbJA7RpFxUa50cpzc86UdX1DCuSIIg4nfObSyhLw8XkQXB5P
6OTg6s6KHKeJ0XODL7MEVbbN03HwblXBu/JF1ChnRxY0eje4YhlPlPZcog3g+wwumInSRoARTDO0
zZKYM2dvsAN1Sti+5aWygpmtup8w7ju6CHuBSb6gqKuYSrS38XUGQzvAjGVEkW2JZIf1QrBSpCHz
BcOMvm3gZ9oQpVZyQk0ojPWT6MXxdjl2zOiIceDAmY9FlaOCMSnn7v72BbvVQ9uuIDL69/14Ys/H
GJ3swU6sNG9yxZyHxSATrP179eWQJqVWojxsLPTqBx+Xmu1xHy0Z4YLKrRNh0cdoVJP4RPnlxClA
q6GDa4rqDyahywCK8OrGI82blSa+/ot2ufmvAy2ElA5fKDEHToHGrWOT2UtMuhdgHBqYc9CvjVbW
7yiQ3apXImF8RuRhO3lYVfhr0EjPaNSeFmNA1Ayb+tLTdSa3d0nYkGQUji01sqtgn151Z3UOMVZ8
xRQulykKNRgm84HmR5FAT0THoHtaxWjPLEFumM+fu8J7XpFntiVAlirKEBayYa/Vpot9BC1tfc62
S/B8PoOPI6cdMWvSc7TAeNqQPfnifcLsDFm82A9CA7cQ20aWQQ3wV0M+f+DdU5OQaxaSTkBD3SRj
tIgthPCdyzdI+paHxnz9KHCcuPlJ9BJbgSpYdFGfhIsnZrtkhEYExEWD5mD0rcvz+clmCT6PN30W
FnDhXymlMRqxpcGxip8jV6NxJ/9MEl+CMomsCUUOYlerx3fKd/x/ndNPtkLEetPw+NNcPO82t6ws
DSPlOqRw3HvevE+uZ+lt4DlxeIY6F/zMCXD/1SYoK5br5CXStSsDOqwkAwtHqaR3WCBhod0idJMZ
pWYR2L4NpqQNbXU4QDuxVfju5Lrpn7olKYXntNElOvQ1U7Td+in4u1X0wileSvdWUL0yG3E3dxhW
BVNMKBLu2AXjmAfbaoCxeIZQdrtfRbAI3vkigWOgfqZb3ArVK+uPck80r1UzoomrLk3QvyVeuNgk
7bwfaElcBem1yDF5X7RXTNsVnOoVP7lyyct6lC+o13BEPnPSDWpQLs/0B5Ntx0yKrN4va7krsmWG
Z9JHZo/OAnKFwPa73BgQUAVwHQvBxlL8H2VQv+G43N7odUSjQ3KsmWAdFOSFeS/dZeCVCMyXd39u
EAzugwT1MxIz8qqJC8NJbDzWKhC+jW9e8o4Ak+js21/QbHX9/DSs8X2iGboc0AovbnlcbSRJDjYe
P5OFfQjeMkqUxPOpk1pFrfYqwVca7xu5HMTDTJYBFpww7IbOxukbRO5FNRR3kOux+ot1wo0BOrBC
PWZYt9+5b/ruZQYHq3zysLwc6Emar+QKh4H1ys+++Mut9ekHHSqpoLAPAjKQjSz7mKOrF0v0OCBh
S1IVVKM0YAOQx5VotzZs3iRf82Jw6EzoJ6kCF17bI1176gT23taRWTENf6QgttApNzxUaWylic/3
iq7BIyv8IjmBpiuCGMaYnZp8XjCq7lfX3IUfY42kS83T3VP3M0pnYd26N/gIIMh07cUr5JbPH4z1
CzMDp7kqOX24dj8PuNtsQ/jpx9jpVNuCDAhD/XkstkZEfaL3yD08pfMGssrON6fSv6t2X0/O+EuW
QqnE2hQ+x7a+wizDOLOO7Ip2wRoppIXoBo/Iby9919FRSXxoa+Xl9GxPDPSqLJsZj1BDFiR3O+Q3
V2NamWOnJ68kGa+jIe4CEo73rqV/ZwinQs+LKsXYJNZQSkHirIx8lM6qe+Wp4z692cZ/f1Pw4Pos
NMrIMukV8eLflo+b/8Ye68jg+EXIUSYHXSYnkbeNjhtSoHoGCzjLib17QbC2edXpL5evz1rLbV/K
aTFm8vYrqoeSGUy8f6pCGMV63L+LCNdbn9BUA7Yh3G2qDo8ljJ0CcsVCCiE8hIQbemXU6B3A6IXf
GPSE1XQUxFJspxP0qPxv0qKNUloSNxs1hUgeA0AxeyxFA15b622YkRZCFZcKE8N7KBLIqGkThjj9
rEwkG3UJubYXU7HoUSqp/S95yCIP+9gm2Tde8hDWzAxVCSwKyGNDJO6t0wjAFTiECs5N3h9BlEzM
oGZm1aVAc624ZeyHNuWhQm9C5+EoUwqPYTnWT2UknZlJPOT+qNQu+g8MiwlQgZW+dOkVnKGEx5nU
OUS1Rknn0vi0XfXYxSY2moA+aZAGeK1F0mxoMBq/7f5ale+lY2r3Zc7LbA0tRNb9EBpf3RqB3laA
P7T8TvDCye3Br+cc3jSItEztXqMW1JmYCaDiKKJdrtzsimyQNMcZ5w8CFcklrT4Wi5aiEpxRDtjv
zezo580mFAKsxq55rHVu4WHEUE9QdShKQ8iwWNvfWfqrZI4e9qZWGfgsVTEJpBxxscQi2Q9VfgQP
vlcXfnosgzNybuuVD3Vm86hjKcz13wT8CK54JATxvnwJ4l+4Ew74WUn+rVdTPElFIYeNeJE4m6IO
peloZpKJ02cFOys065h+WlT8Y7KfM2FgAyRtNE/UoCX8rSlcXY5acmr0Z71kxDPhUZvIqkCdQSPE
meZxXfKQkteTSJnCJ+phK9P8XIftKwg0KYrpOe+PTvpBrTyV93hdrpBeTdKhRJk0UkKBhcp+PxYY
Betdd5JXKZ1KaSEW9zBofbigor3+ztbPKGs7zNCdZ+pHvDJ68wcB9YMR4Q8orudI7NOr3EpUyafo
Wb6zZ9aeZ/8knKXwSP1F+e63tPRBRA+SdlcI+a1RwSOLk7lmpSDb3bsMI/6zqkYv6MNhRRxgcuS9
Cu/b3rJVf1LuuXz+mqu7qG6idSlaNCgQYisCYjTFF77egXoApcDDsSSk5tPOzV7P86XxVojBMuld
DWEWA9yA3xfucpT0USRYKmGxfxJVgcT+wASuygbB4nhiWB/3Wby6oFrX4hMCvhGIzfwy/ra07/ou
eg98auLZm7GiOnUrhFkAGDpjmMrljiimc1WCfcZFphn1PwCEgwADz1AWOVKi6PBEhzpbb+8RucgT
vhYH7QMt19x3VOU8TA8YAEAo9cStVRh46gmJubrNxKXrMddA200nUoKrIGYT4iBRqCF1T4NCETD+
Vn+kQwzlEzwbsIYU2ctdT5gTW2MsPT5hmRQbUh3w86s0nN7maC5IHtELDs6/Q1b2eplukKYMnTh1
rXIW8R8iJNbzOUQs9PKKyib9mstBU7kAHqBwDBVI0iSi5thXZY69kG7CqDUBnEGJTV1JCpqN/MBC
HjxfstCBsoiV5wK7IXW5pefBgpOw9pDXEjAT2K5tCdnDd/TYeXXXW4OThPaCBTzLLvAFZInmk3nA
+TrvvC+eP6HmTGRcsVszpFqjTjp0FF3tyA4uKXm1Skpz5SCq6dMZpOYOqD9NAxeSZF1k7MGZA2J3
PncpBWMbGwSgtRExOmPJd/u+0rCRrxoG56/jPPqJFzDBxuWRt07pdzbNMqnpT7ohZpoFlU3qD2gu
BiVUfqtjsUTxjnu89TpfzkbMTuNyps1GpvZ08rIj585z3G3HwXVA2oii9HXgnp5jG9XVSMI0nNeG
JX/t3Mu7XXlSkYwgqkUderRkcUeKXn4yym8i9SSmH30K30ivCQXkx7uXKAM2yk+3MzgBlTc9SHLV
AwU7nfyXX53XDHfCxZoXNiI5ExYOmD03D9TwRm2OA3ziRNkgIqT3jHtGW+9rpy4+UzCIpOecT9mn
OnB9ZIulkLeB98MhjW/CyRucm/qCcqmYmClpxq+8OmZkO4mkYEsn4NUMX6WuU4iBS+sLUUcPuWq+
MyG4LOAN03Tikx1uyjVoC9Fqv7cOh5c2TxrYARJUL8S3emNLgje8odH1mJJLGVOAwiTKy5J4cYbD
FXf4VRGZQSg6aSqPEZYMR4ivnBKLIKnruI6Sf4LX4qnogDvG1OmWS1otTF0mmGHPpC/zdkoI4M1b
4N71P5f2i6Ge8XRCfwD9xXla1zIgOeVq2jGJ+7gLM5N3LhriDZH5WL35IVdP2RrkJrMKVaZqVJxW
j9IQkdthjWIs9f7Lj9PTokI8iAEoXZGhgp+yfat0eClrpUXNLros203mIjGNRSn8KwELqhdQJoXd
r+PhO0lLAfWCWj04UQZLKhgiCyCV+XbbKyinn+xwEvIkUN4szI9IOEdqj+4in+5F5LiXRa+EcKvd
RqjLbm5VtmHspz5VrltYkpV2a8KODGFRM/p7XVl+3clDJvPf10kneqiWAR4DHy8c0F8aS2Slh58x
YZ/NVrbzMQVTaCd8kgnc2RzIsVK3oT9Qv+l/knuN5vfQX6FxA0tG2UkY/VGB2d/d0lbVWc+FeiiP
k+GFI+rJj4PPFNdxwkUmfjdSCaVh52rFF2WEkuLviA8FBZo4lGUAYDnzKMbrqszylcZxSuDX8Xbe
sLYjvd2vyPs5nFdv3V15+6Vg+WyrbbtHbEbDgSQyTi7qe/3mwOCV25JLVieSwZ2WxpkS6kaMbDzj
We3G6w1fcjMZUy+ifVGEQS1SS4nHFwx5kImM8W7Mx7QpYNU7etba1mKYMEWAuAVx+VbilrGYVA4f
Gv81sflRCgAOba0TicgNqkIc/FfKJrVT6DFXro5CjH4jQRrxeGuJZjCA6YH+L6zlg7oA9qVQ1VjC
d6wOCuyON77war4LlBNDxIsLV4eXX6GozjcCRZHVRVuSKb7ZuK08KgvB5L1TCGbxOwla4EwNrhCP
L3pBSqgaQ/PMn4/RKo6aoxmFO0jyXTY8fxG2FdEH93tVsxVg47r77cVlzkHquGg182OOhViB9chm
ZH6d7De02jPj8AjETgc6+aROPLyirrjzjHYmq2QcY997AvETLi0UaDcSHUpNGqqqN8lvOqrBNP6A
GJmDeK6WV5lWvP7C/wGI6vwoM8ikoiae5ZwBC2UJ9HimTNBb8ljwgQg/vuMxC/gw8cegY5ehul+u
zuyFjhxx8DnljwLx5ewAQ9mrVxJTSDbpx1oz5VLd32MHJueoXXSxcxTVWK3QyZcy5kSNLcpOMrYL
Fq4GJcaXAE7rXPzg97QS+ehvQpR8zn05p3IzpC4GOQGiDVK9vRlGlX4E76ZCQFFT4qPGI3AJEk2V
8d9LaeF4yCfQWgrRbymbA28NsIDsX3p1RYIjykeiBMZQkVd2Wl1G+fxG/b0n4AukwSutco0edzUm
WXgTT6awB1AoOiCWkjIRZYJEyJIBJDNjimQkI6zgEUeh7WvmQ2JGmrpiovV14GAOqfvuWaR7cJYq
FNAFPTCYt5z1K16WQyqMW5jpEDFksZ0flGVSB3WiB7s1ZKbO+5mhXsLZ2AqemzPiioQRvRA15WfL
F+zI/wtoQc26/CKkj0DdlOx5Oluf1nHbG9JJOykpATIb75fk+pe6YdfEcCDPcY0Hh3EiAA7SBcdH
yrPsrYlEmnGI4+9kslaOO92gGa8AJfgyP+VCCPzv28eydKyNAWissL1mL0coqiwVPOepifQsfaXY
JYuVJaTMOoUS9epIQfpgvA+OznlMNQZ+zVsakOfEsr/oAJeVP79xJwosnBqaqAyEyXogC9J2Rsqo
xzuJmMKkKaHxSL5N0zkJuM0EkpZRwAakLvYLkt/ofMNEdRhkxSW2LG9x/9tPJMJfUFoPNxKa5q+4
ZEaVcvIECUo67NLJ8yLSuNVIMek+D8rL8tN86jVt8GpzOSsaRyBBhTNAA6G1VfUKPLuzWgCPyGjO
Nmj13n+pVwvRDgXc1paCCN4NNALcqjLLiF/X/r+HwYa2rVsoGoLjVHODvpeO2yC8Yufc1CIIci97
vYwAl9cw3sR31c9OvIqcOnH8zhfSV9ZO07jRymfivr/XS+hoXZS3UEdfZFYaFCrA5uA/HJl/Cor6
/LcRBVDA9DwS+3XLAHw0vgvENumTmodWpgM+7vRY0rN5CI2+dvcF35k+HJfixh024gsP1I5SxT3L
xrtyubDKNjcRyx0CzmS8k0vsQrkmaJAvMBNCUnkvMHqRnvv1jvXEygFQHZ8x0bUvMkUR4Pg6GU+Q
dyvx1kIeFWCm/jTYMZqawxtVkEI4ArvjBrnuEx89Lbp5/C+uD+Sjgf+lBs5PkguEbGmGPfFmGWCJ
2B18bU0aRbnx4rVLq5nmqcFW+EeeNWkarEmE3PFc8H9rqXTwu/oNAb4lNYnQGX6SWxt0lP3OBhp4
FyB1DKVJgZY5GA3y37ujYjgGqg61/PIXg/TooWvjV6NEV1GLKTMoBqwOSKIDuWtl7cRfsOV+HW7W
jbEddqXJDSLIKFbJv3GISE0n7gGGK16ZVND0IJ2vBz4lIEXs5e11j40JdXETGgESMxp/zpeAg9xg
LmV3kfePzgWte5Jk/OKKaoK2aZ0ccxkMh0nRzwrfEjNxXQahA+HYiJfMJrmF5ZFHXEcyNuUxu5om
VlrKZoCVYEqcUEO8s4YtRPq031oFHIuCeJJqE/380sMcmkuVDV6L/J3VzhjgTTgSIYWEy+Eoy32y
8JWgiGy+i5UzmCGUU62WNKYxyjwqUt3vtsObjZVz+ulG7w10YUiJuZwmYwPYjz6z258z2a11ZlLe
rmLEmV/+B5MAn5QDzSVHrrX5ohKOsRykr71FrZiq1nM0yIRv8ybfkpA499mw/VwPg1ZWYCYIfNoP
MWpQ7hQdUilPuzfhAUkIPozdiA2py3apGpd7Ljo6hL43lSPZTbC//MBVfBj0pzXakWELa8H1KOeq
sBukyAWGDHVMY5+nTmLHUwRZr03LYKEroipmemhjoQA001TS/T6wMW9+arBjvHamMX968jUV3/9b
w2pGZVl3lX+rQgiFtkHvn+8jb8SayygwtnWDbcb3aM+/1mgWz8RhBNZzRsd4wMGU+09pyM5/TqjA
gRCyZfawvqiwNaxSslwvWNMtSzzLC/lCs5S5InfPZK4D7nb3TwZw9ZCtoTtAVJXpyqWAFR9S2tL9
tMeF3hTqcr5ir5/jG8llj0OyVgXtVwYcFn5EbUiQbyiuxhK0QIvCNdrsNdL2nYXD1RmkVr/FIjy0
4/AZzOhLHCqbM6VKFeZ8Tolco7SastON4uMKgWoUiehKSS66dJF9TUH79bcpLJLZWuQs7kFxOkf3
iOlnyGQD4J3A21smI1e1N5h3QEA2GVnonXG+XyRlU2oFiNlvGAnKRHYDB+9/aB8L5ODhjfqT4097
2hTHQYemfceuooqxzoOEIGXbd8POMZ5ujoTLazBYsbJoC36fDGh1H1lUFxqqDEmrq4lGjade8pYI
wXTodjFA5sNC0wkazfrCCljPnmReNVS9fNBqTXQwhxqUVC23BBzuggx7i2Tcyt3ZwIuRjFagarIj
yxPeVB3Qc532KtxwaBRd2Vz58GcOpVh6lXdC4m8NzQwzW2KmatVOOLBP8kFXaBosU4req4oLFMpF
fvq7EABi2Oj4Iu94Ce//yXPDfFODb0weIHR8ODpID2ktBPCx7pB0F0TKKPNJmWmDCV5kpRusEdvt
S3zV2ueDJ1TIo9ZlYikH9/5ranrxFWk6pxm6KmeBXlMRCeRhD9+DVYeidU3HYHfgJfnWv6Tg8Ew2
BKkKF3M+vk/nqDn1eMP/HitRk2Ii3wwwcyfFaNre3TDxhM+iUtjNp4P5OZq7VYfA7TxzXWRR+Hhu
QaI9KjqlvylnOA6MLp1v4vlXTHi3sVn0TC5ihyACJlV+xrFvZzaqGMqXhAgoWzlB+4FPQtCJnRzV
3b/HPR3/H3mRZ5vc/MMKyo8wA5POlkXqnp0ac/mEN6CmZP+Roi9ekr4+FaXbIvE3PwfQ358kjDkz
JKZtVmYGaTkJg4dyTErS+psqyTcIRHjFjyTYdtnSYPx0Xw0oIaql71P9uX39zbjp3OrMurWBnuxP
hFKnp54lfvfuJWFKg8EXBH+wlmqd2RDK5nHIpRZlKlgh/JxgDs9hJW30K/l9Ux1jlrkU7WXJ3Kl/
iR0/w8k+nzIlTIedQCuC7a58qxmvf7HbbFBc0gKsSdtp1IjYkSdxTxezGIPJuTDI6ZCbd88fh+Vl
6/bJK9IJv2svlzj6q5isIGAFAPpGVp/bIIDR+7ihePfdYILdbAK2+xsDZOT8PyzNYvbhhXZm6vqH
4lfX1JDdJGAXUN+vKZWo4ybcJkZ+UCZu6pVfGeWZKHb2hNbqkH0nHEaSJw2jYxg7WrinDaA8VbR2
UxYVLTgofrB8mptxQVhdIx45AdhNhdA0a/gp2ZeeFTO4HVujC8WHSg+2/nXxqzdy1ImU7p5eP2sY
CMF7SV9L3zDFue9+8UHns3acMUCWNw40M8Ws4DeOfn02clxRyio5vXsan6aoGixNXe2hpuqq1Gpb
AAe7/BiVXaA7JtWxLEzhfcxjsdHuy2V82aSGbeUydyGreUkdomI9amxeBS2ma3HMXoh+8BSsNLYZ
kNCaalM8wYyD1nPeRK6OpiI8yYPbaGc5UNfaXDcxv+9BiCYAWZm2P1llZA7sriVKGTJEDRZupLQj
9vmEBkYr9OW60l+mtbNpIVQP8g5oSQ7rZ7+tcG5GPKo4EnuDebnZAJHMl+bdZJxrAMSwxEGAvx7a
dy2d/AusAoloSRVt7QofMZV3bsg4Ho9Ig1UpiZBiLSseDzl3LEW+XjNwAfJYzyBfMLi/vM6mLsS0
SJi9R6aIbvG8BxM6qHs/KiBYhyuGI5eMFAlgzenBYMya7IgMXGVfJG91wqSIMX/se90PaCFvYkQt
m9eMmwbS1HLUGaly+uab5vDnf1ha/zLdMviVWseN/d6/F7qvA9Ngs4rvnbs6NUf6tTTv0ctvbvAp
+nPS3KQVnsR/o+VE82KgPaREO8iZc0io7zKW1+puQWDYRloTDBjAA/Q1j93N+aHCqhaTWOYN1OsR
E7hEXo/nYdcgtRohtvLIelg261R3816rD4dYhcbbK77sSpYClwbeeCMa9j267dRlF2wIZ+5yve9w
BeQlSt7yG/ev4SJ6tQfIn1Z5jgPZUQ7N/EOz1swXCWy3BmGkjaQnLOmWqHGva/eENIkiCqZKRrze
F3ny7lJ8tmVxAp0WDThHMsm4kp19z/KnrfuCUlpv4ArHEva2XNookL8UL/Hosw+A76U5zIhfSrYq
KzO8VH74cGXzmkYGF5LRz5E41z6QEJHwLhKIPPuQ1z/wvnCt4/CW7vKxV7syei/l/5ZmnyiSMpTM
/A9F3uzC/CuwgedXKJvfK8O9KxUV28HMZ+XkiiGyZo5/ThS17PPvUHR1em/h6qiw55MzJqISViRz
dnZHh/9koVFaYcQS2E2dKJsWjOjZmIf3X0BV2lJ2FMoj4sQD/ev7nTliO6tspi5eJlvpGbgvRQAl
80rb8S5xpG6CVMRwyX+ueMRU8GI+/hLV6Tuzll5LJayYn+A6shla0fQdLNUWEGKFo0CU5oBKjc4L
nQcKvmpdp9sZW4TCvYwKadykSrx73E49ivWwXTjMd6IbiM3T9WVcAzCEPZgv+mxdhkR5JIoKhs0p
4nt2/hiqOTW1eeLZVui0l9S9SmKhVNWYrLhooY42OXeKvJ76/pJDoPuQ8HAitNluKxjIzXTAeQ9r
rbhX1wmV8JxH1mUkwsVNh4CG3EbXti+EaGkl8e6dWmrD5RRo1i7BgPNbkiZjMjxzufWBNxodTsFH
x3mQ5LkqJ3/wpNLNE68j6tXu1RTklZqJErPMXAghelu5+aU6HFFGBTGrialOMh4S4NZe67Wijm3s
kVTvEqUGBziMKRrw6AYr2iAdkmlUBRhETjggk6J/2WWiMtepnXlpTP3N+biVKwMSlYsZcIcPpTVQ
78TvpujarfPOpn9C6nV38GI0svFBky7nTzgsoG4hwIAY+7DYerFZ6dxc74i3w7xV8iAJO9JgtCbG
SonxikK9bVi2y0g/QLhtaHMGAzNBNEPYK1pis9x+FNkmQBNGxizTYQDKzsYJRODW6S9bAiG9m8at
dUQCz/h7IsYCxhBm1eTeetBfGD9UkZbmMrPP2oQ99kNNPwSq3L0Btz5lQFpu7iNvwiQZ3qhShryD
6sG0tNTya+7oZ1XiBY9Y8Wah0m1BPyQtrTOAss2FWtS6I8yBcmz4b3JNj4Ixms4CjdEN3sKEfxnq
QBKy7oO2zz0r9JFc9SflB7/gNFGWww48jvn+ZSkgcl7hOOcUyxBGoqE94lDdV/sMjGcCMrq5ga3O
Fc0va7uFcBscvcpoJNMpclyGtd+0LbCNl0FOHt0m8q0eJ8/t2xRaZsw5G/Kbg6j2PfuLg1so3DhG
983rNI9V2LcF4L42V+uHvd5y+ToCnJJEDlR8+uRR+TVEq2gaA1B6JmbQd+rWPCxLzK7MpYmG9jB0
bviyI5fyfdgIX6NsZTjVQ77mCBXziFf4XmvmzzgSGCWvl3+0iyU5bD2QJaKlQE1UcU2eS5q45Xy8
yQiwT5IWT7eU5zpm8TtUKCi46FD2ugnu7dvk0QPrI6VngnhjKGHqQAJMjgNVol1U/2usOthKbOeW
lqU3URfnE1go15Fy48VN/VVVcrEhTXC+sOn4czGErhf00LCwnz9ZbUPe7pQX03b4P1J7CBquROdZ
eheIuhTOEvTQP/o5V5KLMK0EVR1zzR2tXjzexoHMabh+bDACNAJFn+DSECpBENRhbDXXWNV/Cnt4
dyinMu2CQdYCHsDEqc53LsRIfvC5g2hJM8rQjADjwFx9a2CR1eoCUg+ZADV6uhyxdTAYEdieCz72
g4iNc+T7ttSxkAIzuLSw8Z0LdXKXtKIK8bDhaV7RgDKlq0WOEcW/mzKjyUXRlBcoi816kaEyzgmW
8o+p7mIDIh/t4VEIuY0BEJBjDaSVbpak8DgK2KnI3aGLOuDzyO1sPRwv4K5RfXBLd+M6zJZ9faLn
iBL0YYG4a2i53uxgvyggMSkpok+Oh+BEw18NUwav4beme1GqafhRTJjXaNQIurTFM6p43vnNkq/1
KUh4SQrbm1tUX4CXABJcyAuG0JSAzCyEvFyVOCt/U1bIwyOemq0BJf/SV429ClPg6Ov0LHQqGyEf
ErNbtsHWJBoVlzToBwJXveRqA12fXU6eGrxOLLrOaPYmjxeQvbEvYgDa4mEgTEFbB2g1yk1n45eG
w3sxzLIABQ81ZSgGVkyRS7RSz3TUNYvHsA3oJgJ+2Lr8T1i1goaOhvvPnWDf0M2W7LeiGgAKWy8u
6pjEcuwQ7eHiWZmGbph06cyJ/3p06aTPhlUABkUSh983UVHs4jiEyHqjZnHOSbOlTQIUHfpJvjBC
fto1blXjvqxqCUNcF/2q3AFIJrnTY1WGwnc3KJYf3gCBpfCJS4K2Xx8k3n7aSoddShGCx81sq/TN
eJX4IQjg6Jk0sPor3J064IsQci3C4iBV9zq/nuhlCFaoslQFINrH+nd8ityWInYVKXMCz7EgpcYm
wxNVmYkw+HG/Afx143bk7ypMkOd8WNbh23DWQiBX5B+1BzdmPmA3fgn8AKU/ZPK9ATKt8jgVVt93
cF/DwfcKG4yzEvzdRHGDOalFzaOlBqy9XCRHswlpZsM6wEDImgy2PyQQglabiaiFZmRb3soyztTv
2cE8yAfpgzuVnyhWu8D/BBcc6kqDaaPxWd1klhYYmey1jJwn/pKY3sfRQdSYNlOpfVo0VvxGl42c
Vlzd89o4ZeGs1Uhl6K0RMTw/0LArrwislCdY1A50BWWSvgZ8Q08IfJT80RvJyOOGoef9a9qBxGSZ
FNL0OQKT0+WqulbN83/QggLveucMxlV/IErJWgI5hyFbLyCo77sq2u+6lSQOIdjqCy8qktBSMGci
0IvjG6qnNUIdhUKL+2OtxRGdjBdPXz6Q2ITId3kt+vei0D2UjoNS27PjAiiv6jYBIpTKEOWMPVGG
muxaW8DXAGweYpy3o3sgyIuRW+AfYqz/XYmYd3ICAyBUTXIMcBMduBx4zfyHbJ+ODrf5AlQWJDuh
/dyWExUu/RNwdhpa1HcmRr0LV439XRORlnMar7sNfWFKVQGJevUP6L3x1VhQw7IpCNBRAzjU5jWH
7dUJoCXPmLxAVVQjcBhy9gt8Ix6KT9t+kH8eHJ2/Wd1WR/GC4H5rsktA1muGMAi8yrdGUqItbkwp
tUwcEYNtGGjsbAN7o2wyDTidx4oeMTs4arVVXKfY9Wx5gAgVUBLW6+8+SLzV8oIaluPN/6iA5Bxs
jSycwfeo+3l70RFlMo91tOzdWVs1NKvXJ5m+jE+u3auqBV31ETYt5ulnLp+cWfGBZ7b7m97PUXDx
lSNr2B9oV0PLk8j7AOwSlRo3OZAUbYgyIyfdqpHjCYrYFh5Cl4783UtlAnhnOvkHdGrHPVv19cd6
WrgalbQW3ANOQ4FhPQA87lI+6DTISYMeFxaDdLltaYz2pky0m0I6COfMfwgivnZ/iw9KgDQNVo3I
mtHlAQmPdOIGE/d+nfRun1c7saQBBY1JzrMwWcVDAS9WYd0bDq/5w9zhQRkSGS2YDV+1ws/JwB7/
xh3/OU+7btSebgqcy2HcsmaItYRSBO5lUp/gm6+wGWgJ6Lm7Egr0jk+rGOceExRkxBWfPLxiol1a
tr2eii3OvE/MI69egUzyY8lT7GwHPpsGQ/dH4IYY0EbEVdnaXnQbjH/nkCIhY+JBT2tJi4PBpzfd
g1zQMlxmg+rPoetYTio2JdU0kJDIf9v7bYE/I3mWFwcPIgWSjS2/G5qaX0umlJAbT9PXUFPD5dlz
xqd97WOiQpkOkaNb9cU89GZhcrM2ORd6pA5NZIyEtWf7fUPbfzhS0sRTtBJDV+ooEiwAFvqbibne
hCXJzM+V/+l2M7hwGSWuphuDet1kFgkUwdCqgM69xYzJcw/4gm1f5ro6Yk/ETeS55QN1F6WyReDL
zzoH4Tg42oRWzhuruXxKYz7AI4KApv56x3Yl1J7C+eV/LuuMgzbhXcEnrWLIegGKwtP4EUlvZ4TQ
ys5d47sMtGJZWj7JzZowshV5gzqnXHP7dx4eUjfZ2RzcGJBZPJGzvuWFL8ghepabn9YHNsTB7Tom
OQcXihM1/HjFR/W58nMLgiEqxN+qQRuq0nAKhUI4FyZKhYAaXzuYowsTGBRA0abFF8KxG994f/2l
q1dcbFfmvlFs6jrOXWp0Xay0CII7SYqsQ2vrG6zl8NCnLlbGm+wKl70K5JjRMCaCYb38LsZgk8y9
xO6hnUibhbkbyHud3IRlI1MmDU5YguACEFlYqUk5dj+l3o+iCEFTKGoxPcLZE9TNfTycarBXLn9R
+7quzahcMsx7UKvLSytlow3udCmU0kqfDDLILidKCT1cN1Fdpmr2WpSIuoEtdWUnPS+R/dhPTfhv
aRqMNx7Y2VDJHwrhXip8YueOd5wVNnrt5WXKj6n3qayOFaGy2v1Bxlr668cFrN/QaVZxohvxwabG
JFPd4fa7OWZFOQxISXcb8BHkZfYmSQaTgAQhA2yovoTkyvhiYi5/n9W5vu+hHY612jk7G60ZJ1wV
M1KeGCglELJir30OmLcbFjqN13e7A7AyKyM6apvyRu5Dd8Sf7m7MlfbsxWDt0BTwKUJtwvmX4dFj
dObmNuM+mFIKF1ImtPo/kCpbinJG5rdf9/LqK+eyrUQ+/aYNQCOML3aBdkP/+sk9DE+p5IvuZyq5
Sd0M82ugJA6TWVABXI/3D17EOGERxg0gJrsygzBE/TR4HxFCv2vVdsjNxduh28h5lYxDtcPsoyc2
ulJ2OQZ51tOJVzN0tPMMO7IdKX/6Udn4vRVVOnjutmOdcLBv9OBSB/pnkJaTeYvN4JF4FW+5u7YN
2BraWTjgTwwv/dAoGFIzJbA9M1jtMzOJ8tufDs9ZTY4MlSfMq0wpH9XJyjQvyNZmcWkUfgfEhw/d
u8O02TJLBe+J7UUnbnqdS3k7FbP966aX8DLh1r06QQeRF5wDHM/DMTF+4O9O8mRb/qxrHI3Rz12y
RKcH58bs7OmDGaoYgqwWuWOh89PQoYvDNfAy5v5GRUrZxYtE71SW6APzK88oMrbtgnvdoessQiQk
ETxb6uvzkSX7Mf3byV8n5GAehKb54RutMOTZ1aCnIHk9VtYqOmUk3pyRE20Aeglwz17/YTAJq+vP
OZ4U0c/rf7ryMxlp3akrWjkOtusHlNgV5VDrOK70a1ew26OSY6eH5zbD0AHZgz125Lw0M2AcYbmC
gX8r5J7RBA2+ZxGDwDw34pJ2ZvaLLUYZQ9aeeWlrPa9Q1GqgnMN648QsaFirneK2Rr8bP6nNEnPM
nCRkHT1qHO8DOmOQXSYFzgGRTs3x8+qUQy9Z5pl+UE6GNMz60z5m0TSIZQn5gCHEhCijKvdm/wt5
e1EnyYonnBFjPpCwm5u9dNJJ/O0/2MGS2VG1DqqjabzgrJ8neo97hOYQD5xTMXA/deoDkBRhDm8L
LJ6Ti0PJECd8BRr5xkbkhlcRISGjvWNNdg/dRTXgLjVdgUPAqRiUsxJmF5yHnawB7WzP/zt/TuFU
8329bJ7hITMQsTboB1AC9fLCNVpmsY+DOsr4CRtzo8nnNTUEqX5Eb4fG54M6chTp5N32DDlbaT/c
eweUihq1etqLidqAXjXj5oVI9L01oLbenURDArrUo3ABiDiZxoHzZCAKrYPED4CQHylu2ZsTaUkx
2qTWqGfWHoxbjJCROZJ50sjaQYYSaH/mUx3dhSjTOSY8HSmuqKSMsGA/wG52b5APYSC4Dd7halW+
lld9H6k2s7CtbPGzPv+Cfin97ARHyHWepmmuHybVLaWxKJv+ybk8yrbUtYBXwp44asncUFmo70ym
azPxO3VUifNCHFO/vwNvwS79BO1HJxalI3HxabDXF577EMNw0PXNyW635jt6bYnCxAn5gal4rOvg
loBEkSc2cP78nFZIXhLEF8ZA7YNZ0amBdt/AVsB7wyzY7UXLgiwDUweIVbSj4JD8j+HIVKhJTU56
QwjHEjJj0MOp1OBBgYvWKY3rmucnaJKP2c4FnEAps+kFuXAF8mVk7FisvrrAaVNwGNjeOyQcme4n
ogs0JRsEvD0xMjG4mjKqLsPUvXn/Nrkpyy1ogWVTHf4cg7TP0j/ED2VRkA4vjaPEFSIDhaRk48Al
xlDv0NdY5yrz6cyxzoWIgrgRigmzSiXkdt4n+qtLuk5JKZq8pRZxT2MHdd/hq9pFg1VgxVH3Vkfi
ylaOVRiaHa//I+2Qt6vx17TUI61Fwb1sB7F4JaMBZ5h+n+MKFqlhDM3H/q6JVUBgsZgXTpIxAad8
Ao6CqME8tssM2fBgDr3wCNAVh3KAHeRS+8I82M9YzDjMvXpQcTfJ8bRGug/TYyoy2186GKfXG3yh
h8zJ2bPXndKL97L7u2TotzgItkzYczuX0AOcyfzxizO6z9SSO/gyMJgbKgGVki0Zt0ZdDIT74Rrh
b3/U6GrYFrmlBTlnCbgvZe+6zIKbfBizjXvhBTBGWg1bxzk4RYyXlS1ISHEPDleoGcROX2tvxpDL
je2zyCb1WmJUcEwuZaWwWwZ/cwGc58nevuiZPrqzcE3R9cy1kRUA+KpQHcXdzxThibv8jI85h4Oi
GIgZp3bTqbWHiwFMlb0eJv6jTnN5kqAKxW+6gW2D4QeHOyW0PqQotuf1Oe5GLJrr9K9gL6FKmc/l
3I6c/JFY95OtwyjS53TofwxWj5H+JkF/lQIsQ10fX0iCuS1z10FBsQwGMUc9ZbswVqSLrxrPtRVP
nnwqUAb7JmdFVMWLP+KeWZtTkRu8jpTRPXpTzhuHY0uBCI3zUvjvxxFeYYVpSCm0IrXd+CiKuosK
qBaOIqRaatTV1ViYdYLpwS+O8N49DVBgsWEJlRNtqj8ly/lnx4xrxnvsKs5vqRO6t3BHdarE+DhY
nbcl0nnPHfn6EMabch3qt23T12AYncgD/TyjGyfAnSX9IYaLa48biqKA9Flio/gazXccTllCaxxI
EFvIFv7Tjy/FMxm91Nw314ZVlSgxBniKOpLCWaT+9GUcM8i26L2rE9ClwZV4fsiYJwNAgGFZtxli
3d+MPx27tWAgaWocTVjGISOhzK4m/E0aEgr1OJwG+im+YKudMOtN6wPaRQgyEdF/asjy0sifQdbi
n2KacUPIiaARO7P6cgo4zqKbBbd6yv3h8kArwyD8vqb2Kbx6S7e2nL0RTuMXScRt8pv9o87hYRQC
I9sLUKKoQGz85j6DsbfSuVYMzzNqJEbi6TRAYxq0X7wOrmex1mZIK9+TOcqWCCRwzPUkvkz20mII
Flkb8ZprUGGHGbRN1BNMG93qdNdzNpIhi/PH3QxCQ7YPcap/SoD48PlaWjXh/Eh70ccRKgDDSYS8
BIBZf+oC2GjLmtoTJ3gzDS/cfhNpCeyNp2Czn1u0cG01XgCPuPiw8rwZjcmzH1YDp/uYH8R1nz8o
WV3AZhc/OjTkg5pX+ljI7RxXwZfdtGRZiYgzZtEzmaRilvxRlqBVSjEeVCQNJZAZjkUDz41hBPDR
1cRZraMYTe8dhcgKXGPzyiQi3FaHVAQhDKnTLcafV8IA2aLG6aGNZGxJnxcFZrSStar156Y3bno5
/Xxw/GuzP16jKG2T3DudKihqHwSbNO6qKtgdja7AeF+z41BwMwowfXQTcTsGuz7bBJPwPEah+kj2
WMO30ii+ipBRCKl4ZaDayrLOMfe342Z1L74UZ89S0wdPnoOgDPJ3mrxp9hri+ZQPrrnNU38brH2w
ije0W2aEjJj8fGhRQOM3Fp1peIRCGFBzPl9Fb0jABKDw4295G5Ui7cmVvKLcXTyiKXy5YGffMbBl
AudThTtSWMjfxFcTgxcbPxPI8HIBl6KJZcxowoIRMkCATb4BAIxC2hiio7RbT45MCnIXCcvQrL/v
Ii2dUU1RSz7Kuq6yZ+9lnoIQdcc8UeNQhstGq5nT50USPzyW5LANW9HpfCeJFiZUHR73Ky/2+ljy
7nDTQqwJMnQKnQVbx+cYrdEyYjAD1VibP8tckXsiYQ+QlGVGrGvcmLZ4fC+YT/WO12Fr9ijtwdY5
siP8hc5y0iN27SthCukH68YahanflDnQhdUZbjmLB+2RcWH8Sy1+qiL/oFU+1mIlteTbZCUoZ/Wj
qpfgrLnTJEETZVPpkHTxuXJ3U5jd2WRlRbjGYjqYG7E8jSSrqIXda7HDCd/R+G3K+EoQ/L1TV7WA
hn2RHu0kNOT3wdNDNOHasfN1iaSWE2Y8jkp0t3MCLUpFfUiTGpS89dZL38An+ysmnpvx/aFgiShJ
nzKFDZMcIwnFhPUiWX802gVvrVq4RZRM64j5xyhaRkjlJDZzmPtxbFvhayge863s/4w62xR+kkfo
rwkWmGdr0JEeUJjr4+yzYPk0UovQUAdkKzEW2kRhMQyftQoAzzRceE+lUpTyVVIK7mCF9UHwN94v
ZD6b4Gsb/vtP5rLrR8zF5CLSar/WqnBxKzLhAF+dwy3TJ34aNmXyBMMZ0ZUKmyQ9fT4NZ5cE4hA0
kNCd3G4WiRkoADiDahMc5uuAJNi0q2suX1zSLcq+Gsx2ynJGjD1gr5vjwluWcp/+VWM4ZxYA4oKh
c36tvlmO1mm/Zep0xfSW9TAaMzHkklpQtl1auuxdrVBN2OEUru+dsnCwkamAxhFDCju3SsERXf6T
iAk07AGZo/P00FMHGvZAmOafrBdf4WVWgLBaXb+G6g9NfyzWboRyPeiEwDnHFSsbet4kidkeBGoA
YmussbiQ7jZFlSDd0W2t9UkWIp3v6FQVHK73KbyWk6ViQPuW8vmqqYXn+zXwh7PO8KlqoY3Y51J0
gJnv/r1khsk14eH40shI1xwvcYdmiOL1GIGiV1xvLKHxY76EfvBm10v+G5EODZznIHPSWggNX6Sx
rXMl3VVQ7/JEp8YfRxHE3dZhoFzoZ7HZjmSjkwFj8As9yuZdRUW47cXrhNxArJ9Ua2ueUTDKBi+5
yXTIOvl9dPqygLcBISeJ/H0otS4MjSdDtS44Ssyz2JxlRkRr19RhIyq9KwwuL0+CyJEHobL9J3YU
c5wQhqkpy8QDIIVGoT18PvhR33Vrb5vorYz7NnnbL43rxxQ05QmROviPpdnmuGhi52vKJssR3oLk
1Ua2BoY7YgmhS+SNB6nOiNZ62p6jM02bWlmcVx34san+834serzq8JISSQlEyqGWKudvkxI7A/98
i1w2oz4V2bV6XYdHYueLcxglEMMXdy5USSprZcl8PGqCvy8Iytfc/6DlCDTtZ+Vmi9yYd++zO4gX
lcqda6oPpK73u5PQUiF1pWqaI2lw0GOBWdnHBbcOWqfV/wRajSb+LdfN53avVpnWmXdpBvw95JHS
Rkop0FmLpr2JVFkk95bspku3ZTPvYxC1hNQqmU5QihQmSqQoYNnesDWbmSte9S+asYet8q4H8EBU
VXcgj9Hbo+jJNOsjb3GL4QOzjHYul0UCafP1Uw4cLcOVjQ3v+cfULbPW4afe2mEJNx5YFKv4f6V2
rhSz8IrxOb1Mt1RWS0lu1l+YcECLYHqC1laFe5hKe62oiwYi/xRYjxcWvxoKy1pXagZ5Pht0Mc54
c+bBZcu2p6Ycu+yWbz7GRVoMTTi8LdcVbdWHSeTyvSyRhtinC3MLtH+WSEnBR/UBaMS5y/JNyQjg
8cgNEuUoH0cFLmInGUJDc+bg+Wm3DcdpJumx9Vd2tEFdQde3VCGck9TWY0YqmcCz9HX0L7qY/U5a
EqnoOuahI1gJXzYRimazQQLuUc3yf0jxXggZ5oJ75UnOBjhihLpM/K2zQtPKZDFAKTSceYgpA3T/
bq//YAt3hSOlGMSrWsx3Uym82cC6G3f9V1Mit/4nMWo8h13eDxxmlxsDy0O+zI9U3YHZv829uH/2
GMVozKsLm6PHB5roEdfozxvtAOnsTWyHWSXcPMaBk0JEAPAItY7DrCpSWubQz4AkDPZcCpG78MaA
feBluARkyudhZ9iKP8kDOcA8QS2h2Q7DJwQAGDZ+AgYE3R82+GglYz69dHRQjyJmGtbw968WOoqB
eR2O+8CudTRdlQ/V3SZOAYNi0LuNBdWBnsx/Ae+rQJ/i68PWrAxLMGk0n/CtLwgdA8tiqXxCD6R0
/STc0wSn+W6ESNDvsCLqiAEOOXfNGSzzsykV8KzbUMKGOHew043Y/m8peE9XqM/V0jZsKGjIiZLF
MH7k5oBKq8jxNQahnmXMtTS/nQH1qmKtkwxueHsUQKsluzXV7XRufoRXOihtdsBvaJxrP9N6xxbU
f3JDVNCX8l1WCWeGCgK2tcY1YXVmgYiR2S+QCjx7e+JXp3r9idD3lT0wPamRp1HSdqnl7BSXoYog
fXMnrtCiYWyY7XRh26R86LeTjLUXmeiTY25LBtTS3iagNohCd9JYKm48DI5/VJokpckwG44f4IPx
75gC1GKVMEoOA24xdWe9BwGna4zHv9thOOQmzcNEpMxlB7FUNybzCAw30GhQFGOeSKtL1ORzO5oI
zazFWEQu2lUTQDc0cVkJePgHPrNKXkZbsQBjx5AvdAXqCRcBy0dhURO7ahC14nK7K/AZ9+XgUh99
mx652u+wJLMPT2wMM9xifMQOOuIiSmjCt4Z/Z64Ja4v2oU33ZXazhHhd5OaZEPDGIxqj5jgW1jdN
6y90jmzQoxSPqt21f49Z7ziQAJoMj2tdb9fKBtFnk4PKA3FLfT0p2NiT7piAOkm816YLPbIsNUn6
kTkMmxPpnI+j8PplaXqs4iQwBUYBw7mOnCQ+VOity8koCXx1gXD/DtI6MsC5A4FziwyP+hxBRFBx
NL8CnW4FynRVIzBwlwkZ3bgUbwa35MzGlmDvdD4PZXymn3IQO4XX7C2JX+PCRoFvW3sxwJ/27wPo
J21E3jrDi9vDdhY+Q8ZBiDLYki2mxvpDQ+iTChkBkyFD0JpYxNjrxjg6QDk1aalHRiu0Ye4TKRHd
AxJyYuxZ+BaZTtCx2otbxTgFmCDTCHX9Sun0eCIpSm2/GZUvZA1qwH7u2Z861wdN4T10OgnyD5Nd
+0HZT1spjAcQEzaHov8CuROL+DSCbxIZyB5z5Zvo/SmF2i03kE+YRcdHFQmDfCeVBTxiAD7PlRck
SUnB++LHb8Jor2HslmmdxP72sTkJOEZ7Yo5xf/ka4DzEnMwrNCyzZcK3UJnukFAl4kKAEqPQJuTm
hW47ChN7q5fCgGTEQiYaBcIR2vX313+wGLwhIEf4uBoAUk9GzrYkIF+b27fEzhLIX1xStNWCocVc
l45PyZ11TnkZa9ZR3wJhb0asCsSShLpqfztT9dGJW5WJMAAMMxHCZCYdzsqkzaXPi9X+pJ/eSVO0
+3QvnNCaWkWqlEut9KYwAJLf8PsVubFwD1vx2+xzwuP/UDYKvWhu744Z10f3fQr1noZ3jIslBcha
nsBLolgytcAKZMRLh2nujGTA3UNhKgK2xtoYbDAZ5QIZHIv+6uRS9KRslDKaKNBm7TJORlnwAHll
ZVILQ1MZxbjKlbM03f+7DkP1jiaArVKahN4hkkdbjwzzb0OFqecLm8aej7vayrXsydh6ky15/PLO
TmVxPjMeQRFrLf411pgFlh9OszXdVJ+xf4nuLkfmZrsOZDk3LuF/REh1fPp8eIPF2i6kYIYYetks
Ws3qjKnJu8x2kf0/TyrpJwlX1Pu8Zhz6RwT/2t5Teyxz0RkcJKV4V0xTtkq9YYqZplieWFoH9Us2
Zea8gyvG9BepDDKnmwboUAMKhjTtgBmJbsEpIr+TDKbuT7vesiTDCrFHG1m4Kjb8fE0OHeevZ7MX
KphacIl6PPzbEjLQk7GcLps1HrEtPWjj9eMdXGluQwji+2vMsHWPeWe4YQL1LhUfUrSXTb4fMOKJ
eSyxoCDQ1hijAu4onQMhOFFIJfzLR8J8PNGRsRQU6EXwzmhBupeoul51DS0/XwUN2mQudLTvObeu
66QUTwrZAXFzP8kFCPNE9friL2FW6Arksum9DF0WvW2VQCwu4GmvPJtBbsy04QvJpp/wllfHuQ/Z
7ALdkxfuWWW/BwxMPmwLX8JWE8BpqU+GquKQSQeHKe1xvQUn2d4F5cQ1hBA6pQOoBJvzLyVexEVx
c9a/mqnM1eM7AIcbyMf4l0WrCjcg/jlXFYpyFq5CC8LZrTwQ/przEtUYp3JFa5G0hulu+ZwAaUlg
BR4KWAB3Dvlq1fmFcOf/Fal9ZAc3TYN08jnrWQtHt6E/mkZqX2AVE5lVB4eLDniISLUG3K1sXd0Y
vAU7n5WFVLdB/9LeN0tyvVoNusZtWf8hzJqJRNnqLyFlXS3fijSTnw7a3i8uW17fcdtCDkz9ONar
J+I4NGwieAuRBQ4cdJt2tp+EBafLMkytG/jCWhbhM8Wu2THhkOkR270e2Ds9w3wm5nLrRUw3mgxq
ePQeppq2L/aDMokdF/U/TfMgKPvXEAfPc81ALSSFcid41lvRkEHm4M7x+XD6BKw3gezuBBnE6b8F
lVV1pnR/qhqjpcZVUAPjS3DHwKurBR7Y9jXawo22N8JQT+jP3vwlKq9+Io92YWdUhfmggOTTAmwK
GJtGxDYLB+r0B/iae0Lu1RnW57xonJ4Ko/4i7QF1J+XxjkxOf+vAL7x8TZQ/XG/ce1sRJ7ih2Oxr
VSYJD/hY9w5+1R0tW7R7mIaF8DSa+qvpR3ntw+7dTfVnnLoRhIJczPWkB9LePyLrJUu4ylE3tOsh
2d/Oo+FPIXTNkYNqctXabXyzEoF6ZSXXiyWBC6a0tbtFHY92Ig8exBTZrrlTqn4pRzW86tc9aCye
sORejMJxLjPTyPnl6goIUjp9DMqUCOvoCR665qFAry0rO1Reazme9tklrg0WhhFx0cBd4TZEcI4w
H7IQ4tynVh5jccKPclvlMlILx9ZRi2NUos7pz15rF3WhvB/Ol8O2vQd48lnpbiLp8LnJ3zepE9dJ
/zqvMh4HsVD0hw9OETWZk+FOWOO3zrf0IcPhPfaIPtz26xtYoNyDpdxCi3inKPhm0ntAt+RsjaCc
VMEpj2+zMjgWz8XC/Sng1KJR9VVZLPFexbDeOPSdJxeNMy5Fet1Nj98SRFhHj8Yem6Ijau65GAjg
OrfcFJvCTQfxrAwrNCWq/rWX74vhjFM0HHo1FFBEMf4QNHhvevapTxjfNuFq2wqDsxmxUvf3bIAs
zSsBErXbUc3b5S0F/IERBXiRXxHmhA3bGOeK6mQcm1x9S693bG4fX31DLyXvx09iteDuBOs59ElW
ycjH1uyc/zXOxDUc5K6QZPFgAVa9VIJ6iOUnI9M+SIBYLFqpcFny+7hCX38df3UJS6GPl89ZaZqE
7OV2khrB6Qcn1+C510IQJUhm9fAJMNsDe65+PxCS3Ez9YApPhEd9WAdo15Huusjejd9pUPcgTMmu
762phWaSnTHy0EaoVsFaVBp19HXMAWo5cm6cjMyw55CQau4fLO1WulxPTp1IRQp1+ZYPH6LJVR5L
ICyBozLWbAcQIexvh/MfvTPdugV9N7a69q7C5h+G/bAIymeQMoxR1IlMW/BrpyrjvAPSXvKg3WsE
EOb2SkwH7HOphFgfsXiH0c8wT7Pl6Ots9GFkqNnlHTl1kWSycp32vVdvJV6RQlJ0WBFBmNNJmajn
DmeNRA7kl+3z1O2EBNtl+PjhFQl3TeOMaqokt7A5yYPAPTJsJMuJ3Elc/RjXn4oPdwEdEmq8QNbp
RIY2Dzn2+dwkKGTHUT+pY6mI8qS6+fHNE9VrzHqyQqxSZLF/xFLmyDdlqOUHoCSp3ZZGR7MwboTd
3+MXAZeV77xp1Kwv+IlI+Qi1ibJ5tNA44dHXk0b14XANBj9e9y392h+b4BpICsYI/pTyi6IZ/HuN
YVGDExgd1V/FUDKT41FnxL2tFRdsR+t1v2D/XuOK43OqBx/2in+6U8Nenll+rmkhXQXxz3f/HORa
IYakLZeetVBPEeFVAr2AiiOEu3R7R2KHEQlGIPxd2JfyyZkxvkmH/bkUqTlgI9AVlnWjPJPAaKNX
SuzHOZBXk+FyHans53CcVYHaMgf8mdsNVlE5NHsI0FZ9Hi8JoZIwrKxRPY4qHwv1nRsDZvKxfX7a
Rj7/E7oMsxm+Zr2oNivwFjCkAMqOdYgDFsp/G9o1o+Sqyag9rSmtNCSFcuQVxRNkcX2oFfxseVbM
jbYhFHnZME0zxE3h6sXzklNWzUAhoEnEmH3WK2bs/IUYji17wmE0otY87jESiSMVZ2ENJXg1DA2Y
yxjCIeAp+Iq5cufapxWdoJzUKuZEGVwIOYwmMBZnjhNkXjWXgz45RjojbECyqBUFl2blbKbUyagA
L9Db9bvocepPDP/5+LztsQ97rJKcvKsiu9LRnbdgCg95maT9d8Trzs1fXBSFs4gfEMXz8X/wA66p
etbU0gh2Rr3XnOXXAviGoVHSsHWtHhvcG0prOhtjdnadLjKbFkAipknPjpWUI0z1lAz/gKC1e3SC
BrvWLrijM7IyonTyCnA6gSeyTlpOqQUKdxgggG/sPdIcnbHzHm/XpdJd8I5MfVe3L12YJTq/+olX
HFeIWHUm3eQz9X0LNjSvRvnmqAp3Hp6PCiwNM8p4Pqf+r3orTCw95E9VRsyfoAD7nTGsvqevOHgg
HdItn87veaLGevR2Amn26FWI4l+Fh4ARoMMINop4xApukl/pbhEesStBXmnVHGE7M5G8BauFm4CA
ofD21Y5nRguEK7smQJXvVAlYw33H5dymtr05p2LVzfDf+uTV0ipFjiSfKoGIGHpsd+NJbYouLWx3
DrPFYkkd5nXiediX0bQiFQATBNOml53CxAA4xoxzYKoYw/wgE7/6YdlQBo9MJ1RVMARbpMGwvQID
U336d49SF1i4PN3hZdmVLfw6/kNGkcbTTlyXN5+MCVc2euAgct3ul2d1s8BnUzq1Yq5X6CmvM5IU
V2cXY3jnyO+SK5BLsgbgx91h1eNkmrjApp1zMtv3iU1XxD52exmrBkWqY/dy2tvtyyVHfo8xPadK
5l1tecHGIfPlNdWn/Jo7Ll0x/XI2znaUyK7nIfYpdNI7KNh7IlJ9GUSPWf7758m8tHEnhlkRfMPv
0cWnpx4BLtNVrwicnjjuRcNJMTFKcwq/4Yu10GGjuOJ+gXrsbj1T6/OHlOXMgpPxzuEObJJ2FCqx
DXqsF1BDbbrCoXgn8NEgY1UaRwh0j53mXgOUVjtnBCqe2fAWh4YK6HWkUCQmddU26diFMG7tpkoV
5MQ9ufbgY9J7KCvZAL0MLPBZWQZ2NdhRHBEeGOj5vN2ksEY/g/P8uc7N/qQVDczB0Raf6x0r22nA
tHwQE6lh54+NpoOrza+21sEtrXC7wJxlH2Z9FjHDDCVT5UUJ5HmqCR9C11+khOXghsy75nNcT3Ce
JHeTdsEULn/1HMugPKBWf4eAfaTOTVq9mVFzyVreDREOdvsKd14cYR2yI+Cv64JBUtKnU5/7v8oe
/zEM8hJ3NEYZkI5Xm+XpOS1dz4GGRZWBLhOLJNrBeIIwnC4pn2qde+uNyWw1bqJ3+q0WE4oDrGQA
cIcxteXw+Wp+cBIFGCCnoMiI/JVuSsaAbrrVXi5BjLWlV7hNO6VqJyqb66xHgOvKLpThzX/CY33V
sORMspahqet8EVX11L3Ik7mux/HQ0qPF6v/rEz1TJDoGljBkkaqKnzZ0lCb82oZiCPi3HBTK6v1G
xCjwkZiH8dU+k38k0gafxmu+J1Zhh2yJnMeffT2zlgrTPmZuTvn8fH5SoEmF2afk1oDnI6Lv5RmE
VH9JwjOrAD83pCAKcbY1J+/1GD5KuGMkDWsd2eJPahJaYvC7hprfjuK2rjxKZSQpCzSZnxnCyHZ+
5ArKJrdUJmy7RPTwy/nkRQJ5EyD9rHq2dTp9M5PKvu46fuxOtixXYYPciEhtMgjQOtfly1Mb3BL6
I0FT2vtds9iYpRrNv9Lsbo9ejRiVyDrck5PoRbvAcjteqHNeE5idP+pUI0/h4tnbRaZf+5QCCvaT
CPrukARZBVbRLwKKGq+QJR/JAD2eWZ5tSRSR8v5QFGhuIS/stVbCNzd6Xpx2bxtR12bPkGJEX5Ys
kINq+WFCpen5BAuTxhYU8NmYDQbd1OYDcSY7NcPJaQ8L8mjzcBbeoBuu3lTWLRHEBI+X+BQA+t70
1r33Tf1kzT8RFCKYZQDZvlx+Zr11Q0On6ud6XTAApn3hI6RrA77svVKlP3XRnPLd0VrrG+ESpN1n
Cz6zeJHAR/pG1lS88NmeVQsA0ayoOG/Fmak7ka65t5Yc8dJcXarZGRANNlhFgtkXDEhCgUXHY5I0
oUNuAsgJLdZ3SRfC3tpoH3zHAZvJ7C+oJUbYJbfuJ/oM+OKLX1b+C5Ise51rHUA7PRjql+IWMMAG
nB8ixgclZTChT2mz9kYknPuf1vFvwdgNtkQ+cVSz7FEWLlB8i90d+yFJ/baKzIeJVreGsGv8lqDu
cU0dkOesUj6W1PH5DZyQpGz1LXlqR68TQ1qMJ/ojyl/w0GWYBAgYGnEGr1vjolxSNKYSCsLEhNeY
Ni1HmONSsNL0B+2oo4xW+zIFxOZqvZbL9vqVBK3LEDaCv4vguplmvXIcP1DZlmqLIghn4zEj6MaS
V3S1Y69LFKNKBJri+I9/tV2DmF6bQLrVwLVCGW//5C3WyEbx/FUMqP7fqQhCUhZlTncKZSOj2oNc
iNdhqpJuO1PquqSg0jyWyZri29GF2NCubF9FE7mXE5YMoflc8xdgCNGc0ktKBFGrWevnJDgMG7+Q
6yezXhwVWKNiICyKacxKYn4t1F73UhZh/b6A/0duBmb0u88tedAG0HCOvQBqFpegjcEkAr1iYiBY
vuydl4ltPJAH1QjwcrRCEnLknLBDC02592yqGwbdb+E/R0mkzgsHY0FwGdcZp54HRob1h+DaJXkM
tj5sXJwBM9iok3vKfZPKN+b6SnRQ6APxUMOolLmIHF7J2bzS1YEN7M1OwCEt7WkmkJxMMqwbm4E/
lH02P4lpJsSZQYwGzeLuSaKTtVFJFMr9jvDifLEDJxEFIdutcrnAWv35ncwYcDLl2ivqPxCbK7r8
YAP5EFLO3V8qKEgnR9QFY2hWvdj2t0gppzkSU1X+BtKI7E3DnwIrTPgCn3tZC9gbN1KLSqIR/GG+
y8jv3WfomMDXxlNbz8fy5+ovYkQH5VLxQWBvyNdSYP7xUNp5sH2ukd7kJUKCW1qogo2vaHFWZU7j
yNzuB20HPLt8IyeGrIY5RaL3TTJP/sjfQkbyCQf7u1qvyfz6B7gh5vDf8W+EaNgJ5gnpfsYvbX90
6i58ck3Ozi2Gt6tdzo6vjPZcGeK1SsPQZ+8A+znaRmovZfckyixNeJClhsu6IUtGL6zywiBu4XFQ
s4yL+QoODWDdeULcIzrslAoYGyq9kPsJXRj7FLNEkqjbZN71MtS/gGXu/S0CTqX+WR68AK9Ply02
E6zCz/NmwehruyVkhi/K4g+psDWJ8HG7/mE0gDOzcVtX28jABPS7j2Ts/UEr98ovgK7xxHBHhn1u
VFaSsY26jKprDBmybLDvFK1YdTOVYNjBDbyu8vah4TW0Wn1DTNTEEV/grv4xRtx9kgUNrwfEwMRf
JaV9cSVQMH9T1iirPyFLJqNJyje/1oZ1BbXL0lgTFDgt/jvHQU5G73rzhrj4uPOkISvzU6JtcvBa
HYzHZyl11yhhi84wahmArswrvIG8X/LDvtJhcRi3zzf8jlL9CoEbOogB/iN9TJJ3aYwSjOowTOln
RXT+kg+vL+NTr0a7KxCld+PE0SK7Oxru4te5Fhx8C8phxUcgrWmeKO1vlKFyoO2EY076jgIwORMq
2SmaD9q1Yub7vNttLm/sPf7vw1ypU7q6DmzPEekaj709BaV2LulpLVM4wBcW0Xnh8biA3G3ZL14Z
+Gzn0NIVTJf8VIwwJFRydBxhGa0qQfRagpKuS4xj7/CFi/5IE9OdsnC5fVJc71W20GxlnX6tWTRD
aGfMqofBQh38ooeh2wRrccrfztXzCiZ0k4rG8tirbxzM1D5YL8Luk0jmbyBv1jb2TTP8BDk73Cfv
jLTEEW7DGTheaJZdkz+dik9x1/vjRq4A04UmNRFv8T3nDX1oWuDDxxAb5f6lX3WnKHrYpndTdyLb
5OuSfENxcHBO19ssW1q451Woq4MAqUAUijx80QziH/LsDTmhsd4JbB2vyIlo4q+KNDV8huKXkdM7
WBx3EvBugVoBWiw6eRsjMokOdvEckPXnBNFqEDFuBot314MpWTPw5j2knMbjA9lLh1nBJjfn2FHR
ftPd1Yg5Q8RJUN8TzQGXxhQDhRJS2nLVYoKSQFWvPJrqsd0OY9Nb/4Cds8ZQNW7FOSQFAzEmURBb
hqN50Wi/74ulpmZhdctPYSyhe7O2a+7Hsr2GJVg9wQlGNHpla66OXIY+WfBH+PLJQYWch22RR5Yx
GNV51NpDzxy/3atD6rAyV6CZlL24GA5YkQ/hHOgxTrqa++gwHSS6/RA7oC5hLvLl/gkw/eF1BKrS
BZncR5ZMieeLGwrARmRWuFBlVqhLFVAO7VT6aXdXlCWdPJy8Tq6Stxm0ju3z4HgBa9g53AjwCjZu
X4l73ca/AZpOKxq7oZ6jqFdToJhJe4dzYLmLqjAJr4GPko48YhLMB+BIWhLG33SSoWHMD1EywiQ9
rGfq+uVUNLMFePFUE0H8c25SzFfwgdCLyp1pKpkq6KfsAkk6ZcV3WiVYLTNBJ/yCLGBzAyB0Ea0H
QUw8fDoEtGykfXnnDY7UPaaQndtgANiSDjeHA77tHW3+F4mShTFiBnlM0TkEYl1vuhHh1JeSDNhX
mA9oqhNVUxJ9KvS0JxAWeUQd9t9TnQYPlL/46t6odoYFItpEl4yQCq2s6MSzN6tRZW+Q49FzsT3x
CTEJfz7gn4qr71Kn1pNXAinu3sStk7lYDVhgVMM+q8CmtwNZGNLwSiF2CxbBprFPYVyuXZSrYplR
XZ4QxdoA0l/WiM3nj0XW2VjqUzSc0J/nmtxOP4nv3VQlXs9ardwvundSyAGwuLLFlXvT0XSKEx2Q
Zh5XaLtPTz+yNchuqVUlCaZkY4dB50oBaocF/eOvogOdJinZpPKN1iaUf++kqQ2TRP9HfsaOb84D
/zlF22J0iQoJ1/dwHTz/P/T8PiASNESgrLSzdoiOqH1GwcVHdbN0lQgpdf5m99vKKwQeb6Bczmkk
WPwUVSNTNoEiwVG4wK6hCaPDXimxxm5EpyGxaf0WzKWSZYPW7J9SBNrI26e/KSsZYfSwSK1dGb6J
d4nDe9Ot2AKkUS4TRh6ikPp1A4ecy78t20PrNBasHWja8YCK/8qtWo/oUa16vYeLEgkzLBjz+lWU
gdBYsoi7yA9Q3+qfgZCSzl2vfhmvYzm2VFh5NaiWyjdsjGNvDUzmjLlV9plY/a/lpDgB1OzsUeOF
6e/kNbcdxoMVcKlpJtGLMFwmaszEWdK0XLBL8MsHf9iOwnDK6ZVnkqE0A6Z5DH0vbt/L661U0+7P
ZxR+0ql63IKM+TjyHAF2DNodHGx7lLYFGOahPiwP+X1259q86qTKe7c0m3xF66h05/S/ySTbKfuA
w06Pvt5NasC6N4LldOm2+mbjKzZ6avrpozcsbFGvosUMvHAbgB1hF+qWAdFm/k4wESGtMLGHUvnH
+3uT5QtuG2pHxb9OiVPyjoYsWq3WCEh1hkgfCyNqQu82/lhVCs6Pjc1UcY2jtDDKOra1neg1JJdg
P2YzMVzUGVDYjlKDHXkjSG87fOXv0Wmf6q4NIPvS8lnQC8fsXcNGfusmZtfJoU2SxuJIrARYR3gA
sGUWIiZJJUu+c3BtT7nRkJgGv71qNq4TaV2v4xy7Hiec9uwXJexMv4KAtw88o6kNjTNCGW3rpM/9
svs8Yg4oQJ31ZJuNcHvl/iJB9C1pQ9GBK4cPZvBwlP17zni+gcBd1wDQdg8ztHEddK/ndsKuzZac
o+TsxTtcERx26UJf1leakseQmDAtL+CtHu23UyRwWJjFZeWF1Rh8vEA/xvY1OxaN7I8Sg/VFabrp
D1CH7kERgaExCy8qTakr7SB46DLUzyqWctTdGlK8WCwO/8VLwuS1jF5zIMsYIqZwi6ca+Xt2tv/8
ohLd+7+VUZnn5yIgIJZIJU1QjFvvGTmjeBO4AIZh0gO+tI6uV/sWBqKw4m7yr6aY750XZVStF9vV
itnfN0uJvpNghI1YAx5fmN9GvSIfgJBdLAP7sCwMxBFxsVg8OvvsG8VlbhTqrfwrB6FOV6X0jIM6
Ewh67/LDoW/5tnEeh55Z2WQUC6Kd9IYCGwDpNuWIBUxcigChVAZhc8j0u7kK0EBJljneK8eLMWXo
MN7ZinU90FjbzAMipbQz4VU1VqsRxO1DcjSHxMie8QizYXzywfr2QIewhI6SxtzAo4dpP6sgNQFn
er40Rqy/lL0VIuMeOEsCQgo95cMh0eM/3JQzZFzp3mzuDfh79VxxDh08S+4bmjTHY8rwQZUqLoiB
r00PlcPcgtXVr3a23EpkbBc4H5AJLldRZ4qDAfR0O62CldDzxkQ77+ghxr4wKEEnhMBfoSe2edzV
ygV2aVrGMB4iG9x371wI88o4z69R0/So6HXLYDoG7x82uQzySrMejLiWEnp+Dyvw1GJDZYKGFjuR
hhJ81TiLJhiH3DfSjpmfJyCU9LcuWlHBnciXOMiUFUPT/6fMRx4HwTupP00X6MKLRwm/OOMweBtu
UiiXB7bVP7HHLvfySj2d6Y+DtucfIuvpUlSDq+rIBfVIJfCGZv33kjQGsS4j/fqn0PIxLP1FsHah
UYigXCPZ7tTMvL4I8AcUk2okVqjhfXvE1+PFxHIUlWyBVA6LXQ1ABrvTb+5ObBDkX36Td7x84kL2
ODqYMbzEAssKP0f3Zq+b0YSJra63BbCT7sqTGmUUerXoa6kVBiXCwmadOloMLLOEKQJ5QPbSuOp8
C4Nk3DKjFY7XGpvUVqVdS7ZgbOIN9Jplx8RVto/LAzEB3cldP5xdcDBYrt2ENfRqERyLm9hN1YEY
fZUAZiXXBpjBwlltuM/d3nxBrjH/Q4G3Y7+iOsxDByoQgMrApg6UBobmHUzsI8hRqGu9dh7ya/da
rpXQbUIcv3z+v1dYq+ulNKrjlvS8R6UpyU2Co6YZS0nrbu6eigewooOkTcYQkidjhPt1xWcYXetP
LEl08vZU9obmfAmvCfZ3uTUNFE1LzXc1FPZVQRInVkRljAUYPnljfEgqKWvAE89mZeFHd6QgbF49
HL+AcMGt9Ez/bPxzns8yA8MqkXnq9KjeXB2QOT2oGX+6NH/X6IbfnYwMHcE+85+OVpt041K/ISxU
Pbz3Ce5qqXVLZfGisO6i1dtvouVd2W4+k+ApOdqk0HedKOPvX70WSFnmiBNzvgaz8qP1wklqa+gB
8zR0jh68i5qYrOk0Qu+HChGvDjwcNApQEQIvGQe+/6qwZDgJX0UQCyjnISHBi0yaA5kpmTkaFdNa
6uoQ0LkeR5bMS/Uzv8bSKcgjav8WB01U+gxyUDmwreAaZD2SICDiGPbsdmBiDMhe96J1Z9Na04v2
7RRvuep7gyZ9wOTycOFprx1wAIm1ywrVAMM8+T0OWlCLMMWPL0sjB9yAdg7nqqbjRsbIMUwtsBVI
I19lRho7c4e60wlbD4WQSFAdPUkIw7CZZUlA3t0G2AWU5NMyNkB2b6n1rf9xpBVlslZ1+OgOvfQy
nZeR1x2WrEHPx8sI3xJ6aOwbsAB/0SasUeBO73NS9EFA6KyVSDNaDEUG5zdlRPdJ1lkG++0W849s
ctHg8GsggYjFobo5hz7Dij/syIH8X4AexxZjKn+xDAn+vcdjbdtv6xvUFHglj28TwKxmHCIrdu5y
dAGQ+0QoHjAt6pbgE/VOecmWulIW0a1SX4v7q5W/8LZ+GRH2x6SapoOuCrdzhUw0bYZQfDkSiQEo
RarKvwk1VNAcziRHZS2DeIYQgWRUZvXf0QH5bJcTms6iBKuSKiHye7ytGvS19/mgewbkeDUdwz12
udeXo4fWdHLw+lYAcr2TBook3HJXxyut+WjqkgKqOALWBJ0+BNQ/b+PYSsG6THw+kpEinmZEyvr6
zkDb8Ha2l/DhsCMUhBDLDxSjbxYTGwQMM6vAY00+UEPL0aOQBXlTLemmo9Wq0WFZuELAv8tW3872
L8gNcpXeTJaaeK3UxF8YmAj1gcknHlVzLV0KYjKNCIiZHWIi8dlnMNzWL9kKWulFrVU9+Vb78bOc
/6455fX0qOkfSDwfiSjG+gbIliHOT803q33AaOdcFGVm9fMd0Kc8VcvGIPVbuIy3CjnaGBsITve0
jHIuz1rirnT9ejpbZS9jsDVFrFBfxxUqa+PURsJroTGgpMps6igGEbWLZunrvHSODYs6jIHdbNRZ
w2SLbN/w1y82MSMHge0Ww1aPqvQzLK5mzQ/RFVlUoFwP1tKpW+Ur9Bd1wYrnoYMNH1swtUJ6sLLD
8ia0onC2+ZWd3GifoFPkW/7GjxJm6X56V13i0muFpbD+PDWRJMR5TQbMaq+JTwYszF90CI6Zd2l3
hh9TdvjwX/sxwlvYr8/RCPQjpvaN96eTv4i4JHl9p3tV3EicNaUdwbp5mVLD+v5Kzx/gpj7ZAN1y
/yIRshpgnrZfgpxoiVS9SqjMY+SaKvSlP6TRpu3WB1cQiTF2nP9Mns6b4UBtKEy+DXvm7kpKqjG9
mQgrGb427VOqPdxXlpjeGbSa197jjrHklc6VvB4w7YDvY8U/Ht3C4HxVgKw51FkTM503CExqaF0z
QFDz4oHGTqe7jGgeYX0LD/mz5huaXwkpcH8BjJaaY+xHWCOmlwBb3Q58dHKNcVTCBOMbhcvG4lxU
7EoIXZE7u0ROZbcQsXiciKaSuMkBL/ZHazdPsnkbm1IJ3I86VVJFnKnFzwpv8d8sBo3KBQYirU3/
cIrYBkriQv4tvE7dpYEteaqa2JVIi4QelBssVdJTCAu0nxWlfAezdL1oA1D/FdMF0FsfZisb63ga
Am/2mUnTaVNSpEo9mzsZH4ZK61ffKwDwxzxxFMxpalHucED4707RcKCgYjZGxoCuSa+oRAxrcv17
nAFXS25IzuE/SkIInf8I1CI4IgO8ZV7RI6xEJ7krMlbRIp0z9gYeBnWqIyRMQ4ijTW0XRtuTPkQg
Obm/jrB3NzvusU1gmPIKDjPa44mhm+jQTDb0YuQrB2QShh7W/5L54tdWNRfKF1BcR83oddCN5yZM
Rq5WGhfjgYFhUcYSC21he82rbjt+7tk0l2I4smrxCDu6erCwKx0KPqRKGKJazaY6fkGu0tPq4//F
kp5wFNCcdpC5ji3olF2Oa9wddfhZIFgV53C7YBQ/uDRjV4v6xXQQl48FrO6ca3NEZzhsY6VyNS5Q
agdlcP2qCCAK1c8tb7yPnndbf20b6VBiP8DhbdX54uA3KTM1eRjKfGFa6k28u3WSrMuGWIDI6Q9b
q5w3NbRQR2AGgk1Bq50u/qE12ZuW20e9piRKi6lJGDV7w9d/zNnKzF8HrUJmDteAGzqygkf40Llw
EFJyqMm1wcA5/fbpTg4+I5Es28jhVyNXfkL441+UYjdjk5qc8XTNOdrU/fNyukHuuk532DljG2AI
RWw4u4W3h1VkWpEnffDvnntcfFNH6IRUbwQTkPDqexlg1IYJ/x30f+3PZfZsu3HE4zk55YBnp3UH
BtIJTWQZ6ISJ/Vh7nOlM6ixiJ4BUyXtze9wH2QccZFl8qpKHy/fOPlhmK/5QLqsb2gsjZqX5sFkr
XfceyOwYH6A/0VLCKGN7vzjQ8EvMFXeWOAmx5WZWDHdR6VW+kOPnzircoIrUXOPLO892nLddBFBM
75pd8WhddNTcthXgOpz/fuMI2PIdXVtNhlgifxuNtWi/ruzTIamtBmLfOQkkbExA+h+3wcuDa5bf
FpCXMPv2stVUmEO9pIlEaOZk5JhE9AjwJKE3Hg29gtNPhkqLABGEyshkqFn0tAMGdR8SbKceS1fj
QnEz+dosbuzBob+OLQh68vRak9BlxJhsSA2ysb51Z1gs3+4nwgO1Uyn8huKfK0IK2jI+oK8+j0+E
t4jPr7xb/3zz7Z68Z6XrysC7dU7W8CyYbiqBJq7/qs4HPnham5UnBzGJBCY3vzix6kUDRpuRiDeX
jfh6MA3H3pHim1l1S8lmbDckEkhgUPiiHw46Su19me1ahfWWB4ieAPx/Mhd98o3+EaH240byY8km
hVk/sJx4XMUrzfk0Vq6q3iaKQElAsGMQlGD7QjVhUzltPbelPfA01sLQOvE/Gp8nqfzYeCr58uB0
g8hrStNEocQLtwE9GZpkpZzZe/lDkVRYe2qgqM0m5gPfVALkOEgkO1w1k+PbUpJi4vJerUcCPV/+
WYZe5mblB7QxCRMv8850U9s4V83pDmc57NIlMgsv9x/080FRZn2qBPeUsKrVKZ1HAbcGKc6T1JMB
WL6y4z9bAh34A2msqIYHmvLCw7054qM5KtNjPO3EYkuH4xKFCSZ3KjH2KFG641R/KXssBhMcLZgF
dQyP3O7kE0NB/1hpjMpihJaCvU854FYjzN9ENUBYQjIy/FfW8btYP0RgpLaJlf5CbrqELGUacLR3
z5iD4J38JV+8V/PBUk+QQkrv9BRI1t0MUxEFW7df7Ywu8nDj/JH2jg8JTeeABQptbtAMBaiHgWc4
GFaU0eEKeZ8mKUALj7h4x+bga5+r5kg0FiXIk6fr5Z67C36v/pDvVMo3O+VIqtVw8LIvWp/QuMQR
lwPNunA7v02Twjbb62NG+nok460FZKQGrX+7yNieWVWnb2WKAzmKFvNRBRY64IJDZIGqGDJCIU0E
vVikFyaKVhoP7t4jvsNrmPsObpj96/6pTIceZPb0NueHaEqim49tLRBDU1r4ZmNoSFbzyPI8zN8u
HOo5dnrEsIXIgp6qEDTpEpRIAjvygxlovXOhCeFN5WkW12k3r/o+qDmjZwQg1GPHCbGK/ZMpPFEa
FXJuIEi3Uujq+aninQfOCZVBYUZZMSadCWaUcMc7R2/KuzyWCfr52Gt+EmXv36LNzXasp0bKzG1X
Cl3giDcgeKfYSiK5SGWqCQn6ELFRU4eaHtV8O944uqcUpdWkynWHXHXg5QtuT3PvooeVZTq2lWTr
LixmNfjuOXDSTwtHgMJqJ5eNz/7J/yzfBGb27baZsubxFkkANgp+HMkMtf+LTxYl4DvBOnkBfpkR
aY8s7gcoka2Ffzut+FY5SJ6ASRNwOnahL4d6RLAw7MbQMw0xzIHZd981Sr8g6Z4N6SP3O1m1W7nm
VxM1qxIGXzOC6sDElQWnV+sNyJN2Fh7+Xt7p7OPsl4x7jb/cDXadJbPgTYA/SxdIO0MBPFdYm4We
cwoa/GED2pQioKv/n1zlmFmUWLu1EFlQeYlV96c54jpuZhDRejoTKdQJE0hKDWoIG0En1DERPWf8
kYDSnHbYJfUEOxi2wUoAtosXYsccbR0La3aB8d2CiyhVBThCSdGn66vGo98D6jow0fGTZvPbi8fb
+gwPb5aG5K+GzVwcb74s31rd79wjQuexQb6TJjTQGcvzcevd3AQjutjhmIBKTy4VCIz16Ox5Hdgz
tHA2zAUD47oqu7THR5eLm9Bv3CMR+yCDzvVFUpAW8JB2vGHEyZXtkmMKpNTnuFdX1M4YhNK/eNWb
mig2rzzDuBQyKFEOxa06iXLndw8xD9AefMgQl49/J8EibHAT1RZeyehyR4HAMdtdi+9m3HfNedsP
SVvO3OgMgd2P1JvnId5YDFdP9SkMqHvOvBt1SxVaaFHGmbEDzAXyUI4HOVKFszzpmIWSoGezjMsA
wroFl6R0Kl/oQPIiLkM5m93WDp2A23JmsznpYHxBPDgdtIcQVoDLvsp1yYw7Vl3BofqP+adR/l3B
ajh258vB7BLltgD47EY6BL6debFfsGcWCZjH6lTeONQPNzH2+R1JBKkcYbOKnaY4tGvQTc4XMu9w
TudQ+0aGe147ZOWZlVPLjG0gLIpuaxclh8dJ6X14r5SxbCvm82lWFLQX5H9roD85TnfcdtcSyeXE
uR5/Xqwue5DCmUxaPgueojrMF8gHaS2+yZ9Jup53KMKfrzR2BcTIW4oZmMpU7+gR7em8Joqc5po0
J4x8FWOzCIWYvtKjpcikEBCtFp2Qi+KXpDlA/NNIUBTyHKIuj3dJ5LuY0puu1u2RXRDF/GKqLgsP
qWc3rr4Qyubmuzsugeuowi8+/LREpSrh5VKoffvMD5F0UsZ2qK0Mv3fxTUdU7906VQmpNEoH4Knz
Cq0nu1zB1zwAI4FWLlDkF3Gsxcx8KOxv3fYyuKlwB50/ChGTOjcrtJeCIDHWcw/WSvjqGz7T/Z9o
ozidQAX8z8NIFxnyHC2M2rtz1yTSxSPkaV+ttGiOUFEeZUCVfr72eilo9H8cayTmYzzBi8ioLycU
uCJP5ltksMc4Q5nEfEEnHDtJqR8r6OBjbqoYI7iuz5ePy0UBNwJdMGyqv6SJX6And4f0hpw5YWeO
18q+q+B7D/ZYhYd66wSBIbzjTWf0lMYEZcj5/juzR4+Vd8JjjMv9ZH4w2bfls0YVJocTFGrOzOZf
1PMTxdHJKE4UTT8cS8Uk7li+3Q5zjBK2+hAn2MLCkGGG4UuDuOH2BRkdIIQ1KDvi95Em2jVxLEQr
JdfY40G9UGItg75JM4RQZj3Ey0Z+W6lkQyMQRAlv3CBdCe6b0vBaxMLLFPetHhzUozySYyoJpxjP
ziWTyQTNkLm35i9oKniFW6o49DQttbe1j2tyn5z2m7V2+zVcP47kkJwFDOG1SoVeKR/6dLBuJEv+
D/ahZOgJw+Z70NzWsY+1z4O7BAwrEyAfY4CHDukUCYyFnCWPYtMfyrQ2rJ4MaAL70TtT8bS5a5j0
KVJBakWwOvmpnnyy0e/5H6Wi6rdDoEKUtMzM5F4BEYH7PRL98nq92QrMW3eLovr1zJf42n6P94uh
0JiO64iCMj9d7pHk2VYTDsovVHag6I4Yryi2zsdFpzXscpbIS8RmNECeMmZPUUJ+0+KRk1/q3rBP
1WJkHLFVAe84eEgNqSKLeZCCh098k4HYUXGn5C5dplH7FAjSYAiXGT4F1GtQ0n8Rq3o76Xte1TKA
8Sjd8+IbCpJ+tIa+ig1bTPmJ/7tfWPrx8B0eFbgZS8Ot1ggWAumuo8m4Qnhin2TYQPt7NmRPb2mM
vS9CC2J/6qHNhdNJBeONyCUsZC6XERpsiCbHv2MZuUfBDnzj6ibAljWZuGLo94XTa5kc5BJaUR8m
ZMdNOwgS+Jkh//qz1RdOLEnflTC3czf3j256pV/v6E7CEnFfEqrCGmIUu+oVW4VklcRvRNSrJKoD
aoszOSmR8bFU9A9YYWs9v4J5/vCAmIfJ/JCB7MON4u484NsmNfo5BN8DoI1+8L7dZZyUX5Mpfw0e
YI+3ID4FHM1vz6m48I34MQuYCPVpozfCPnCpZGjpgtIzPRai0Spd4I2EwYwmxy9uVZaFmqo/Sg1X
I4EaJO49d84gmd0q71R1ufzAK6N4xP05uQvkIAoiHkoXG0ts7mzrREnj0XCKnxUKVq95mS0S43ov
qXp7vS+6wGEx4/DxRYoCp33+jTe17ypfoNcPpBYU8FI6nUXsOfI+2ED+AN52LjyTx7qJpzJe8gjk
ZqLkKEUeIwUaJsgUzyH6Z5IFjMcsTKPD/p1rMjjPoZw5zBy+9RmyatlhnWZLWtAlxyabOSLCjKCP
chSDPcgOfpRI52dhegO835rhlCyXLXTrg12yX15tLE2CnHanKXtdbemg/LX48+MWTntIhb6qq7J1
nDdRVb8H5+dy7DKCE8bViqJAM8TVx81THOO6pMFVP/Rr6KPvu5Ap7/FjmLX3/cFoWSJBRKzWpZj4
zTWmZE42GrdvShK9ZIOMW/OcGiKLQO/Hmvp0eQxERGDyfirfHj91eUABHmhrwe/PKtmo1klkeUod
ogxrIhACF4huVXILmWwkyTDbjgkFhewiqYIvPYagMl/iT8Tq8wtkYbcwWBwEGpIEiDQOt7jnXCQi
2aLnU5JGehXb/scZSUNw3EA74Fc8NA7B5hxpJf6++P/b1/7DfhzObu0T8OiHi8SmRfqfAqXbl8//
199PoqPhwr9Bs8o97cmg8y5oEhCgPIOSUgxDZevGh4D/Z9r1oIWYZR7UXGq9G4cDnTjW+pNCnpBU
Ei6mbgcTJxvSjuaQXKD8iMvn8TUx1KJMtINPW9ePh5jBG5teKv1ldMecc+h/wWREhcbgwzYPY70o
XOGFudVWSMo0kb9ZZ2P7vchMp58AGMoZK1NOxnyYchHbXQN8GjY47INjPn+jop2KcC8Skb4BTW8V
7AEpg1ENGKsl0LRrbc5Ut1vybD2DtNZ79/kKwts4r5p5CHRF5zZcJf2jrnNPR1QtYdx5krSuztEM
qjNb5/sNNV6+YlzDzswVFInj+H/qOgLQuFXN+T6GYXGfZMfRDX55jTxWw1/e8FDI2rw4fW1syV0K
NlrxCqBLPGv2tnGhRMXZqrJ9w/oxYvetKuOo1yElCjFpLxx6n6HBOQYNArvr4U3Sig1xgKyKYZET
oXCXPbLOq3PmGfjnyfYwSu2qXQkwuLgpffGXqprpK9hn29/i9QXmUjSns9lFxbFmJ80s3ZuBBJq7
lg6FNbRNGHmsMA5VDNv6lrIBKrTxKvLgBr4G4vUMvWSLG5FukmMTVyPkswbajrhF33Y7f/lS/LNp
XG4TwSVFsQngE3TvUAV7mC4c/gxlpMh5oZariNg51JrQQpb4NtXQdDz+uKH7hsjVWKmUtegD9Ynr
+3kjOm4oqdNKjcgyRRR96bdu9JMDCtvhCcz8ZvkPovEXlTXWFP8g8eUJBg0om1Fok0A0KqGXkOWb
sZMHLjwbYlVtWBoH6wakMW1QSYrepSnHvHCOPJqp+m3HNv0k4R2tB6c68B2t36dMxUOWpuYMQqC3
djQUnjLKAz3BYCIiPr4FPyM8SJzdn/lewMIZYCKpajTXFriGAbGsfcoVCru1cSivHkI+ZfvLxAOV
87cxc//U6vIiFu6VN8OoxpWch7bcbxFWWnFsIFCTAoPNewcrBZxrEOdp140ITMG7aCeDh63q7hWU
mC5KtgK6GQNjW2jBvqV+KiUgMuAO4GX6Z/ticPdh01Me5Ge7gz8ABFTphqMTxL/8+BSGbzOz+5LI
lb1LAnjqv2c6pLCgVUqQRImk8El6MeFtw7YAWXpNQ0hZaWr2+8Td+v0y++y69d+0cJt0p9fqM0N6
rbpTCWXRf8R65i1W1md30lcO20iuLX0N4hybcZQKRcdpVWkmpLw/WSyOwypIudln7YSXnNjdkx2S
IcpBu22FS/3clGB0or9mKoFMACLlogCXMVSnV5Y6J9y8Ic7PDI0GW1JeULO/oPU7+6n9WTyMbGfc
wsrvniZSN2DvNRVVvqd47uz098BE0KnXS6HsjhWYn+9qgw6ROLIdXmZWVqDmtc5jeAgBngnLnxvM
eHucH9cDuElqYFaHjaSncG/8dOsEVFG920uZyVz7wg3NzouMs0XuoQ6IA8hGl/5avk8EHTzueUGL
lTJbaAW+33BkbyDOiOORkVpIqreezpVCbl4Y+NoBcjy63q+I7iXEXNkkY9PJTcAQVzB/sqH+MxF3
8F3zm+2uY084Yg+J7NmORYJr0W34y9SrBKHF3DUhucpzOcpGxkUmnnYh+VG+kfJisLP6Kv4MzrR2
BiT/dJOTtR2wZtykwKix8EE3cB3roa6njIBW6YfmayazbYgTj7Q8v3Oke9UjTL5roZZVl2+N1Cpy
ISoYNo4+Zb/VFYm4Dx4MrKYeE1KIVBdA08kJRi5Cz7ik+vbTe0jgyN3nYRzKHcmffbzFDMb91PRE
gaaR4Uhede+ISuu95SODqc9G+KoCuDHBScq/uKBC2EmZy65nWJVgtJGj1bUxYVoe5XxSLRC4OmjB
dRDTkCx2Z6nxJET9cui5vGiVdZlmEQzaI8O1PR6mg7bT5+xIj5NEbYJCt4hfDdS8sO/Fwkebd4rl
Q+DN8HUGZOvRpN2GK00ksiVuOooIwlaRbaz+kvweoSLuMIcUPwnsCEJEixloWg6wJK+74UMwfyIi
s9lIGFtI4H1TpxOvCh3OXUdgPhQd5Japudu05qADWf7FSd/eDuFR7BFXzUUoQnbjrqghov1eGxU3
cLqF2+INLAcqvhQyTd1Zz4CHmPO9lBbcCEUillugpm/98K5TUqXwX3JCpl3BsGUtDqZiRoXtk9h1
+eTedD1dxv1KclI9eLnPKtcpGcjYqBiom2O82uyjA+M46wfa35S+WIbbpfkugwRM+tERD8WqYVjC
FG38Q6Z+wfh1poAxw0M59QQ6vMNdfLqpwgc/KwmdPw7oyxhdkhviiEavERJHahW8Zch7niGI+GFJ
MWAgG0LCXVt4qm3HpEjJOa0WxfRbnmD0rWSoU26UCLBULKZf0C4VzwytvsV+F622o1YfoeF8OPsw
bwnXOVYOzQxcbmqiSdNjnL1oES09Fv71uWIZD+p/orzZ32jsrFT3w5QZHz6i3RwW7EJcEVbBN4Ko
tZME0BSfGpCKN368pEftmlOF2KueynsB3tHGprIfWv5Qe22MqLT+AqbcHNi6/x1SLBdHExQQv6AP
kTOWXClUcMhSJaSHuLMpS+3gEuvyeEs8V1EDvEauYRtArdfaDu/fMzUGJCBDXrTsi5BZ165qNuTT
Us+n2TGxrMmP7h680daXfVrEv+yHlXUfffE3QM1liqG3lzA1kneOG1pEbfryGFl5C7wonmL0Sm5i
C3Y+Pmnv4LYxgwFxmnnhZjgNjJOQnOBKT28zh8u10zkd2RzN340g2TxT+vW1152pDh2LWKHdEmu5
tBg/JQwK92c3XB6MUBFL1I5Zf+39H2TfbZlJS/GUeAMomlk6G2WjBI0/LBDs//2LWTuLoBTCbXU8
lNxxJxhsVOCE/abXe7OSu5Z72xLSJJJi2FxjxhaadtcmgvbaU6vRaLufM5T1kqnJfd7c2es31V4m
LqQAVx32Y/4dUZ4mmlAaMDUQyJntDIBBq3PGw3zTATweEL7kXeQVO3Y7XJp4AGcJBzTi1tXgScXp
FTdSV3wNwQSulec8HbsSBNRbEwZvoaq54/oeilE+5z4/wRpKUfjXnOzjqcHrh//4byyGjm6YljV3
jc5YvBr6RvbLAndoHmbtwFayud84TDv9X/4mcIJGSqJ3bXyqVBrKrPet1J4rpqwxvolnx818ed8F
ldTVMleUEfeiF8la3Z1x5udLNGSQzWwwC26t2EwciNQXFtNuVRMkKzzFDyksqaj2cWtC2U+gRNnh
1pq0wCg6zhVQsSP9AUG8/Bc8i+e4froBtE5mk5BGdFwXxzWcfyce3Wze6oGgpPlf3Rd9delNq+bH
W3JTQtQDKzJDwOIVsiCNL+Bv/o5V4Nq9kLnSPyJzmREIJg8sSHCGNKGkoOufrV6ExMFBxk2UVeNY
TG+eS+e0iha5IrMevh+STUVUvEtNBvF+2XmEOAAWr1q6cjOJ3MZJ5YwEffFkIf0tGMeWp5LsWqZY
oS6WXIaksB6wWcl0XacVp7LpKq3H3hFFxfkm9Fcp61L4JSjlCJ54Ne56O9lK+uvlbuJLg+fUZuRH
9X3kZja+z3+xaFgzsnJSdU1/TfQvLrFXXtkNQ7t+skShRBBmExhzF9Ns01bdB3khAl0kxpz7w3YH
2xLOXEdDktocu9a9jm874WJyMm4oEgfhpF3q5rG0kxTA5NV/oeGuJIBZZQm+Zxaa+qTd5GI5k4ie
fz1dHJU/YvJkb8pZatMXaq7g+4F1/RoCBDuA9Dqwx59XG2kJ8Pupg3Jtx6nCb4qNUJFWiM6SQnF0
z4pdUTLpFcL0hxOMC48BZDY3udw+XriHpym61SCtNOI1FPDY0b11Lc4DA/MTCF058gl4Lks7woL7
osAiKZVAHkiCuwdLnhNJDQ6gSc4FtvrVGzyIP74gAj1Bc9/8cezOnpNQ7oXO2RBL5YuSFSZ4hD0O
vfQrJA6x6I6Cn1i/JwL5dABPi0zeCp3eN0b4n9inkb3FnJ8I1+6MRjL0CxO1s5C9q3ygOikp0kwR
2kSwJcVgyJw0ThdVZvnIkf3pqS0eD9hQfWAMAmbSIPGyvzaAxwxPR6dy6aX/CvtdFz2lhAQKrFyp
BgYRUsM6Oi7G8FML5d4H80L5qBxoLZPv7r6RKOwL/0JiXuA7qVWJkiCQLZxAyXSGdMN+3QbKhXVr
top2haxYcIec30VFtxX+VX5cD3C98PyXX+54V8aNNezFxLclkHOIgf+rIPnurbjlTrAvzN3n76oJ
ehizv/U2H33QStN/USs1Qo8c305TKjRymxKf2dblzIJwUWHW/suEA9YPQ2qck6vmHyr2v/WMIi6S
IHcmwjp0gB3Eevv2JHT7sd3SRfWCrFq+Jqntvz4ojn3spgNlqeP/lKzCtm5cUS/F8/i+zQFkfzNa
sDx19wcYga1B+XGKPymGA8Q5Rp+4I34dehae/sH+B6w46heo5oVA7R7fF3nuLJLgM9hajH/r61me
gX7al3/Ttfzyfpwx7jWowwnjLn4YrWV/K5JUb835Mx2kE3UxICTMvHCBRouC1iaP8nkn3UAROMZw
4eNR0El0p5A2EKRJM6hsnpmmY78ExHoJFx+vnXjNreHJ5TS8QoDZh4np43qTVbcsgXW5PTWnqSnx
StYtYfsBKT8VaoRsdAWap2oAZEJS3tfobF75Fv1HaMP4gz/75xk040X8SYJiAxf2wLl8ddMtZDqf
twxtQv4cGfj1grr8bi1KIm00BSg+s9tuazPGb9RMwPli3t9rwn6v4NxXYpHCmlaNKCG9pQF48Awb
jHfzew3S1vDl4utSuANufL0RLa+eaeRajpBT1q8xrXR+0lEqK6g8rz8gkqRj8ShVs9btxUFjsSIK
le1SwlRunC2Yjkwf3KXoH6qSMNgUKbiF5eleufFrpFKoO7MHz19ZefsV2xSyC0ZdDIuThA/t/zXP
qcZlizbBzdQ+L7MQW7pkTPhDC7Afj8gYFLsEbCWUHVUI59LFYzNTNExlIQfRL893gxNW0SfGDfmE
fLsAgTXNRkYSRxF3oEKjUH1j++XHhA8I8edHZRhGR1sVUTyfyU5oPH5UdSyRMsvq3ocUZfGOkplD
YsbV9UUuj8M8kt4kscnT640ygG7Dw2yMlmKDEXbWXJoKhjm1U+pEavuIxrKsWOLZUPcn+yXdtFxp
DFuNtyWXpd3vdQ98yHE9OexQpA2AOZGhG3jNobhkTnQvfRZWylGxhF8DKjIBSkbEyWulGSxvaKoV
WQoUy/KNMxvJLQ0XxMg8YwM6LWcbGLMldYBxnQXlYvgNFeDdCEekLstf6R7WTbL9rYeMQtrYJUdv
g5Lgec2mnu3Q7zwvNsZu+eTbJ6pDOnpzy6P0wM/PZ80zfKU3fvqEUukJXHD6h3zPItPmJFuIyKro
mziFSWiAmIWDIIc2nQYOKXjlT07JsjhXc9FRaEJ0dKqTiTtmzznFWdhzvXxf/7baRKfMzD15iKds
aAaw9xfZwHz7X/IWb+MjuHdIAOKJZutbHQw6s1OCHr2KBaz0yhMXXtD6jQXIg/NNrmIU76HCvpJw
fT6WSJY6hHLKaizRoSgZ0NcSrvUCabHgP2kkQA16afclY6XGQ01ccvrvKphGMs45tc441buKKUG5
C79L/wuv1QSek4KxYY7tqkMtic0WzfZ6+DdLdyHb1ZfZE7eKXyGQqYm8ph671Q49JA6sRczQdFay
f7OVK5f1pr9wOebO3L0L7CAdCXHHmIU9gEH+koj1VWiRnPS7kq7wpxQ6x3JzFk2OyIHWAxYm9EhH
Ee4zeboRQ3AiHAHM/mOg2tNg2/4NXQoxnCP+PgyWT/r5o5G7TweSXJCRdQcXRG/2GmqJA3209Ikm
d18KLCFx6npXVsS/dEiQWG2A3t4dB/KGrXkzbdiZzI5dEpyZtZer2KPu5A5irhoHEzpXPsHxHf3s
x68HhjEt1B1mI8ainHHXjXIYoZ9nOZhuQsrLLjctg4FtIOlvTQud1Cc6AUIqDQfgZv79vQZFFFNx
oUj94FsnM2f7qHd2kMEcovFFe656FJ/JiAbRLhkY7ZkH+le2bngplezKfrzyAG1EQfuAM4pVPXoY
8aNJmGU5o8kYyldRXppc8owLrVwTUis0cqsanRfMJnAbvFNF3GSkxevzMGW4Q8k9w3hOFZlyE/K8
HOx01X57NQxumx9xf2baaO7T8le8Vvz/La4oHcv0qLutrejGH7/64nFlnL5AsuJ5pVPUsSPqTFDr
eoVwjKNLcPwF09QaLR9HUejd8rGJ3mYUyHYnepW6fkY7vPVnQoKFUnGWvEhvlPS+vJZmjmX08LLh
e0JN9kMGWvZGSzHxTprG7RTLyNxEbd5cH6Gje28bbv/wuj7Lyz6gP8YSJQSOIQYAmOCccXBBLKk4
du1SYMtzCFLIV+NOmGD6g4dcipk4lY55Y9BQTzxftEWcsA9IfSFICqBQKDlrS1LV3f0m2me279GL
AVFTdIp94MnhC61CajkKKpRElN5Cfcy/m4ElFTmk3XehIsfdujFkq/7jAmFg88KlesdmAG9MVH6G
Q3rYa47WfBIu7IBLS2a1pAX1uMvjMMQ47yVpn2yzlYhZJI4e8FxXGMo69zMvhMJOwuVkNekheYuX
7vUfvWlFv8hzY1ES1jPoc0ADtiourC8rxrUK9phUcFQjxvjeWV+9Cb8eLPJwm/z3Z3jmvRWr5egP
YnwuIthEDIj0VPjtVT305Fw39IJsOhso+mMGeN0sRirNfJEN0aEz5BxN/EHC38OY4JqlDfRCAajW
kgDmA4r/5XINDbL33QlYpjtuLOvPEMEgWgPPNm0vU6nsiHPU0I9HmxOa0GVaaovNX0RuUlgGJKUS
ckb0n0gEec70bzYgoTRG2t8nxpM3j15r+LVGuAxbn/tBw1ciCFmOErky+hzphSVGrUvqA/fRQW2g
TbLvk1/Gmyfv6woKovJUN0W/Yg7gJtfVh1jtpfuYKW/GQUksgSkLqujukEWKNFgcAxZm66MtXXnB
Oiq4YHFk2oTAXBQDrwTwh+r7FG6+ZGCb0bkL1osr4a3L9wMKoqBQJtf/W8CUqMZkG0VeFLku2WQp
Rv9+8Usktw6o1luO2bRCEiZEK0lOYnAlOV4mjv/gcH80o5FjMfpPTtQONMDXOLEeRiao8ZHiF5KL
FbYsypVK0RoV3ALrWRAxE8B01CViry3TfFz6p1s5PPk+5Uw16+UR9jNxF1RztO3qUWAPZ1+1PJsE
JmFFJc9g5UbnL8MSPWmU9KDDLN4zZX1EElZJSfWmaVag01ttPK34aMJv9VGpyxIyUOet5ir9Yucq
mhakvHjJEwvPui5pz38BzaBNPRgjxMx1/E+tbaNK9AmfLOclngwvc9GqZM05pw50ps2ViIeKQHfg
HGRM56Nr1zaIVd8TGgRx1c7kVEJi4DtZ98Zu0Adch62EVVns/CKkOqLvZLjcN3a9o7vYAoC7WWVC
eB0jJM4jZq140TZZ8VL82I2oWs2ra4G9vIZg8IltlbSBfy+RiUuQzvLwwpg1A2mQjWOatnYWdNpI
6AdfgsVquxGfdbRe1/GUBYDSgiXN9j0escVKCrw9nQnmwz2u9gYqw9GSXyBODK9Wm5KU4F64chMj
5v/x5Kg13+0HtWZa6mHoQo0/28eWnE/uqs6zrilviCGal+JWsDaGXKG6aTaqz/xQs9hYJPi2FIX5
QQYfkelf+v2eOMYAPmIkan6/RpIItQhTvnxnC/kfeBEGw4+yYe2lQsTVXRkmR/27WnQD9yZ5KoK9
NRG1chSO3EhwMGmqSUnzj+HDzSy/cmbosNvlroJsUvt6KbDVpc2V+0z6zdbTxlYejaC/xdl0Pji8
FCjx4YcqFcY190+kadnUOnp5eXZvV5SpTHMLX9fULm7BqVzoUx7aX1LafIrcYIBGDypOr5L+Fu1/
Q/6Vk1qgq8+QmAQVgBPRpMFAb3j/8P3UsLy+KeVX9t9uLN10d5LbLwmHPJxk9NX6lX4glsph5mVX
BlifX1SdM6qgKBSAi71gEta6YWj1MvRjyx+cKG3mh3FRXLiNRLb3NsXO/mGoaweE0SernPZ7vAjI
ltAjksJ/ry62/TbHWxs8nYUHZKxsaAoLZ7+PNH1bSjrgHtJY4MMZl8mHiHqKw/LqB/k0blAjXF0W
Jiw/RuZPFjNr2i84R0vu5mbNz2zdX0Rm3E0h5fMaixkfFygKkPG1wz3qJCBRBxuPBOtz7lsYF8to
adDWTvX/Vftg5E+en4gY76AQXgVcORL/LDjQ5NsQgd2VfWNCS3howtFYDmPL3Wz16hrjsy0jOfEi
6YkyHlN8niiBtjo0cg29yd4ETpCxc0U1qOOE+dSRq+BZ8r+3PCqOBpmAbJanfXLBbU5YtMFC9Yxg
WmoWt5tGB8Ou2lDw3XP5+z6Yb6Fx4uM9BEfGppaNfJN76o/aCiiJQNA4HexaIAsLWOWBZLkGBdtR
h7a23svg8RLvkdY1v5wUaicSWd3Kt/2YR3VqN+sf295iD2pwvPvHpuHVsfgZaUqQMHuX1vVSAraA
QOgd/iRUegs78l69BLV65OkFsg/b5Q8nc25PYRihq3gInLYtkt+n+1R80S1xkg6O5n4Gif51Z0Zk
h6IB/VcTbcAdTi+xG3hhyEyTycjSNPHpuCc62MrzP7GaZXjjkD5MvpNfsaHo69L8a6IOWvmc1nEj
sgTofR0MdHwTnYUVr1fjqWHE61munrn2NyeIur/o/JbVrJw7O3s8rJHSsoTSh0Bjrq5iRaSfi/e0
OkHMHUYp/a3FiSxOzKFzpqf3kU0gI8DeYHeKCiGACPvIBIat84/Rb2YQvKnHBo/JnFJyyJB7LEDI
wRSVKxpJwIIhnUX9SYSgCOUjT26ULCc2CMKiEZzzrU3k6yTzxd28l8GqhrKwOxlwm9Y+dYF1VtxP
ROkAOXAb7ZgGDUnyUouYFq8kuAuUyMdqhPv305+XpbptcXN7ePrr9kDP1TEb2CEZ9xaeb9EWPYbw
Kmjzz+AkV/Hmam95byw0kGtx0GQw8Dh6PpcqEqg8YQmUp+in5kmSxPOrqb2xBzxYThvrBimt8G/r
9DczzYP4IehJ52ZsK9c3UtlL/OCHA0g/iq59Q0GdZoBHy6TJ9yiRolDZfK4kUIZT6fAv6WYkzicH
mCcMtzKdgwQFd28lDrJGAoF+iG40dLu2ZlyVBu45cHLhrAm5Kmblyev95NG+JYk8V6n9sF4gtXnM
ct/AjxgJIgNBYNKfZ92Bw5rlCCryfYg996rnxzO+IZkGg8MhhCq8h4rD/AtalIgI7xwOi+DbXhbW
jm3kcXeEeqN9ymQNhdmEWGAR+pCZPkMXrCSO3rgxJ5maO5BRbc5H34oTBDvLpUk6m7snscK40C8y
bvR6F8t/wAfwFTK9erJpe1XpW9zd+ecUc899e4UnRYDIx90qRct5/PtM4hP2EwP+n6TeFrEUwlH5
6PTzW+09n9s4R0x47LIhxGcNtgQk7u2xaoJQ/5Wf0QNdow+odXANm7HGIHNPnzB3ceTh0r5eT9cz
wX6/SOFLcQ6Q/rB8QjnckXrdwdKeMLmPFa9VMQYvQM/04xs63Sp8bv0P2T+sdKwkjKOlxN45qwMv
Shl4al9lxEhzXnAHY8Nd2hlcnPptXd80E6N0C8PT7H3nlBbjSo5ZvMyRmJG1QObALWPVX5tgUs4+
HWEy+VMvSrzVyIrFsp40PloATiuOJN3UJhWwJGeV5dKtL+tJfp31YVdwIdFuzrG50sIG50r4T4do
1fTXpG2YvHQKx0wmaWxoLrxlmneUHoR1n9Ze7IQ/RNJHFnclsTnPCoAxjbxrMdOIjZgH4O80VR1o
eETlmhyzIOu3ndwueCMVjwaZn/MIQXIK5AH8N5LecQxGimaD6OBwWD6dSYPSODif6dODFyl0HP8D
UpQCV0ct7VzqTuM9DSma6i+xfiYsttj+pm/klhFTIutpUO8U6cwB5Kh0NwmyYA1K0xxzCz5jtibw
E3YGTLI1Kk6GZj6gJCOYkv97AYyNf833XcJTdwdGRNIAbhGd1y3FvycF7cm6ehboLnV8g1lZrq+c
JKkqyZV/9HbQyxKtsNcFauori6vcKs2JZCB4yD7G8lZmscM4jSAC5Pv+Zb8O2wJy0EMAy3+7rxET
+FeoeizxD8YNTemm7NUMmmJeG3VepEYh/wrIRvRr69Makjd1vUKFPLsvWCrkJv+nbHwMdjGDdreI
fGYZjDTQZz/SPJam24fznT3wL0gZOMSMwO31qhCCGFduG5Zc/rxQgUVI3GeotUZfbivd4n2YQASb
2to/iPRvPwnloLP2LYtvTCeMBM+cqQ5fVRG1P0M59GfQ+tnbLk0X7IWXva58o+qVCiTp76t8lMXQ
bg222f3uSr91kWUZF11S8y03Xm9pSTc3H/+LgyngXFD1L6zOGnmMs/5DVg5krt2+YctUZ3FG3ZgJ
j2KhIk1Sz8oVkza6yqXKwO3r48YuNRGRlwrY20SaZ3Qzr1dVU4aIgzUuu230mRnC2NFGkbCAHe8N
Nc7aAdqLkvVnIJk4reZK6MN6QchvmPkuhR0FpfERcjKQNbLa9q72xOZCJFw+cKVetDXlzzQsrsFG
5pJcfNbCLV0kCC10g8PgFj2S3sYcvhI+lq0lQvNOFb/l6LhDhRwFSXamwB0VrLp121/kksCjtkUK
YxWDEYPcLecX5N334LE6dYi3EzKx9il29LCcafIIq/aycevg4GCXWKLEVIo38W7G3m5P9zCay37t
7qAh9C+9aNpWwYEvNnNr9RmWjEELrvkD/cBbRj24G/cSYx8MRLF661PiXl7yWUVihtkbYyiLgznO
YTf2KT5WHrOeRdK+3KOc4zDW9xy1Cu6pXjAYaAjFYLGii97nNsd7RywQbYkjdNOq4ziCHE+mfSZS
3S1FTwYs/BONUKorIRD4iii7uccQZpjaI5Vv0zMf9pMOLBNx3QuhCAnO0NtgRnP78fhpqzxtbtfU
A38oOqJ3W52rzIeb5arJdR2oKmkeYzvDceoVRntnTUC3DXHuUnxjfVFzgQsGPv+P2/AvgH0L+a46
zIkP8HzKjuH2ZJ44ZOJdEzfXet/YEU9f3RAUXewyEAkW9R2i44/99ofQgiH/ml29Aorz+2AE527o
JVq6/ge8aZtUF2R+Pfgg5Ost0lOhILZmRx0OCrPMLx1EPGEIPBfclLMs6Y9kugnKZ+DM5s75XrQs
6b7pG5L+ewYnhIkTohIh6jCQJaNerDor0V40oEJWB5Gu082mJon8zU+DbeH9anvtAI+RmLZIgHIs
9Z66NuSuAQFEo+vUMyjkBLbmjcxA0uRGbMpHMkergGCVycAN1EdkwG/hCT0eh3vKNP9B7ePxQAMG
oSBPtZYAnTRHfONtR1VfJy2K6pEWjVd+L21A0hO6RRPDxUNxdoDR1Ne7wbjFHPEBwDGlCtHJ7aLC
ud5Z/FqjoIVrcHRXgjIP6M3YtlphOY7PfjG9wItALWnx4gnBhgiN0mAo82gcd8EUWbZi1WRJigKP
iVA2s+S6j+MvdJ+AvNlwVkcRNMjmy2EnBwzl3rKY4q/CHmaSrtkmKQINHep35UYLvb1aezlit5GQ
looNGuv0SG42CIEmqGuSXAdIFuRuSiqWAxHg1nuoJ6rUem6wvsNevwVOkFqRzBpOF2bAW84asEkp
KkDEBOUEqBesS5ucZ4sW6OekavV0Qh18/KGhJqttXfgF7YXZUlrLcxv+roXMPxvUbUSLZMvPYNqL
9IIkuW0S/idyFcctAxF/+519n46hSNtuZ6TxikRmvciTule+FrJ/GWHEKfsxkSAXyhm0J6Fu8ojQ
28yrulyRaFQynFK5XoAbNuTnrOKlAbqG1E8vlKiz3yXVIr9y6KqIYRSU7i7TL8/kMXiUo2kaTLPh
NdV/NwOXRMKs7sAKtDXD633N1c90Aog7LFlmbSHGx3yz8YCzg6BsxWKsU6uSn8ZjEydPFnhximtZ
/hh89clRN0BcgVDqefGxhJGKq7+A2OvKrGLN889rgZKy64NNz8m964zghQcwFndOwrFVvDKasWjg
+SeBVYkiONdax5NuUXcYfAVehUNx9svSNmLpgp5Y8K1T4jvBlbFD6+kaQl1pkQBXbFQopAiOP/xx
IRStanGkbxqeoT0swIiVMSh5IL3+bhVbmi93pVSv8rYq9Nz4wjdIUCJ+EFzAhSaTBqGM/gXttCFk
/b3pXRQIrnlWI+pBminVokU47853HLb2Iiuw8671jfJXd+PBPeBkD/fXutW8FEvl9DkhWjmr6sSx
WqZZuWN6Mg9CGRNNFQqmCDHIrUtimtyUGYv2h1LUBM2aO484g49bgaiZ4N6s723jdG0IURqCivaN
ytUBahrkkVvN8QSR/EFRyYwcdhMBHkEv9cHpBuKEi4ZEUX5AmVBWsC5nR9qAnBGE9fWz2Y4/FulG
1u5GPJbwdqd617qJjzpSNNbZoKkelKHwgdkHs3j4OCGsEOlvt3617gEM1nBfYEEWu9VEJl8/+OLk
qzl2BZZfl3/Wt3mQfe6XoSEZr49ESXNDxMLfoNdmIZ2ThJpwXLMTh/+B9zHNIMw0gqn1syB1lMZW
WHr6vjOq3H/UpGxsAyZ8sd/NPvmKOYcTHOkJT5HUSrJg+3A6pHbSdpsLnkKJ162yM1ngZKm5tFMY
+h8R9QVIAqSy88pQpS28hOpRUsPkbkzaPnliaMlvNRvWBciHC3O8OMPQw6t1q1gXLDjw+FT7OnRE
Fpv/40Prx97jmrI4Rp7D64MUTpDoXq3VFzH+UOnzABdwcci/glo/ETaV6BHgfuD9fai3z+wWabTi
IQq9V93RAe5p0GajlxvmmMgiSbB2hcBZUs6WBQWPxnkc1XnbRqfuAQ+ix9WSIpgAwzi5wJWGgorG
OgdIlhr7LTSS0rhUIo8p7BnlSKwQ6aUgMbGBj5ISw36/1nfQYlLYmbq7FCihamxiKusWQqWwemFt
yqrIFqLrlKGbyw8lZDIdUKOIWYEAHIfnhQYv/KmozBY616y2uHTjOtMPGpMobbK+Rmm+Dtc+CQIc
jawzcqZ9spGiZTqOJX3SsI4FdpCnIAQEIosCD8L9VpY/sYzoq+1ok9lGoLU+j2agG2ySREnvAgfJ
E//Q5UJgX3Up/CBHW02Qucj3cbzqwg0xOTMh1dhNVgVV6x1f8VdUjRJe/QD6Wz0ept54A5IQ91pf
sHhT0+FnOkTxCx1JLlqx9eEXlYoosF9K+l56JV3tHfBTgBaxY/m56xA0srW81svGFLwqay1JRp8m
a3v+U+HiH7wr1X8TIxx3C3yG3wDB2UJViWua/F6nc7RgHkK4Hl/p+BVwk3CQ76JOAKT8npxqug7k
e3jR7G23eeHFqY12ZefeS+kdOKCAeFXp2LFHf+8IxfSCiU+Xd9yvaX1g3k3ForFESMYvR3/IBlEL
Kwcycjs9nlsvxDY6c6uUoH0+3t9hoIv90qRXl4rbf78Cq19U0H8TA81WWuIQMIzf6Oz9qbh7S/EE
Yf9PqVsLi61MWDkP4FcUK/FiMMQlVCePPBXscoK9FTbUHI8ItqqrYKoMhvh/nvFRBHWEYbtdiUTh
IJAx5f9l6wn/nvPYiwXad5k+h92wKzER5oEwlZIwMC5tcBonKtrnsKMrbZqX3RVWluctRFnrH+AU
deErmd5nifYQm1ytVAXXQaPF2tZ8eo5VovFQFXbb6nrtXfXwiLlFmmhqPJHxRqLh/myOxWogdtrb
pRY5e++VWZNPZmd1QqtafHddq77ShZ8HVwEDc4n1jFw4kBgOkkb1gvMEiLsSKZv5Xs0EqsPpKb4c
Rg1vqiFV24IU93sfKp12qszR8v9ETHyMeU8guiV6JpXDYVB07kbaOnOukaSj+L5mYU3aEMKOPvnO
nb4eKlOodQ6g1xOz9NqVtnWlntree59VxcU3+QsriF8M3WUDDXDGArheeQrcad/LI6Q7ScgrYI9q
oIhuZ3Fu9K8LwUPQZUrj0ka4b7qyXgNvPJ6LugmcVaUJgfiXpc4Q9SsPj9uLViq3JqInvR69HHNk
COml6I6Vg+JW18nC5cRvRpcdvsISCi5yI5G5plTOQExsYk2nNYadFmTTJswvtk9vNkt6shsrLglY
GK+tsYkvSfPyz4l/XWk7+/3smnp3pUadxKt2NmdYXoVvfRNby4QKM5BHd0B44B6lRyz/T+fDXYaS
bTOXKIpsE4eRPznAeVXhf0VYVv+b90gVxgIBzanTdbolXXXFGKTEcKxu8fmSeT53AvUV1yfU5NRd
xOF7LeiR+FArrOH1Bx6qloRl4PJjU2SeJfXSutlwmC2WaZ9wl8dvrJ+Kb2rnM16kpvFJkemm0yKT
9LendXUKRSY4W9dvco2SmB4dhppio30tuaH3sWVxp8TQtPBljmUaGWUqOanmx3uTnn7Xm5pYclI7
psNjm8R3gQfKC1o03Wlzm8ydRs0dipvsHEMSA2/dlWaqRnYLF9K9KIHBLjs0OlR4vPZoiTuvaGgV
p+lbjd8JcAaaLzeWM7rJ7lRZvbbPB3KTJGic2gbAOxqY7hosDkHLpjTojeKO2FBK7uTwCWaPsl4a
KfHut5eliQFM/+yHC8TjNEec3n/zmUD/Pie38AP8kJb8JOvM7idB/+Csq1CMcE2yOoOUS4KMW3vx
p5hCljBI1VPAmBMv1c8CxdjldrTfyKS8CrLcVS1WGdPpLiGsKmkvX3tzRfymgxO5QotOX00fHzfA
k8bgVslwRS0TxNOKe90afjOm7VTobX2RdpeFyL+WWCpvy3T6Btxnkw1owSh7oa6mhQAsIQNfzF2E
M9IRXYhGZWixU4m3NJcg+ciMEGEGWLuy3c1S2A/r8UU6dWMHb7Obr+kfBO2Hm1rVi36azXPWU881
Hqh5Db7X/PqrbVUpY8JuI/2g38m0ckZhbKwp0dTMmWyL4yhEKsvV6XLjmd05FaABf+7Gjq84ODtD
TmpsrNaYxpMABQ0lA2+tMAycPAwoaIpQuj3eAvHNm00JgcZisa1NnSalQePyIPlQFPuMnLT7FJuv
3qljJT+qqdL8UPo7QI1rUDTQ++IXlZXqIvl/3GRqzf8B+NlW2Eu+P8LRnbR/k8smgCVcbMiWU9Ym
HbgChKZdnPi4bMb0C0u1fK1zgZrp0gImaqBAktrBSs8+nKwvp4Xw+df51jjD57D+jf1diPOGyOcX
2qEbGX0rOtvDeETq22IYKh4TBlZHoE75osXgwQ2cGHr4zR6vyXBIvKRZVwu0Hd1DrnaKC7BryuGT
Lll1dZwTVIAkrC0EYlP8hMcZQiRLFoKGHbjgZi2T08/WAAPV2pPZx5LdsJMdsPZAUYO13czxGET4
42dmwOQXpFAMOGGSZBrxBLn+OovvGTLX7E8lls3da1GTmibjz4xi0wdixkH9pSEV4ZADk2XT83+G
SjW2mO3VA1b1OZn8JdoEUsrFrZWecLAf8UsFZDa3f6UbH+tonJniwilYLvbYqvJ4rZA58AtbL7Gs
J+/ksrWaYTUSsiVlkv7tfRaz/RHLI1jc4birX6LNPwjxkWBM0DdRvViqKCfOnENSP2tivO984yP/
CyWjNOgk2HT0bTCoZ4qyYI9IpshbwavY7HLyPB5k9Q+RsXda1OmGcEQuw9lEZWMf8VUaVLQoo8yA
1rQk+rzPxdISRpr1s74E6KLIiuwk62DGbpXlYQR3/SlSFD9piYF5aKgocAQksZ+NfqAxmmjVupSY
ds1Npr3ASO8O43UuhTCb7/ZvX+0Z96KH6VhniBns1wSXHKSC6oeeGJXK+14VjGDusrIjtHJPXED2
P7Y7fEDHH8nH+bI0IPO1TdB0W/SGdBLovwIlVCDDxGxrPRvXMUfMAAC4tj5Fup0zc2VXfkQQLNGj
0Tp9vRk+DXikEZodop/MGmVnNeVYBROdrOe/Eq19CMO7kdY49xv3Djx87l6kw6JZLkj/IKF/bZM4
5MDGdXZQlXY59Ya1W2dLBzGVfIRxf86bGX5DChAIS7+XHodaJXe4lDH31IZ0Fg7GfO9UTDvhF/hT
hghtIGJ0ANs/5zucTrDS1hA0+khWNIQpDjjYnP51kkQ+laog4cvJuiPQ51OCfOcfLKD3fsivrIMg
76WYyCUOtDWJy+uJW1zetp8OVF70JNIX3HdhL12EO1BZbVYPNotX6zDpVsN86YBGSHNGYyQQ8Xzh
tz073LkrxJpYEksHHosjtaUqrjEnXIS5YvbuBTQx4vV09l5WQtljXsBuT0cuTTFN4UM3Ag0kPLhG
HTu4nh6TqOfuZif315BTnDnuIkQQ9aTacu9KHjPyh/Dcso5OxBZCjp/jM4NiAWEPsdnWiREjeNYV
k8rDIJSUjYblugQ6/QYJ87Mwt+7AmvgS5lT6ikRUXzHQcmm9bMwKt+EPwykciBg4b17ysnArSSLz
YNUMgFstwQMAYCDJIJiLaaWV6N0JZEosk9ysQOGljgpYwcdS2WMFZk9yPblMdESATYMa56Wnx2c8
S4W4LBwgrZXD7FMcTT1q+4XJ4rA1hAxznpwcgokrENda8JTEZtWLINorMmMpLf6O6l7bzUMqVmRk
LbVmRyt+F9CdFbb4yu6h3Ih6V3rV+smQ9qlzM84YkDiAsR/ZiaCN82WGlzLCwQdDniEXdmOzl2+h
hxEqfbxpUNNrDJvKz4J27p3Rxst5QvaVHGF/3S7ApaucMjYqJCgB7MZpnE7FZ/Osz4zPcwHI44QU
Ht0iil6SwV0jGZOGpoQeQrILOZgnMyDBJa+oqqzAWpC4VWsS3V5ihttIUn3Z47/c6mE/kdZ+W+Xq
1hrXIwJ/o2FM2+ODhaGaG3GolHsn8VqEHlie07qeUCpM7WszFTtC/+DJD0eZzgUalISTZDsGQgTz
9PWneXTm/wWAlm4SbYGgYnrZPY6J1iwnOyRvhpfGy/NiBiJMN4tv3YYPY3ttc54xRHrHHdq9BUvC
YCuri2xR9+y+BXJFdenCky08qAvXAy26D4v6cWbenyxfShv3z+MrZBr2S7i5TB9pKwGd13GDJQlY
+kx2jBZV5SK9WOT1xczUqHj2Y82IXymW0yNZkdxXMXcbUQmJpV6yNpOPU2hTyEXfiQDg7x9mymdf
XtB+063PJsxyyR8W5zPfzzrtYCXlE+QwJ+SnmdfKxHnH4r2FfvzOfqgecXq35u8l+2jehShcOLM1
5zS7I2sbo1AQ4VRZkzgLrrZsqiq1s/7MNZoeD3RqFmtVll/DIWEfFsxjgIu+WiwJjPpb/o26XXYt
A4lGxW+ZGxb690QmQ8k9xWiqQ87Sjkn2nnyyyUSXlRMA5u395DVpXixZwVUgiX9RhzQrTnoPTuF6
jZQmVb9ch3Xj7B2T2zNKMcf3tLwG6yMwFtA+KSUcaYyMtr7CfeSNqfGfeatimGxuHy6PV4tVTTXs
wFr+ku/T0YvLTsyVEOmyaTfN1iQKS9GuX0NSSIWkL4r8EV47OJqo+3oe4Xg7st+9SwVUME9l++iN
maywzeITMA5elbOynEsabiI9ry5Cb1DJ05jSgwlHgzqK7+v0Dt0RVX2LqRUm+x+8Ph8v26WI9CBS
4oWNeI+EW8ZfCyNKnN/5HToiqjLkPRiyATDrplE1AHxCc3eIkcsdDJBovBNWFjAaoWIexRd62/2Z
XSHAA5oGJqHXAOpPZdG/bhBUXIxkZDz+VMxOqK7/3dGUlsTebmKXUD6RPycz8i9QpNFFF3xwPMh2
0MoWPlxpxORMSMK60V/40jv2abtn4cAZF9ypvIWh0bnKVVG+nUniSUGdJywX5/Q+rZGIF5pLVPup
5WquzlQwScBHFTVaSwrQ14ziH/B3F6DSxnseIicFkFrjdQFUbeNw6K9pSI4cgg1YJlAnvUODxf3u
8oJT8rnOUS3aTE2VNwIE2xcRjEjm0DG2tUoln/WC1FiiCZIvzEuJUqZaFErXNPPPSyyZitGn2zW6
6LpUade1aZzeDTw+VbGSIvlXLwFI58yQKHUwDtgdl5t4QXoFeIDCd5zs6/EAUnFx7vgKWwR/AB4f
ix9xPsXGxYpHF44SI/WgTVys4mP7rirkbOcRyqe04TiLJirhwfgcomRzcdkCQka0FkaMy/iOhRIW
aEkzszne/9tdWinfIUNbqEbPbjoTKTtGUJSgnuUuUEIcAu3ZwDhLS1Jru4Tomy/ieE8jgPXTfaov
EeS+gH8EIBpR6OHfCK2TqWrfNrpTKtWZWlPPsyuj1+1qhdpNJ54hRIiW6qBoCZwP5oBIGFEin80K
w88XrZXKjS8Eqi+MWfVMmzYZ7LgpReJholj0X6dKMx78BJcdCGMJDtYd4wrAjsfqkR//43CawmNc
skZLP+GnCi0OLMCoFhLKDhL0WJ6+Lsa96r8iLIGQQTpWHylXkfcTPQT5KJHuX1uydFLOcJjJwp/i
Pxo83Wlanpyx0FEPrZO56b4Nxu2GnPuuDvSmTbXXIbVUEKESx/QsvEjHVAJqxQCyA0ifozDC72me
QF/8uQgGxNq9U9at+KAbPfPQW6svvxr54ELlcNN7R8X2as0NiM8tSR8Ox1MIEyymxtibz4Yc1iHf
2BwUdYvP8j518lzKODqOIoAdFm4tq/2PpGFT/lLesKGz/p8osOCXOdw6THmYtIi7/Dl8A/DClqtz
X2Jf7ZNihdgGdGw0r3Qqxx6X66GtvzhyP1qUVPPM8oiTMpwn/vgSNP2XxInlRmAv5p5vqzCwQuwy
6P5scQktdnrkzEk8YIoszZwQWAkMYD2DbUqpudDkZQUACC6jMTB2BtCQIdd+ab6eFaxpOBABs+JE
Xy79UOcW8aoZIVVaxzQ+1nAXWJUAq7P3dte5Suk4PIdjhQWb3Y18pmmyeD0fL72GhOuCdXeVLbRT
bnfiJjur3HdoeztfUs6UHH4vANDsfkOV1gNxiBamx2I4y+1VrQOAnWh9KOmQ+jLfbUq20UhEJu3l
9WAFh3Sa2OahS2WztiJFmXm/Lz5gws8ZL0DlJBXtcVGVnUahPbTDpz5yZurzjMyc7FPacwiSLq6y
cTeGqWNWi/KOV9D/f+/Khv71NZ6jkwv8vQzpiKF/BJoqy1CZOc3tPtroOG+8ggAPwr2KvoFvq1M0
jU+6uZ7te8o2r/QsgwAdkt3P8UMr1adbxOVyYZXDtacrbDMY2OcXqgG8CiTmahXDilbe+svqg3jY
mNMHEFW56ODufBEJyYUiJs/bKuN871596qTg8NeG+DgPRxWkOwPZPqGUqLmpRPpECCY8ZJVSm3cJ
rh70bR1dPeWgTrdzsF1JEE30zvQAR2EEzqbJp3PvkEs+UcdPfEukhfs4nECPqYBd6ttiHTtvXNI/
1u/o2S1y7iSWzyPf2JMEkYYt0DcGRDtg9PdtSKj1Mx2toxH7adezCrE9saBApE+jdqgY1AaUll7m
2EzSqvolf3oqjVVgWRy5Suxp2yb1X85mLNbD0LmjwUG/2RzqUK/2TuPYDkdW6HbYGBIE439JwWsn
aW9Pmk0KOODUTLOxHsvXa47oIFKD6hbF2zAXCnqJZA9Zzz59U7iY272Fj3XxxcHI3fmO7vq7N77d
7jMWl6YGRnL1ClCt9kjveWOE1uh16VfQZ1H4Lci0H0mHnzD3UBLKaNw7henRVAaWA10/9S0QKzR1
VhIv9RCATwTprqvRYU7X1M9qOrsiWJYDZ0b9rrNVTfAisnXuwyOJqAyRWK16kCaM24vRyzm7rufY
zvi+Gag2i7MPLVLhJl8oZjdAZ0QkNGoO00rRZhjHwCDXMDYW1Z1I7wlEM9I72ch9qIeaq4fBw5KA
oXt9kJVWwNsbUS8hB6dQgP9xUp7kT2w2iMdbZWHyELGl6/p9+388lGNNrzlOTAIWhAf3SLHAFJl/
F93m4VGNf1a7hHNEnOztQBiG8gAchEyDMYMIdf/93AWBAKadHo54Zwvb9ic+DXwwcYwlRDcHqZFi
ckDof+BQU6EBU0MA/2ddenFY/hseyCKhhLLs12iGYenhOLDU5c2rabMbEJDQsBZ1e9WsL1urDrP0
IEzrZB/nN7n2Qf8a2lCYwGKOIObKwAnW0e9kdplr+jzkuBgFPZN77F6o6R8YXKKU7BwmEBCSUSSM
bk5yU7lT05i6eeoJng4GY8C3Ask25EZJKDPvIGJdHPPGNmhp0IpdwMYgL+idsVNScsPJ4VcR1JdZ
1H/v6r+STkF84DzXdEuABL5url90vodUX7GtR1ovuJJB5r/XxvRX82lvEWNxgfQvtXpvQ2SRlMv7
OgFZm2UCaBOX9jXEYsCg5zea4K08MMltx1Vmd1bRS6UC9My58fGjuvb9AZFr4AoyB4DGSdNU1G01
LBJ39C2KMpFSRTbUltGyJU/RHvfwArpNraMcFyJkTT7V0tIiVFERplIJ0/kxiDvVVGyn+MNnSFqZ
kW8vBMl42/7s5qPzFiibuJUpfJmj4cpDM8CunPvP9gek1MhPBVmemmKDnCu4f1Q/JNjTeX/uI2B0
ltXPBp65NDmIjyMYxDYZZ5/kuuKefItwNSa7OscFuR67roAEepiZrUoecKwPF8TjiVEzhXarHdsa
haISKrDMQOSpbhuekR44FKjnzNhL04TFYdLs+Cs9fsTnZcHa3KKxIIxxF0D3aEDSqTzP8buYVeAR
WwsbvGW64tmwV7v+q1Lu2u3GNcvwSD6GaStHcfgKLttrNaE6NyTRs+VJef0TpWuYuNppTZLazJUc
I3F57Zcmtuj4dVJj2r8i7gEaXXMR13cZ8puiBYTVptr6EdNoxkTNfNQk8xcK8EP2XgAdjAYVhnFZ
vWLfFC5K8YAbdBxX8voBfgwQQjAGpCPbgGJ7GFJfXShLITAwmIU2se7qK50CP8gHe/S8u+3x5wnf
g6wzN1rWQZ+Q3e4HxYQ/mR0W7jowXRP925iSIwYvtTWthirStSRjyymriXHmn3bs0LAz4UAQb+/q
JWB2OFP9XFU1DdwYE3Zz7TDES3GhMAeWW+vbECgmajnyWGjlZdHZny4zdIeMMir13dpepBUwJOQr
kAvgfU4aQgpxXJXl4l7i+e8NpfViSmBJ5SbWDDzCmUINy1fINAGsklFLo4q5rDqyQYddFLUFYtRc
Si+NWn7hMPYsQ53lf3O3YDeWLlE7gvGPNMBN77ITQL3rwloPJO5ZYsawapHr/ZNHBif/wrMBw/1n
rN/qtOwvfPLWXlRkIo0iItMjtC68FzWwDnFnHm/tmnatZJ/8wPrmuwoR/HCX+PRQYKSqyqTlZ0N6
mqxsAAADBokWPy5Hr2n2FIi1eltWun++SdCxJJI7BXS8kk7aBQyFKuF+xfOMBNVWt7rvRYjFoeng
cj+/ro60FHYS5UtbUhLPJMwMEUj+7vnywDK97kYbyvwiR2fkX7SVExLaNVj2/PGB0074ycSFfILc
U8Zzen6axmuD6lhtQxSFCthxUDwTUEBaLoyWZRAV9f8fg8jPnIxINraPqv9eI59ydc56BdkalBfX
Bv8bhFclS1GatRaBgNwHJxcxRRo1uc5hKalHutLBmPBz5dkG+mjkRxW3ZHQpAi6FnJcPzqB9fsos
l4C665qADAePF/9GlGfKkKbChbWs51v8U2JmG2I2Cdj/BZbthExyA6mKWn2aEh9r9qXWX4xVX97O
NqeHyt3C7ktCpluaiMjhIHFPYsme4rbT9H3sl3QyG2Nml2PBzdZDe9pdDrISrIc35D7NuyAfmb7M
Rpoi3egmBswEukG62PcFbLWShsM0/JE+beWyHBzFeNj/H70sSMPRxsUwlr8VxLAp0bWV/3WtRVYN
IfCe9z6mkxp1BKxWqGCg7nrcM2npZqYHg89KYqeyy/45h3of+7UAKeN+TIDNGwFlg3cW11cS66p5
UcUEOg5mMZzWiU0PhlyE/6w6q7JkABOZ5fW5xsw1udba5FJMoCVLW1dstm0E7lINfqd7I7XF+eF7
4HJM5rjuYwljvzacW+evylSj4yulb8qNLlOV5+S44xMKbFrK21viKRcpI1LhxGcz7cwJy40WhdI4
qytedj5GSpbsXGMe1rM7TiCj1qM7SKa5Le0A4ST6pOrjA49ufvETC69N7MjJZKd+maDFb+HS1Rf+
uFGWoI+nylxw04tdqKoEqv7HjNPae65XtDNXb/3uQPdsbBz9+JQlaW+oREnTVzZw1Pup4FpFCB1K
fuI3xLe0dPkKDQIfmzMoLfwVwoFIVflZ6JgLXJmFz4gwsxxhwK+G1M7rI1FeWzYmt89CX3ninFX1
z0qSVAONFuyklrXCAaO82RkVuqXfpwfTQAMTvwJhGAqUJc3kCIzRgof1YNVWTMp7kA7J/bKUmAE+
jlWXQCP54lCllWC4li+Ow+TAgPsWPLTGPQuju/G97cjp3kHJ0j2XxufRYF+nO0QdxP+o/lbAXf2j
Hh1gwfUIPk9sTzTqeUdoiN0BGAzCpuJ4OsgK/RSW9QrZ+aUBZUzhwCHli3EBjZQuX7f3RfYG8IgS
0nHrf90NO1cms9/i1FaVwEEhgtsIZiLYHVoTxHqYLe0cwt1+0K13ufDdKYSSTpSHoiHVwuybilrk
jb6oD1KAy9SwA3lD1hWvCFONCm1jt8DAFSDI6gJlsqjspvP6oQAyLfVILynVOgAnMghQW7uVc1VI
07hBM5q0ZwqRDZuCuKVH13HLJm6KVEnyW5/GbBvVOdmVzX3OWmLFM0tJ52drwdQvX6b5Fg227GD7
LDFobzkaGWVaGAUGZyJBAomG4FHyTBbsfjk5vmY4nc3rQK9ZZqyJ3fd7Aier3Z4BUI7VLIv1PgO8
l8/Ew+6OSVJIjdo9j6z0QxHd49Q61O6XNPdqEn7cLX3OcQm5BZxXWiOuqLgAeV7zDyStP0Jbcpap
Ye5pAbOsPFtb9grPzg55QcpNs0oS+q662zTpCKVpb4ihsnsOLTqSbfWldQyaux3AEYBH7qdfylhr
1TZynQivvTG89i3Z4mLIVAVVxtzJHp8C98T1zmL5dIttkQw8N95pHFRmXs+BWgiqgv/wxmhAJX4a
lKpcd6Ykg14EmZV0c22yEI86/46Mr5X119d9fjNQNg3sN74WBCXkSLeoOK/ydKeuyl/zg6B7gTDm
RFwB7XIJUtl6Qn626bGx2R6NnVEQZVqrdd11DQc3n/ohpKEAMSW/tZLqMx77aZYImM/q6yd9P7yT
0dtQRvBxa7H4dQa/XaGj7Lo7m0P6FElMmw1OwaTEZx8g/jHv+b1gej1lSW91C6d1jBjLvzQoxFgk
jyAzfdf+K1FUd9NIKgU5R9mk+uAo7p0F12wVvnFv81isYX/QKyfQ2dUJRHulMB/GIKgBGx325pZr
eT9ag16s6lxCXeVZu6W4VrRgbaVEEKkGoxmMW+Qz2AiXYk6XGDOVjUh+87l6tskmVJdaKNCbb/5K
u4l7gUfCmtYqlKOUzmMyBY90uI96plk8Gy7VLUFqlS4Y5IFe/+kjjza1k4POb266OOFrXlWHz+aY
Rh78R+pgqWR/rmecz/MOXHViwvF2umC5g2qOfovs53baWlHFNYA2J/w4LUjlECcbroaif5k0fYvj
AV1M+ZyTdD9355PzmUopXTrx9UQ2QJf9AJKOTTkJRcqb72cBf29EUgTOQLGM9UUCKm1sgExIeqGg
1ALRW66EP1LYYtUwGBsrQVrqm1ZpojWqHm/dRlF1x6L4L3X7dcvD3Jq5l1ITrgHl0zkjQZeFVzhZ
9KtwJ/TWAMPkhAr+OhgYV896kKFIgLndd1UhK5ZgHzGIT2sffc6iQ4uLVAZgl1jTmoRPQ67XfCqg
IJnpuexwIgabEkyL1aK2zHWOAb9lmb83a+wmLjMSpSjz9AIPtE3x9i+9HQ3G/5B6na00lc4UWu7K
ULuxVpQARq87CIMuXI2swSSyfQig7Y4yTJlbIW18PSSZlsBPujwL0LBxYvtGug+5edfj7xzZ5H7F
cwSrvtMU20Fz/n+jRTzwXwhdhYNDGJUUjjPM0Wj7eVPzu57pzB84FRzpk757KkdnjsGOJWDPnb/7
hFrL+YsWn6LAsi9jaFeYXdBHXzgsNkoY14jkPBDk7R4XSMOZjgw23lDU2Gu9XPl9mnGmRG76KCuH
VLF887y/1v/Yym3gAw10Y44xqnY9VuWkKl9UkBtzUp2l2btQQ7IXTy3Q3NaUwNod0HYDPK37YOcJ
ZZzTBn3gv3ZY3dea4sbkw3rstJ60BGHk2s9or+F6/cSOnkAjUwDsO4yiPsTZZfanFVMD/rKDViFA
lVo0REeg/4vJTIc915eH8qK+y45lTxrVCfj/S5O4JUvs0fXVTIVA9KFZ51M8YypiH6yA7cBR7MVv
dyHGro/2hr7j1qZuRFgOMDvhx9XyI9Fy2GDIBHLqtlRoBrb6mv5sxUPpVzbUxrJ9Ks1/mQVAv9uX
01mZlbOzXkUz/F0w40dZEX2a7soFCX4PMt+3lcMOky1o/JOH7jIJJhCGd/kDi2VSH/EMb+enlewT
zzshKecJhOGt3QlSEzCpbMxGqTwYzcTOSppQ6VCR9jdZM+rQmjsUxQIwhw/w+7dU+7m8WS938n6N
FZTvTBhOL5mB0BAb0nWgFtKzp8sp06IWSmpng4bAxSC3/7nV3v68swvUBt1ZCh9EkuL5D4brLIRQ
CotxusMKaJdii+DpTTZpc1N2IiOXDvV6aGyFXmnO6kAW2qC2SwhlWS1vJ7nBstfcWTFUT4AK8MsG
GXa7EOWPNTcGaiBfwWZVgi3h39fIEHupDdMnrGB3hBNyqhk9E+QqAvqwEFgZxRv5UP88Px7ACxK2
sVtkdkzspNf5WTlzaPEEH0XINW/MTt+EQdOKcwxdf42yP0JUUyhZfaXMBpZl9i+LTHwYRcuURAO+
MX5LBipBTevrkreI2/zNXScn+Sy47xgdQ0WYD2WI/BEE903/fjf178/2+iaEnAdWWN4gxzFfN7/K
kbq4HSA9Q07a5ZacEzQjt9pS6dMxYAJkBfsFZ61mAaoaK/fPzoikzltNPACHQJ8VzpFyO3ylyMkn
YeTwI+kWyvrDsLXmSY4bNqxmYJWoYjYqjb1e3IXYKuieIDIjo+EGe5xfKacLvPuvV60oST1376Zy
JIks9HSMvdfhn6+zYNcd0K7f4qTzH9Hf/Z1bERJD5AfqZx1Cp9qaQudDnuHTEv+mYo/YYcRGirL0
VhTAaetbNTVUHKnW87Jpn/IMd2EXoAsIlvNrCOV27R9KyO8cYW0sJdSV11osL5EXNBOUATs4VKQY
PPjhgbwtfGuNwvVIEFWiNBfjz9HAvauSwBagztqECKXEF3Qh255YDt3kepbfhzst6kXqLKvYh0Kj
0ldYAJliOtSYyg2metBwmFiI6cfgyUBMoXOb1LM2XTlZFSv6/vb4T41FSETgGN4lGdaTeiebxMTn
LIMkeGGVC0NsIt8KmVqoNWc57i1aQ6XG57MNN1W0iciwwV8oEopU9JW+lse/Q90KgI5Dg+ym3WOU
7p+JzjVPeOYGhcm192I6Wea7ZQVfCqZ1B53xmCLhcraRC+/4LqgB/sTJkgT3i6PQwspG20+u5ncS
u6L6zBBvvFr8iyEduoauXXZObL8+hyOSgelN7LOoLTj9cX5DJTvgbW9EAjUCFI6drsyWW4AW/k5d
6bCKTpoJFtS6YQHV+ny9zGuyOIwgT1dc3TkJIWb4XRMRf0ncuUa6aOO6tPnsxzh8QyieUNcQaNXG
GEj7W3Aqmx1xI6JRCycq6MeUmnFeeyDPaDTn5t4Pnj4S2jd3jsNRRWakX4AtpCtjIMP8Wpru7gZn
U45FRMoK6v4iB9fE4ST2lgTlW+/zXFiJ9z3Fyh3Qx9H7OdZmjAPQfQK0Pu5pKf+/PXQ634aGVJeZ
rof34fPLEkWqMoZMt6N/Y2uYbHDc14toMS5yIPhKFJVRdJrKGLvj7QX0Ds7OKsLtLB+axyBi9xX+
CQx4whF4k8vcWKbeKCs3aKhJ3nAS6UA5t9jHfhaa/XEdKvDBCeY7tHoaNLU4Qx2gQrMESzdZW6kL
ikZWLfFgpsBFlJ/x6KGNvW6662OA56wA08vBVso5KnZyzJNabrHE/jaFuxrvqix7EtV0v/imo/Zy
6Hi8wxtWIQaMOcP8/jHd+phFzEXbuqnvkjpDL5iwY65okiG/6CPc6ldQMChf7EG3woKNuHsSCxnZ
f4CGRVafgL5wE1sYtL5CkOTKGqR3Sb8NzygwPmt/z7c7q6nEsF1IP4Yf3nezW+Duga3mvBlHE6fZ
yuEEJgg0WQ6rixWiVd+p4I4zXFprl1aPdbrSsfcEuQc2RahKZIHIFxGk9oZvlIMXwFYuLlqsCW9Q
YTdTGhwLceasFxK0P+flavU2M0dgRQ9VNxv7SJismBwjL79Z/VAX5UnR+RfQU2NjcfVyzqPYbznq
KC1TyaDXGFXZD99x0b7fdimNiGpf+sipojCfmZIPJjoXahDr5ZDa6X9kNatIxam/7tcpnT/GKa+6
VNCkz4NnMM1yXzLJ4G5Cue7dGl2u7tfnpPxI8gbimvvAStqkNz9pjezkEnPFTXv8rxpmRGV3SftX
MaJse7vpPZFgChwQyJggzkWeKxWejdTD7ag+XcAOa3gjcEy6tH0Fp9sCG7AQit5I+ioHmISd0e0z
McRzd1BjO8Wp9iVnMigmIAAKPsBLY4SwmFJp5u3dWQJ802uAfT9XEDgm7vGf45W9ncWZFgECKVvS
OWRFAUD6st0mS2n507roGLWtiSzJZNP35VAqMaI+MHR0RNyhgIFgd0ptd0bZJfwcTL6gzH/2go91
wsr03x3Wv5n9WKb5iR5l6Tv9TXVpdLBDUbgcieR3W5vEH9xmic8SbWKoa53iUVKAaNW2+Gr3lhB+
ibPQH14X0g6dwrZ9J/EJ3nbPZRZEFDua5lUUHdtKWonnri4LMSO3/t46GDG3TT79VUk+YZsD9BfC
VDhqfP7d2eHKmtcey9xJ79jTddAG+T+savcFbdiL5xu55SHNUUqhdW+3U+gIoPYvPxI4PkbMMNBH
XAvJfT/OGvgXGRNiko/ufVViO0BOn1ot+KV32UvcBmu8teg9em5o4dbVnmTy4LdjOQ1ARYeGMRs1
8J7Obd5T6+8qxZEA+epNKo1Daq820CuUkAoOOtxWlCpDeoQZpDGdlSK6Fk9NE9dyPF1aqiH2icOJ
M7MqcweYOekpjqydJXY5Zj9siXHpdP50QR8g4s6skmPUjx18V4tlbP4cs9TsTLCf/S9ivfK1UVnv
b3tTDWNtvtvdZcLuaIB1Kl4Pvvd2bzSA9xVL0Y2Bu8g/1qJoR/xQCB9KZ9kQHBTwZl7J4LWoT54v
BsKoVDyp12h4/L1vstqdOxpO3sffPFN8C89Q9p7qG3jO4e1JCcxD7lpIW3zHAvhDO6ZLFuPLYoEf
NF0AH2EoYQcl1UY9hOTLB7XuZ8FLCItoOBZj47Rhies0wbbRbTuhv57l5AdSgtTfOZr8kkRDul+8
fshImjkJT0QqIGOb8Pht8YrAv+01IOO1C5J91NLc+BUTd1R+NMDFybxOXa+/9USElrC3lHJ/tSOD
GQUVCy2BjS70EFKOLmYlCYMOKgeWjSFonZ/sgn8qGWLCzik7q49jBYAktFHtRxoHeeXj0+ylEcZ4
nXq7QnsAIdbLk3a62b4whPgKXtuLyRlCF56egSoRKED4Zgl/S4tM9865sk7+RSHfF4RpIfXhh3c0
Yq3MyqC+Eb+Nw80iafFyxrGL+iMRPnCg72QBgUZGlour1Zcw+X6JugUPfuIuymFys4hD/IfGrdlB
2XcnkPh9qTja1RTbntM1myoYy1G9Evf9ZIaDTI17QglLXV4Sbg9Q+658VmW7Zh8NOG8pJCBqJZ/P
vpYCN6zqjTICucFdqF2oJiP8aAf5yA5B5yFjttBr1cUx2XhjuKPgVVbCVCqWhwDsfhIKbUS2E0t/
7h1GPi/QrJ+4J1zKHoNM2EPTlkc+SaNtdQeOZstgoftZ6gUiXKPbDW9tn0WO9phnU4T/Qc4myQPK
vMhAaRtgBVEvLa9ApTKUqDErLV1wMZqikUZO+o9mHEmmsL8+0g3YnCoBagZeDAHJM6JCQVh6iT24
5anftMhyLX8twG1sw/Obj3dW6IGx2JJp8rGsFebqHCdqzw/e4PPLr5nsWp1Jm1Isgb1+sCgOT5i3
0U0ZnbkgU8pAdthwIfJbWDG5rc2r681dJJMvwpsp/rHQwSBzilacVx0J5SDKdQ6DWVdDZvI05yud
iKmtawNRCSU3oZke4DEE/ZyNiw6hFwZfO8gCbOR1ACsvATe38PYMCSuLKPRNxlPPadE/EcWX0pSf
iY5UkBj2KNkhWZKNxO1QwzPTuHfwyQphjmbiCSOhiGKB/Q1d4zoMMF9O59s2oJfqTcCwV5WgtDKh
CHuKVA4phkO7KL7YwbEzYlaT1l0jSp6ifWojKAMzpzmOUz+Hg+AEAzymEcW16yf6LE1AJiTI3Q49
9IZ/OgKEn7qMdyqBQQcbBg6HhhYIRwC1i7kxa/RbNyMhv9a9B4yOvjOUvHan1evzbG3lgWOQW+rq
J74VQJHvcT/wieuUt7FBIZ8C1hfuykYEHZEpvj2sjRb1Btthw/7R9D9UvfwPTlZnV8mbl0bvHOeq
poXl1PUCfvdq7rQ4mjCMQNpMHfXOzpl0YxBxeT2vCx5NgZ4WwCfySYM+JADxHM2cY6mS45GHyjTk
kHrXZopt3eqnjGHU5lxAOjsifGnFykYbRZ8MeFtLrB2yYiCq4PNoEU8kHUfxun0ySsU5uQrbP0Gc
yBPqIAnLnfjHzKV+LBvwVxDtgOO3Uc8E8Z+S833AjXPPVQ+1yxVSII5y5gEhSZWoo79FmLh8lDy7
AjeVfWE6FdhJd+FEM0aEFHveLCjBkErJIDW9Ofc0/WqFJQXay68xtoc6FS/KOEAimP4T00l/I+jw
dbpCBeW31I49Sph5Ot1RAyYvRxa6kLTFKmQxws98srG5VQs0ULWy33+ibFgoQqMSMWVcUpi6yje9
XPPAC3GdAC9THaO0Hf8U4Sj0bKHkGHgU301m1yu/vjJhZpxsfQUZucV06AfQ08+fv6w7yWZiUb3k
gqU1DrO5+lSE8NmclKoYIKbYW6g1cD4oPFEHjeaeMs31FyoVwUPTVyc/h8a2R8rE7bYOnpCHsA5A
TXTXIj2E73g+jRukeQIroHVr8yRCjdpyRDYHF1Nk1Ietc9hNQgdaoZHrGNKm92YmE77oVtRk3rH6
MA8c4g8RFasPaB9xLB1CCezfnLEJ71LTFumUFGbI8RrHpuvYAfMt8QwjtpELUME8uPiEyvK1NW78
Wa4OawgHwcqZjV5Ot6gfu8qdV3oUel59fD3AXPH4aQZkUKOYTsGjJ3Ln4QLPs8IncAr9yaJ0g1Uc
cIwFESnFpOUs87djZylICNPSs44jspbryXgT6EzErGg7DyuIVihPpY8OKbOV6BrULD/4jAzmB/xY
A99n7JnpioxoQgOWf9PCYJmINO9EkvKflfrldLpucTS31e4ehXDB+ejUptTxQljUv7CnK8fN5+l6
mq4qeBmWT0qC+1OPMamL1BpFTl5e5+CFqaBOE4342FrKYOjBIICcCjVa/6xLu9sXyAGfY2UDGqUA
ADoXu4Vr9PbAP23TOAov06HfkSOUzLbq9F/77PY64csBPdJbJwLebgAwNpeq779WjqoUThymjBtE
DLal2JN+vIvER07+3jNxzoNQ6AKARgX0n9eTx+uEtwGYr5xpUqlslajEVng425rPFEJ7y89lF9O5
unAsnITFlfbTlitJdMpOlyK6+Y/xyd0mIpqZRkAcBvVOvvwybdVXMpPzPpTaxZ7SM3bRKQbU71Wg
BmRJEuWWrX9MZCz8Y0L5QfPouBO/HvEfWsECy+2xzDK3GyXP2oPg//MIidlAIi/y7Lf3YHOK6Lvl
DSZMccbN0jFVAfcmCptlcdXx/0dInVw722LDEcztBSeDpeFur+/BY/Z09do6zW+FGUJD61Pnqjbz
kMdzYTKP6dJiiKMzkBfRP3XZdGHBkscOKYHQtp2iq29xb0Y5ePqiXhbTaOucm2cbN0sOmkAaCk7t
VY4wR85R31NgDPO1ijKwQ0S3+a/bUoERjpBFIqIuM98tvy9iUfJu+kMWaxl9eF/1CIANK0oRr6S7
4u4l7iHhlKEYQJuIhszP+8FJx30/QJDMyXT8Ov+1STK4aTuD0xHRADdNWhEVDyn5I9ZGYbwOKctv
UtiawOK1Ulfx5LY+0+hRGgWKBqu6IUzTPImJG5dzrt2WhXprYzWLhAlo0LMH4AUMPDRP8eD0/rO9
I4tZcS3a3wF64DDZKgvq8e8+oMtF4DXZlGz8q1A3kiK/Xiy8v3vQGeluZERniA6U3WQ658ijlirY
HfYN5qGOw6TRVInniX4YT+SqlMDNA2LkFmIHN/JgdDe9idVn/WpwuKfZIBjRyO39oPtUEyFGWXEn
L7b7awKXYqa7GodlkXKKcoV6JnvGgGIcoZRwsSI7SgE5bL6GTC0Nm5yt2Gk00Cy9Xxa8rg6/zvDl
QG2UtNhMdjTpIMuBC09iaCApY8YVvSZmr7ozCNxHrxjzaiz4Dbza+lAH73Xt+bg/bFzauYQ8psXF
XpSAvqNaQsR4w+5QXTpSGQSPktHu6BBYWlFNSo+L1YeQQGSqN5TPxl2KkH6EsFXk6N8HurxQJqiT
O6Xk5Ef/InRPbgzS+FKBjjmhRB8fYZmgNvXqrKc6Q6jL8yeEpdOGc5wmtVXe9nj9m5LIXgBOMpb8
MbE1SXjXYFqXNrWpTK7XDs+Ji32AJcyHNf5/Zn9PSi7Y6XFxunDvXk4Ynvh2kL83I1gv+ehqKA7O
2Qu1PBr41MEpjgoIaZTlQSRJjXUlhPs4mGx7M8mcwLJE9yqs/RBhU6dK/KvCRw/aPk+53R8mGNiq
jOI62qfSRztWHGWMADNZ9BjaAzngSTdCKkMRrMdItcLoZPPjQjS77yoeFG1v1UbyGur1XotIWyDJ
HspWzdEFBJNodqt63VE+ZDoxnvGjvceu8n1GoBpgt1vNBnkcrsQV13MQe6PTbTjYVAiYCLGE5tYl
97sXq8nLxMy51ZtIdUWVcCPoIE9+D1Vc4f002wshTC3dMzIXxzFo/b5p13+pvpKDzgvuzehoPKoa
IEk6MBKpbvQ2zDY8lDo6Puvmc5WY6jrca2PAo8jSUqhfttgZ6L5sRO9a3uZYnar4BgVGrhfCiYqe
3ygrwn9HZFizLUL89gip/lemRtZ74rIhX+PMhefQ+eMEQcqZiL7TAMfzdBAeXa/TwiLOBA/6KJRe
vOzZyYJX/J8fbNDy67vc02US72GaKKYN8MXN7EjpdnhZWq+4PqlxegnKsUEBglHnGDfeozXyBigT
SmiF3H6V8g+grvaIR5hB5rUn3LVc8yULyFnX9zV5l+rg48TsBQZYjsDlPCjlQOLNzO2GUpQ5EjDK
AzuDYrionOPpPE03b4SbNk55k2MzlTF3ah+R1AjROjDqTzf/CYF+ImXS0Z0UBYYiq5cDj4y1bWyk
gXCHUDwWb80lLuVLxkUFnGGm8H9DeyCnodav+ySj9FcyIbxVxQQgpY6Al7NZNbiespozadO79p9P
mpdXx78wfgnJBc1lwETxrqso/ayqS7oRWPSThIXHo/5pEHWMDBBLFEMNP5UW75fvEegmnxt07uCN
QTaXScl7wNFapyrGaPLzrpyEx02+ySuMlQPWAXSyVXqDopkDaEteT1ZMstWM7L4ONCye9DKKr/wr
QvtXUQ40GFuUwdf/23h3e7ElvfRTf3MF2Oo/rp5o9gpRwOa4/1hbiO8q4uF0P6is2WOPT1Y10GK0
neVhM3HUtmXE0cGjUjL+dnEIiFutNoyAVOjmKkGBtSc0g9InZeL8tyIag1+8pddzmBiYs71u7po0
cJdknvqhQWIR7ITugXlKOSv1N8s67F7t4DSWzRPk8EHI/Hsdh1dmJK60auMR6DYwCArIGc/p9IIn
WGQl9inLkU845HgNZzoytZ+ylufVQg3zadxz/Pv9YHtYz0lH9bbWv3eC+Yq+FsPZWupDnOj7Dtmq
wn84XvmNB0hxgVDn93dxApef2Tcvz1jKdurKsmwNrN8/I8zxJoRcRZAuVbnYdbgR2sGDSx5iEbUR
pNvYEWu4mFv+LvYFTyEuwh+YHids5EArdUkQz2t0pIRmZmGbKqNjWI1B032tVRwmbVax/Jq7EPtq
5tmFE5fyYvTJ644mOPBW7Lq0JBtdHByfaKne3Epeemp7FgvBX35s31Q7J1i02jk4JD8JzX9yc0L9
m5hMFjfwYWOMxh/mvLLbC7E1GE9fjx1rKlnlcvqZGNi06zKO8ewPuAuKpj0gJ1qRkgGluodWMbgH
cTPcd3nzbxhUsXqvvhPwp95VHSubf1JYOubet7sG44LUEFkLTQuhBTMM0w3L+6G+gDTpZJ8qAM2d
UiKqRiwCwmbIF6a0xE9uxSh/1LQuVS20oSyTDI2e9Xs6STMPG2rr6L8I5z/pXbbpj9kzK2YueR+d
j83P6iIlAf9He/w4npmpPKouxJGvnE1XwibmfIW4ULnVui0H8bzo3KDRLvYz+dPJ5ebrjZyZtKfX
tRGMC3wp7hPt65MnHYS8dnFEqap8+rADFNIK2fut83qZai1ZC1wyjMsCHhyCX5XBuh74Ud59ljLo
mP1rkbaPQEp25Eb+5gomuC9yIuINNAXEwQ8txEzuC8ej54ReBCFU/KdGlSUoZ2K+U39CKjxjEaxF
3TTqPU30W/dToPY+GYZ4Aba+qpCf97+/NZDtquNwtRCDRXlbW/OWDgQb8DPHGgpa9dJzT1vLFM8r
jMQJi64Jsy8M9NObluKig9QbOQNN9A/ax3lzDVtNxQGRTdOjAW2HjBbRoZYbzxKyhqeD0KaoULcg
1+vs6RyI2r4mxmfNj+NNGL/AvRRZlOQefsslbkOXdkeb1Ye4SC9XRokv/BXqxN+dxjVsY9bsc3Y1
y43H2M5x7RzDKNLOHRq09sPn5f4lWY2wDdhZb8FWZMoTHDif5aqkviXIs/XwUlORdgDtbu2UQbh/
JmcCQPzgD3djcKEuZHgpIxDmA2tE8B77hQaWffkHdzIMbTqFgPgNDLZ77fsE47+9viDSfuduJbrf
xdks1h6dbSQjPIQXppGlzcARKwODdEp7e7W+JXLffYNiV1qzDfxYvUW/Ovusqn3NMvniFeI/DNnc
GP49FiUTlIAVA/O5OX1/Nv7Fc8O9rJhs89033UwDhXFxHgILZ17XVejZm/HAAiNWSHmJ6moOP2vq
6qlHR6ymHGGUTFjz5BU96eUPUjMH76lU1xFHV4jGPVV1Z6nI3528hx+sE7OI2YV3wQ4hGUnvcB0N
I/OWA3kpxZWyyleSykOjJPyA+4qeyOhPYVGP8rj0ByRUXbLLX5S9OjjHi9B38RlDMEM5qxesRhBb
KDJDp/cJ9yR4+9aoaaxNikCMsjTcv0yM4lg1uTFwn1fOJUs1Frog+tXOPzyz5Cw80jRj61UUvfza
Sh5xrdKscOI7M5tX4TjD98X8qoMv+Yt5bgGw0dySBL/supD+z7GHLY5LlafmOh8xE3m0LcKoxsoy
JlG5XRnb4Mb3f8szqock3ljx+Lt+uBiVSONr10B8Ch20Gds03NEjEq6xNq9gccycn25nsczZVObP
hGLltZlr91EdBoM+Ce0pD/E/P4V/m8HcC/yfyKE0jHGR4NWfWpKCru7qJyfI5gXrwiBhuzTZUQ34
OttPksuoHQAqZope2A1Hq9lxFzhSL9j1242edjCjKwC0NN9P1bc5jjizxIVN28wNvoYgVyqU1AyZ
ok09WZ2wGKpZ+P38kTMshWw8mxyPhj/Aeu+8ftqjzWw/SO4gOQgZ8TEsdQVSbaWwguK4nAj+9bCP
BOcZPNLCbH/YmlZpcyMpyqundvvJvkKqf1CxJIg0Qggx2bK5cSKQ6HYnrdAgcNxbk3MFFgbBPX81
Or+R5bRQG+sRgHfB0aJPd1pfScM+Ia97KhT9D52WxLKx6jJsm6lnuQputvzg4+sRsiCZAWl3JnPM
tC0+UmL6P8z9czD5Zpf4n7kmd0PfFe6hji5GcaAAXo45wKSmjpAGNNsL0uHt26UAj3jwK0LHlLww
g9gJTexHWfmBsO2lMB4JPTpVpt5hvGZb5TZV/T5WRV2lY7cx1QTHihD9HTrxP1xD44HeCaVEJuac
5uaQzBf9holYvz4bYAgTMHhs/v+aPKeMUeymXod0B/XlJy6Uat0ydC9lhFBPG63NMfjyMEtbBNOz
qHD8hTAPP2FMGIIscddOCQZKMOMPmr0fy7IK2ZMqWTM0GJ6gcVe+0HW3yUb444mvzm8cDoDP04QU
wongpMRaeI3kj4s5OgRYrj9mtQfRYC7wPbXaE1r7h8pmV2urLPL78lorg/CQXJ0zvffY9v/poWUY
cVtM3bpmJFd2l05dezupcu9C0scNRLgNuVzwKaQWtI919eMDdwaJWMi2+gEJAIZP1GtLpMUMzB7b
oZ98WIpRQsvOO+hqr2WmGnLIu+tgKFv1fnErbk2nzIQEziH8ntMfTDcaWH/hGbB8qXvsxZkztXs5
pUC71CFc3ed5LAhIg+xwlW/y2vcbCYQXlYeXnXBCp9kJfA7ltLkzgFvF2XMRWCEBbsyySzzS8U45
hquLrzVNnVlJGM9NvEVq1bM2CkpvH4MOhicIgPnMxPrNuGyF+cbkL6gtYsWCykuM9ATC6o/CnEE2
d4xESwEOBKVgAWv+scDOyRn90yl8mT8dO8D4gjm2XTW2Ohw+8PyGNGeAdhbJ2aUApTiER7VuCVKP
d/oAGAcX9euudCIDnclYFIBMcj80vnzSrG16ujlhV89pX7elyqOn2NqtZRvhklKWzV4PmHxp7E1l
mq0MWSEEiu4W1bftz21iuIPTRboGXcugkcccWuIeNo4RmAFAcsOXgSs4S9P5IxMPB6U4fmbjnfit
A7ng0TZbIcBlR/OoQN9rEIfny1kvS4fisWXuPX3O4eDE25vDNabuSI4CPEiaH2q8NYup6dQWmAuB
IK0fRLvqg92ujTJDe9Uj0MCbamg//rXhmDHbC6cKpxVfj9FBYWdCNIy9SajZqPDO7KquAtlZyfi9
XGYPmyWuU/+FrVTqSKgub3AKDMcfrEkDq4z+9KCoWykMLXWSx2nn7vIsLfyfWAWzqwSJ1+GAlszb
U+vejzdzA3EFYgXA9ACKdD3jwRp6zN+EHfGpxx7fhQCglBdC8ZoXM4N6c1qtwhASWYgts3Erj3AC
R8tRADJrmO+etatow8r+Vvq6DoutxYZFn7Y/0dx6w2hXzqDEe7y5lTnl8cEFs8NWOrwj60CDnnQa
mKUkdoHV6X2Mb3iKFZQDZgMdszkjaTvDLuknm1E/kYG0Qw67RhXBruc+ecWiy2qrIML2yamnzCgn
BXAF6huOwOe7+KyMHNEuIi6baxpp7BWhYphH3Q2cBDIo1Lb5r5alLVyC7KUQ9HO50IUWJKIVjHp2
ZJJ5T+xKtoveY9q/OT6yJzuWK0HVF5KGTKKWDZLthiG75jzegeKyxqu55Q2WEkh0njmO4rURmEn0
b2N3JUZFjFh0FUlw3tcp+0bLiiqrxNchUhhMBCqhgdsgZawHHB7GlToMUu+SdJQHy1SlOpJRTZ23
DtJt1YM+wbGpZ8MXo3eM3wkwyo7qEns4s7rUEf+KP+/srBvyPzBSaTnWhk4US6ZVnuj6Y27gKYuf
Afh8mYICueR8j5YEUD6m1Ac5vcVZRH2JzZQv8FNHCUg918qWnlDDOMf+QV/Fh5+KpU2B1lcqR51S
0voH/fR7leoIk0mHtukgTM7505eiLd/iSA2hIEIZy1bN1fPi1DBHm5lYAzMMIBWT+usX8O364skx
eETDEexEyxTAWgxUXK6b4W6tSAGEg8czjgTnGrPe39u0TIhX0PtCZ91UKbQlBTXCOLfb0/Ff8nUX
RSn+z4rW64CTblxexzG7oqxdGfN61blAE/3Sap2Y1pLwi9WCoXL8EDvV0LLRvOtMv+0/2QMjAHB9
db0GOaefjyKsSO6YhN/sQumv0cZQUlf0lQisFj/xZ1SRDxKB9wuVC6kgpS+WQY3Qgut2uclZLRcE
LQSarYx8hO6uNOEX62STTuIbYa1RrRl5bhJKI6Lqy+aYj6wcpv0AJeG0TQXXiq7d9sk/gqQgVXZ7
f+sPi5lGWYlXGvQLNgVIE9nP3Ws6WQx/Rmd0UiHw99GPN5XC/tq8Tk4s7GpmPfbRSWAAXK9GbTo1
zQ1RkVagUgx9hClETM6rybZl3S4PF8WbCltdB1Smx3oi6Tv1XD2NEoLzHgI6X1BS3Zs5hkdSO6Xg
dB4gxwvl5eHHwyATPUVUu1LlBkWOUDPVEOd4H3zJVg6WtQvA3niFYadDsH6Z22JFfGJYt1nvN9ng
vVlMFnVMYEC5CDSKHn84ULd4+gB56fg5qya6WXhVy3aTbVbIHN1DKM9yxX9CXsO8f6ti8zXi2aKe
w7qD+0kDQeoMzM/5g/bPMuFHEpjOh2XnB7CQp1Py4iM+utxhRg4pyOw5GcCeQSFwMBI7+dMBObxm
t6biPnzellW8J4EtGc1nyPXEdcRxIaypnzJTNc9+ae8MDJpmaSfrdPC8Ufjv/rv/Q/nLmMSIdHTN
/osnKp3bXSVdeQdnqHu05sKmegh22XnR7b657kcu1mbw66F4k80tNEByxgNQx/RB6sp3mgVQIGZH
07iT3KqRLsntAZYXRBm7KH7X5aWByFZ3NJXlI1cJYJTm6GwhZiQ+ckl2Gh/NSG2+6avywPNaKxdM
MOaIq+6u791M/PJOOeNVoAYvgENIZG68GL7MZwUcoI3r7+MV+3zTQUbaSK7KbNcqQdgAiohxjwAK
ZtAfHJ8+ieQ+QKtG/kopEM5qpHj1QZ5+0PwMKpcWe5I4Y4f0VhTaULl4M9t8d8NmuhzB5LHpjQvy
mGvNtxHa+iG7Od6yylHubx57ur/cSnLR5yPxDJFGoSnpmalHr3CtrH+MsUjp1VbsV3nzcShdHfVX
hZ84eIM+U3OQzFS3WdTRuIDDAMqZuDbC6wbLEqFqc6/mV6e3pwgu4VUzwYVI9uWUvKMqddnP0klC
4b7HF0kqM/gKwNp7vR4g5hy/95KsdcocdgH1qRZJqzU+ak2WXpuiLfsg/lv7A5zWKKN6zntiDr1q
U4g+fDGnbPsRqVU1uIgOlGiEZ2nFORN0JQ48k/MaWf2z6/TbqNZ5+9YsIkT1SWbK2hLk7i7b1fBg
PXfcerV2GQMYcpQTMBBmsQ7fdvjirxgtdAiFqUxpQH7vwA9PGjARIGYHKxVSKjQ0MYywg/YTXWTv
Isle9HcceZBdJHC/qdDYC1q3Z9Q9UMdawcR2kz8t3yFB/FuV5ujaSYkM6/Hn7iKCY9T4nQFGUJL1
Wf1bFo7qVECB2S0qtev5P+I0prHzsjRCxuToHnPKxawrWGZrm63TtsC4/K8OdoKygSaJEKT4Y8yu
VZk4U56puhiRi93WxAZ00HiwkKN7QINP63EhFyMOn/PAkxC2AWe9tefb2j0w7lVe/wAvXFHPzjak
ztYEUpB7JDBHBRpJ+dthbnOcEN2pBj3XZTbcdOWxPHoaUKv09mxs1Jcu5AmbyZ/tNX6R251csxIY
7dWecbkVTtJtY5bCqCFMbui/5SRciTkWszpv/jybDgvVuYrpCuQLosERUFKp1vzIa0+ac+SYUq9X
ASVi8SU2P+R7Mz9fwbj8x0e4gbHPOb/BkYz1LG9khv3l2Ir5vFdeUXiZeAu8dje0m42ydTrYzTO0
LEmRUndJZWV84uGfmXPGVE2R30FXvjKK7ITJzYBZc0KoPoTDMPMW3TsURGF1pvm0xPaTsuja4TPG
ZosWVO5wbfXfpFRaUr3bZz47OmhopWyJJovcI9pLR8HB15/YUwQ8FS8lJ8aYM+IYcVshdmzc4T/I
AWIxzSl2Wq69yhP6txtgCnbJR5IULxfA6FrlCu6bjHenCFxOcky48nzlQmkbB1GNLyzlkgG3nqYG
1M7veE/9tNH6dLdjTcz/tGBy9LuzmCr0PJDK0gr7f3OBnza8hV7qG7sdcc8vYi7GCBAPHGlsoSeN
rGN8sXyjERj3xsrZvPTcFV4/+mT3dmqyoxVwuovM7dnQ+qV9+w1NXKr0AIH9tq5rX3YcpK/BEHgA
hJJuFBetMmGoO1Ja0FiUp7Gq9/2/8Rk6+wKLVlwaNdx4C5Rd49BM56keF7bSFYCn2KxcPq6x9Cq5
1w2VZSJDniRz/8mxwje6A93aDt4JtMYjzrqKiiC/i1Yz1kmwmrCmurWoIEzNbfVsLlwfbW1676Bc
cMcGZ6EK4WC97pYFrgFeTs0UdsdVjo597hK8DZ7bv0k/L493AzrOw+a+XgOKF4y4JMi/5wkoVCKE
SNBQyasOyb7T4XZLDeInYPOuyuxuG0Q37+2kEcmhlNBMCl/1huvyP0IzXKOd7CWR6cSCdkHiJemD
xwis4pTFY+S3ASIlATrJLI3R0SJVA+Omk132o0blDf3t8R2TJzkoWSEfObjdoezu9Kv5EMXV9RY4
lUQJJk4ucNESZ7tI6oOoJPfho0VNi3o0toVHzRq0n3aBP4C1cPdrZQaK3Mf2NE7HAUR2MrMkooUa
bAhbTCTqCfPf0kuCEeLVOVWC3RsTPAFtASYHF0ATch1dR9e4H8lUlC9isHW00K4odkiVvjCemdjg
hvr+lFU3Y+hmpVYkkWvJ2UE1gxV2ybYhYZ19znQonI9F0XSsqGdTyg/0OcDw4auyqyer9AHAIZvl
z0HZQ9LggOKphdzscczf4QBywgRAXUV6jITrz92b5iCyhhM2F5aNdXpcCDqgbwj75n14fc/HalvA
zx4ilEUvuDclNZQi+pdu5fpS/PfewQr+MAcxNuIRXHYUVOLdfJhIL6LkbxmaTJjNU5l4E2GOYTkd
S0nmNC4PPA6VEOGohSdU8yDOI1GxVMqZWsz8c2uZCDEMxWXC6zEu3xHXn8sBtSo3iOxEaoDwPg4A
94VSO1ciyIKgNErdmv8MIt1i/xFH5aX4996YT7ZH8uKi5vuLyvJxPoIANRWr6CVBsoodnTQyCR9N
8DjZuSkjvXiXHUakWTIIVho8Wy0zwe+vs4qxXfov2QGN3DZkeWH+UdIAmfSmfH1EbO+puQQwiVjy
d4ZtJmf1J2NjjDJHqBLrz4Xq6RF2ERCSFj16LiUxm8EUPnF7jp9GO665smrgpav3NgJ7GSOsCQK/
60hIv/afqxwpDfDItzLEbMaLlMPfiAb+KqQhUOjEjYAQsc8Z7a6cFsnZpzKcnONOJrmbvUO/D97Q
52f3qU+aTDoufcstiaEb3htzruNbG+FnjMesFkj0UTd3rKDqtx6gXFqj8w4fjil2fcebcKmAM3Wn
7RwJ4kj52Cm4UOR4GjpFTMZzzcEACiLoKw7vPDADrtyy6aWvQFpCI+Le+BqUdd9loFLGPZ5o2nAm
Qm99UbpeIh0gJARmYBPDZIUdPqnaOTtblnLmdc5FVnkPL7D1iEwvUpC6A95hWl+jaArFEhIr8f4P
klOtqbf82vl1qVgkmucb81MP1/5Yd0fLRXUY7OCJN5w0mr6vy4x7PAJp7aRSWt9aOoFOEkOBJ/nD
wRC2CgraXbzvDPLmydvVolX5Al8abJoNqm/ST1FyvGXAhDIVCKG1RDUbubSuA9BzFfP7Cr41Tfyu
j7W7Qhcw/WJYKjRYmjoFLQXc0du/gy/HgeIA/ypEGRKY4qSjxSCpNgurMzadGaSC3v7G8LIkz5bR
J5HqGdRpXKDG4fbktlhIQ1MFHFq439xMfzwzGUsM9ztHJUPktpQlgX9JXSTJvi68MnWguWi4SfQC
57yQtWw/4PK8gBtZKo0o8poJekd/y7VQtbeTELE6mBkFY6VJCqA4vXybgYtjftdMYth8tMzfuA98
zRq189e1TuqteKDoEA71BkF8B8HiIamcxdvPH4voERLOZkE6S6ix8DIihj7ADVIS5SC2D0ReCwby
8P1+lKi3K31hjM6gaci9J87829FFqy3ygiMDjuxm7h73+ahrnuDE9poC0ONFjxsJjG9RFsW+3NGA
uhhM0Yfjan/ETSgxrd0RJccFVDbVTKU7YD60hNqhZE7/rZ28oicnny9Q0ldTtr82SHc9xABnj9zb
013VfeSicb0/1hWaB8I+o0xY41OmTaC6yrJpphCDWuH5GDw5MmDSY8QoMj8XTXXB0jZXbVk7c+YJ
M4o4/8gWSj6BIjNAahUK8IuI1MPKI/MfpNhAeQ65+FqbkHqg2uX0qnWx4xlwWIvH4iSHgf3keeJu
0uwd0oGF6Hr2UFn/yix3SqgTCMEXOcBMi/gEIAgQYETMTyEKR0MbBBwdpA9SHNIorba1uTaHl8EU
BnVOPX99snnSEiYGz5HkcAQ76DJ2A7lNgIfFQqtamIK5v549yiFZoAdHdoHjnKVL51zdXu0aREso
KrdThP14jht73wbOhnyTiNMIL8hX9WnWbZeHsalEr7BV3HlUY69nZGZ8NtnAC/XeaMq9OamVBwd4
XP5RmltskpyG/GrQVQhYfs5Fu4htUaD4/74AaTfzxspMJtfBZIrFt11BeRkQcRMLzeY6rZ7vB+NN
MbPivd0rwfwgKKnycY86pLQ0M5XjUAttJK0cTs2I/mLkwInpTK4FmgMGUMWRiabGLAKgBrACpqFy
dhbJBzfOopKVBAbf2tbgfiGCCh1R/yEhd5+ZydmJTETa1FQOf2zfo8S2Zj0zDP5ROQ8BQg76WCw+
cmcNQaIW8RA4ZQbE7fPEALl/967evHyCeMSg/B8wBxk6t7uYNkg78JBdPrmx3iE81k+Hjo1Er0sZ
aCcx9p9iEJVI57NwYkZaMr2ipujONI/6v/3wBgswl8zZ0EZboYR8gUQNR3asxTsvNOCp4rmgIox+
zf7b7cPP0/AZqDhxVVAi8qfI6JGcwMQgDNfnc3OdLzHDujXcZ01etYD9ogq1u82YVvT1qw0dDJGn
xYxs2coxbKTVD9cP8di0Gkh8C34SsfHwD5Iigf6xBodUbKlfE/EuoCqX19UgODRG37y5G+KlXvsV
Dx6SbOKlk2726DeaAikDnBvW9saO7wGcxoVnzxTUbBruJrJVx2RzFav7JoaH2YgfXQAmVx1wqjcA
0nN2tWg3jgmZUZp0GjaGtww4KkC1/5RZJ1VcNxbxLB1+02fjUs9hVhV7gB12io55QwBG+IR/y8Vb
POLYoxyh7S/LYclnImEP7Vc98e3cEfKV//kANsMqoW6EWfBUFRApQwMH0o6aK1xZfXsuAaQNyV6/
E2AYrMW2k5W4SBF6FP2zgmcrSpOwHVToe9wqF4evenzre/zw39+Yk/FZrjGmUx2T8ixpabIDa5aV
fg0t/fRZj9DLifrisz/yEpHwOjcYk0w7K19kBIJfCzXRjUipHQskyr5gdVkKJvaQAnij8rKTID5f
VZXiULSpF3tguHVDQ4TpxBcZUS8ivv8dtefFbdEwbxBXG/CaJpfkWtJXAPn1RvUVaZL2MK4ZpKfI
CiE2YEQvtoukbI7HyTsuBF0aP3bhpHIFojHktISuTxnk2t+yQjJFKWp/GRpeiqiwAOdS+e3a/aKX
Xtu3W6OWfIxMpGMPhG4y3DWQznNHeWO/US7bfwa9Pye/ZUHgqtfcgILCDroktufMFo9amQqX3L6Q
yzK1sZDB3bJA9cc8OR4qVU9J6pMNXcXgDqa1kDKiv2tJm0uYLot+qovupsY+PoJujioKFz6YMmvQ
GnStk83v1fK+ZCAlSkyv27vuqFJGunq5sW42ckZ8O79KDSKhDtFiDtzmm/OmCQ8+ddmFRFayQAN2
2c7g/3UJNpckOPGeT5doarBNA7iUTcBdkl34Rr9zBuFd8KFq2ce9OODJ1Bf38Y7X5feHDRvaK4kw
Kj+/CF+LPXXg9dtm/IYNq7GTIHu7SPvExONnyCsbbkafk9+ZcYRuzroWd2QIcuHYVdBhmd55Groi
mJhY7gOiYTbR2yOF2wKIGWvmdQN/wwNBnLSxBLpgEPIoRI2AZpd3iQjf6ey2SV5puDl3ZLTEpg4S
qqnMdb8oGZLVBH8QNwZrF1SQu1VsTmiyCFjUu+2JBgEer7IipD+YLvcsMDRS6Fj61wldFqq+pE00
d73fFVpEo7viBw0ahCMZbXUFB4SJH5njspQcVjeZt5eYKJ1/qnbDS3ElwuC3Voveij8wwEtUUhHL
2nq8o3WtR7rYE4S5vL3PkHWnls8D3LNjeReLaSPsMN/ZaIYsrhtNr8FZezpaWXY3TRMQhrSvq3IC
k+2m7N38b3M9Y3GyANRuEPqAIdMRfHZsgu5OpJKVnFAZn1MJsI0wjZ8MUCcl3xoMIfjHXkZFKDy3
Y/csbXlfazJ9VumweMMEaQpAp9400L14kopM2iT3Pu72AVhTXAvMiyg7JaDtifNCdcsJ3cWQ4c4+
jKXl1P8RHBiGk98ax7dnyeWZIRp5E909Kfh4xxp6qaGOlCGTVqZgyJmrjSJupMuF2UQx36nv/wf3
XNHUeqIwX1msqCQvMAuQHzpKijElujmDvCWwR2uGQ1VyE/VrF37LAtPe33T+rMXKaf0ymu/QvhxL
Qj9OOfNmPKlRYrsTnKIe1Ti6+P3nlcjLZN769WScQ3yaHarUHkFk7mOe+qk5PWoocueYMc2E0Tbn
D8zVzexSniR5XafdOMOR1VbjATgLSC+TBHY+nNieNg2bqmUuRFct+0tRNEJJX2ZE6eWgxAWX8iC4
stjlb0bWzZ2ui5zsKs23VKwItWbUPmyb1B6OR7U+/FCpT/Qfq51XM/GMSCONQhS/RM2Qw3bvqHIR
TLLqjm60VNcJ/LjtbpM3Mn7ElpNiQLP+GDHAQqJH15Rvk+WSZlLI72Rlc+VCDTgmJcLmXOOoSQcE
Anp3qNIOXrCubLQM9X2B/lQdaIHacLMF4WsCR1UJ3wucOBg4I23xSkeVwT3jXZC/kr2DX83iIkRy
pwbZ3AHm9c4ViF7qSptE0NZwkNRc4Zw4BGsT3Umzcle4JEDKNIcWaSUEiIBYbaxcbHlrdqw3n7Eh
C/68espUakoK8DSM1IZC1BVuU5jFCidH0iBfCiTa1Ro1SZHT+TNs6gHPubtOugH+upjUuCTMPKFE
bVIhFf8kY+ArdkJRkVKejNe00qP52TKNrh0K7Ay35N38NuM/RA2IQpjvNOzVSOzB3Aw9Pkm0aa2y
5ovTQiWkUwhnKTautCTMAVAavOiHkhLe1j6Qe0OjAqAX9waYhQocAVWUAuWEsxZw+bvWFKWozi0a
Tb1fiIVDfMnJlmj9TfAGmQECCKBbnkiMZ63qikCBIBPNJzoId68vnYglrSXtoxbIaGn4Ago3noJk
gDnzktpgQmpAK9pf3LGRkejaxo8Cu/XPS9Zposc0tZwCNwXLVFA5OLt9NDRuHnzR5lRlYDLOscyw
lTqkby2RwIZef7P0Y+iS5XUyinzvAEvLq0pNucHiWqtrxyBo8047Xsar8S1I3ZL5WkrJj6BgqSSr
UTNyxHkuP3Qtjs8qs7RkAd+OAOp3apGbUHvMUPbasJt8WUMde1xFNI7HkH9zm1seC0kaq+D5LrD7
USyF7eAgySEZEir6vB8fC4qhYW386MNr3YOfh6OA2Gcj9sFWw6xvQUdiKSdf5Ih8wmjXpaz+/LST
B+7YB3EIUXY2tgvzSukwesVoLA0fmv7KRC23p0xLGPJCGkoGSgSohsYUC0VetdYquA4BlQbUNeDD
z1nH3LyDG0F6z4lZUNC4umo8joC1Fk+XhIebVeQ9NVGDwXpuFcVDj4DmIrfXBFkOkvElv2i9Q2tq
0F2pv/iM1sMzWWXnZ5+Yf+8o4uGrY/vWF9eaqUGN382wFtV5a/DFLfruFDZeXi9w8agn5+O/lzpq
OKoCqvnT6ZCzb2gzwiuWv9TDsalczWSb9ycK+XC8Hmvci06rU2gzx735w/GL4OkFpRgqF1czQyRF
e6+wxpE6XuRHm5dJiD2C8mj1B71X7ZBiA85DaQSoJblGPC/gTMUdUn0zpenXfxRcbGfq+CEwdIhU
3swG1e4WpMzj3N9G6/JwQGr8eQjzFV+7zKZlZ4N0VFSHeM/+JY0HbFQ2IOpiiNXXpNXHI7Rn58G5
tAdszvXFByEdqSbCBn9zJAAhuXCtNo9MKHO4Ipt7v3FVe2weDf0atb6/UKHNW/QCJDGimo6rNUd2
beSWR0YC1f6ou6OMvoijfNP5dWs31q++pUCX+hTnQdUza3sIViPUO+cGKm4H7kdr70crjuS8M9yq
Rig0b87SWazQetDFYfhAlvYdhB1gLNn9GzPhALORSfpmDprERVszGMorB98KkaYPJleXKDvns/UG
hKrUTnN8FAIDxcu/28K6FOOwfQKt4lUnI+c4332q9I5a7s3BV75THZhnJEI1m2EderQKoPiKuxYD
j8RiE48PVAb6unNOnllTgFUwVH+4+Fcv5y4FSaJcLyPsGqlIvGJQU7fnmszMxm5epuGu0x3tzf3l
N1VXZB5YBhavAbIwa67lK00uD3XHJGcaGIJTZFMVSkm0Ro+q+SVL9OcfzvLTeDLnrsvfQOQ4hibA
gC5vJBaZp903KWwCOVhrjBu38w/eZOjFLInLNsmnoz9CysCYaTcE0DcrZ0TEyN5OL04q/bsesmUG
ruippiYuMu5A/CY0Hako8Fz1JPUQoBI8+zY7baFqCwvkpVcHiqTc0MKUGNuac3VXzCvd5K2M4J0z
7NJvp5aU/eCCpmG9b7V8a5zP3OWmJrTWqCjXaRdSkDcGpCEsHRzP45Er4nM1vBaQVoIdC9I6/Yl+
fj3WiYlbBkzci5S1FUAVshxe7qMJFISbSgdtA5hmEUVFRk+Y95wQuoFcNKLbucncVAD6rxh1F/TI
OqnShi68/NdYotVI3VPEhFIOfwe/3jAJVWrgcA3yQzUD6VTVsSf5o1mtreB/7nfHNToWNVTmen59
RiMWL2IEI0FjCVM2LNlLytgvKoj0MzuXQmdEFkDxv1vIKn73YpehQ3k5fehvULeBSXi/SXp5lxOP
VrCzDMHk1eSDmYAq7yEKbvgtHQ5E9VgNelDReZzrsNEIzgiN5jNinTb1OoQCJExnqaF8FMvw6l1M
dI2GCqSk2XL/kPjNEIuDn0jDjiJpeLgwtAZTnSBArMCNPS/Chdwfqo+uAE83wJ7D866C6YTWKIKz
YBjK7SSDoE6eCX/oCktmWKXL7NHHEFG1PqWLKBZmGg+0lOQwM1+pLJgGd7Jitw1lwe7aS45Tq/Tr
iZGoOasbWnP2/KVK1Uk2PiBLvZCW3RWqGjlYd6cqLDd+XfiJaFzJTUsLZ/eoeTWZHC0BmCgYZfEk
JZAW0zufDOOEc+vekJC0Yr5sv2h5yAkFP43VB2enbLlk2rLBJahJWImuwtoHeieg3vhAv7fW5gOY
tR+pgYvHdHmqQoV+3RRBJNtqWzVW+jXfBfp8Pgjn0cTXLF3FFrU1YoeOHhYq6Q4+Sxaflv1SZUwT
e6KXYPUC3YuCyS6rUnM8UFWUry1uLqU0k/p+la0YTy0nMamQ93pkxGNVyM1UmH0QJ6S+HA49tkkv
nXEyvMmpcKP5RViIaSKjyEBg8qx+a1toT0BCTdJiJwXEnRYLodJxa+TcCk9JAhKC94vjWPq+nvSc
IJ4+VRegfKr1n3ynfZGXHYOsHb+zmkGHlNAVbGbrcoOR5UdCUGwfKfIPwofWkOraF5m2B3y+BTiL
1c+Das+CnUL9iHnBQFspTMFEDScnZJB/XVwRCAvA86uzl50GwlWA+JzyD+ZtWnSlODuUoWEJxgX6
pCoW6Zi5wCyNd1XCI1RLui+W7rny5t0jvGFK0zC4jAfGUzPIGb5kxKSg0dWb5knngxRqed2/jn9T
H/PH61bkJB3WhFLOBc8pPo24foaMShnwuPUD0ZEljk8nlIeJti+Hd5ffWc5SwgWT947Rl3kPfauw
2Banfya8fgugtUVsTN83dBkdXGRjOpCedwl6E9LLetIUuOLqmv5wnzJab2QSt6+AfV69yO43megs
b71BMp8EujlGcnF/kA46Y4aSsQrRQeSQ6TdxymawYIT+cjqzVrLOaKJ+HioQfQqnOKMA9YzMVhlG
hGsSEg4y2zFRlqvyK0yKwGcgYkrG+bxCxz8ji+SAgYkhkzYANi4EfbNqHHWQE/1XmRWv8QE3rxek
aekUhckC4oRFSMTi7ydu6FHdc9A17+jlNk7qDhk1iaKS/125F05J4fYd6/M/iQx3TPOPBN5Vp6mx
KAKNhjrVsTRlMOtCUXAQpsbbGzxywLCtP/h1UkI0yUytpMNofI8XwEsjbBjsra3o5Df4tuPd1jnO
o8w7QchDXQndsYPniCaz+wECkpyTa2q4Sscq9zb87vaCleYHwLx0qnDHwdnraXFtZwDkVjPKyn+u
P42mmaQueSVweFLwbZhP9MkQsc9hqPf9h95tc5YtuvBGqBnnlPclVs3QplwmTH21OOn6zlY1Ez2S
3HDuP5Oz/xSLr0OF7xwASJmUadJtYKgk4TdpuxGCQHF/RK+yLD4453uXbp5WofP/stwo31DIdbVh
sTsF8yf8RVJRikzjjUAmDufcWd/sAMRckLX37pwfkSh1OJ5/99Nb1x482Oz6MI8A7kSiMagjmqJ3
6J2GKldbsF5R2g6vmbpdMPsts8p6Vtd5vqE571TkJpI01sXPBaCveAVl/cxk7IxSRarPxgQhPJDR
8nLe+O0Jj7bezQXD9X/u6/IcMTJdSX3vww9X2JJnKI4uHnDNpcfiH5XhorwIYuQMPq85lqGZseIx
rOVb6WViBmPs7g5lDCF1Zs6jmTqQmtzt7e2b9zrCKtO6e5tuR8E5KTvWrr4PgvrI2ZvQt0wANBel
tlwl4rmezLuQowHJmupknh5vWtAHPNJyCD/utUYgrGxQoMEn7ThL6puvuRPR9Ufm+w8iYESIB8wi
8PJHvGMc6dnIXQZu/PUlsyvP3rXse0aR+NUGYKLrQ2jmhKv/uu2bpvEY1V21czzc7REtP2sHGFvj
yTkz/3ToId/RmEjqRfH7qNc12oNS6yyx1BGccT9NhQQOxZCCMVOjTg+gVH0HbDMv6rOlWje6t2sx
eOKH955tNAMx5d0UiCtcxtxGE8JDX52pTmqaWSYNKnIN9YjcreT3c9m2fKAaN0ma/1VT3NV3i91T
YsvuQNbLF35NeiMfa2+CCxXDnvMH9anEl1X+Ci+TGS+n5a39PQla2kGOeqPIxS4u7asFNfgwoHNl
EXdI0WsCpszQd8wvZAS3cFXIScc+NUgz5yo2gQH4X9TVwZgyb5ae8+nlBXa5sD1NDpR/V8jGt9b4
tJBeyFo8dz8xiI+KZ9+PLLdWxzRRyN+utjGwjOxl5bvm1wu8MRhF1pMRujY+qsrSixkqxHEn8Sky
W0YURLg4vBIZJFgqWCNiupm9vEk1W3+aYvjYLWRrCT66Z22DK3elZvbD2djd3kp1VpPxXGsYAXaY
dtNc61kT/GaURWTjXSVGKYMV0B/yolOSzQwA27kVk+m3MXOGtn6m7VVLZDallnI8g49vgobz6DwT
HlwvoBZed0Tz+5cMXd6BHVa5dD4iTekP1afZ0NN+zVoIokR6vpYuJ9bnnU2EQ3xmvOPyBLZZGWk+
k+UG85vTVyioaXq1Rt2qUhYVywlmA8AE8UfvkU7LuJDswgVOKbMRxkuap5lfqrWdzoSQ8MYBtWji
u/x4K9+Fl0pMFXE7WR7c1oQDl/ZM5/4JeVO+1W+b2/PEOkvnSyG0B0fSgAzzOtHOF//DX02Qsyy1
yDIX3fVJ1UtetgEnyKrcxYWqKI2p887hZkMMCquL/3agNoBYhAvEDHmtrATAeOyFcW8z4j5cAfzf
bji7PZ1C45wU8BJlfzMMQCrsAYuoaZSEeJbiAiZ2Mj9SYQTFYFsMf0tyXR2tjfue96rQWW+qw9q/
2A3An9F1PYBuOOwraPKwEhCoHGailmXGz+3DjkwrOdZ8ZLThWWOXUVl3Njy0sraPhcmoAp6q5/RR
EdAW1vER05JE4X5qnb2fjoGquguOxg6oj7+R7mnhm8E3I6gDoHTD7YzibPo6BPPwJc+uQcfsSrr1
EM64VKe4icVmWFOZU5ASL2kf6WJtlBJPNAv2/HxY5vevjllzbTNgoE3SIHmCzRN1SqfDVkXUcX1x
rX9GIJ8A2dErj1KPD3q/fu3KgmTKE14U8sq0sAeIZpZdxe7AfmLZ+cvWGOq5xknbq5GotF0F4NIN
wKlPqea2IXWT9Db7Vchz/grTFDT+WXViS9xBrJaDvSxfoVnTgNp12/uN4TunTaLq2Jc3Sgc9lHk8
BkkCPsEsD0Siajegq8Nl1bJ+rOkiUMQBlkGvG9Qpw8sTwbUbt5xlK+qu6Na1wM4D0hC8faTXDNqz
ZtauBT31CcyYJ+nGQ1UKUNXOlVy4KHXfnfa9/X6ZmdvgiJkdgUdDBM/PkkKoOxb8fEt6htq8ANts
LIuu712E9+fQVaoPPEaJ8R+dug6t44Xkg4alN23qLgB33cKysdTrcgTVZEcwCIBfZOyOzR0xx4Pl
UjQz9TmSDVX8WNvpc/HynPh+7sW0vDOnB3IFenLydLFNyQDyYnVMaMl49ePZ085lbITgotP+s/iF
ebW4OGvcBM/SxOu+i68+OZskFPjWH5reNT6Q2GvOLrQ3T4pYy+8u3AsocQ1RLht+kjejPVAzewdK
cEpocPmdWRSuro4+QOFhotF2LTOPRKlaLJSaD/9GUdVvgRgbouIlZvk8HHiGgR+L1A1ZzpCdGLgU
36NCRmRky8h5qnNWvNJxVdJqFo79ekSWKfaKOOjqntkjuu+UdTkMojBOJTn6js7aMYKrG3AfsB0/
1Poz6zsiBfM3Ee4Kajc4TOqbtGD4cec1kjNCalQ/P3L6p4NdzmQ0YHU4QoLHnW8SMn4Y6kpeSLJ6
9vKuzjYzPqVRbgGJf/lm21oDQOBBOuGmCZF5a6uBV6BF75z+aCLYqD6f+UzrfRTJ1RAJ/BVSGQO3
V61+vIdD9tbvZBhDtuFNECIGjxJMTRKifhcV4spM/jjyModOgc5Lt7Gev2AWtZSNGOVNiLIcR+5P
wQkFUUnUyK350jla4QXWSiUuSPmpdL5L3FrD1rbWdIhDO47i0aSVHYPQIZKgylrnjrE5fEoWTL2G
qEvZgcyGdYN0f9EpoWFlWS4gxQtFeQZ8K2i/VFJjGhl5bMMrifXxNLIXIjnfU1ilhFstnyEIYhb1
Ww035drO93DVGNfpwTXXq/iWQgf7pBSaSnYW1oDK5iOF6CuVywYO5SIA9XXnhfuZ7GfcMbSxfjMy
toFnTQ0nEqf8YdXcpGtVkrHU9o4lftpQJPbe/fC4tm5ivINDXP3zgf7tEKAU5dNqzwihEwAxC52U
y8CVp1JBk82RqIPewaqHZ3ssjh3npWy4o+fLQG4KkuS/fBmltzHgubTczeX1aud7yOubNH3WETB1
1T5ITt1xSErbbtkDg2FDtKpqoSOIoHne0YUnL5bhbMw7aNRhmGNI96kv8uAqqImc/sQnZSP6/p4/
dWJVSxh1QPesV4jY1MwEJaXGVuuYN6IWb1g2/E6DFYDyFaV0DM2EjhJppy7ZfD0fN+yX/9c/nU2A
jN2TacOjEXrWn1vm1HHK2ZB/BB1AsDUMNKDrcbw79nqOntvAClCJm6Db4FbQ2xHgItZOmhek79BS
jwhUd7CPZCLHWRj7VbRw6IXjoBzLsN8TqIpJmKeaEcPsYI1Rsl44/lzASronrKfd7WcshEvW9Icy
FM00iqNkq1f92emHfZFxB/i19GeSeHse4ho52lNQRVdztjgsLEcLH5ptg2RswEpklsKwLHIAbvrS
VmqLfwhnBKMHjvAU7hST6AoC/54ZuEEifnqNU1Nr+EnfTkWy0m2+LKzPo+ZIUbguXhcRftmcBpms
deH2dBup09/wj0swRwpzqrUPpeoSSS7dcSj0EgjNTm7PdTPjJeCOSc9U8RJEl6tIxmOp7XMHbK+z
OqAQV9WnUD7crHkWWnPv06qnOaIe7DwO41AqK0BCPQLZez6RNuA27oe3NCw01+sfHfoZ59vLBBUR
8kYrgt2RfiKZEAXn4JWScY/T++0bqmnBWyPY+O3j3VKgRCuqhlxs5So26teLS8Z6HDhid3oaszNq
jANwFiVobrLprCfd/EpWG3sYVBgT8zlqt6aaGetiPoYikgY/yfmU2EQ3WbUwTXCQ+r5qO7WJAfmg
78e0ZTlQV50eCJtIMF2hdIDYMJ1+AY8sCiA3pdMOqdSqKHW9N8zVMdBQmqbjZgRhGz2f02c946YQ
1wDxBqw8PYDx8mYqcdyR2ncV2PxoahntMqhabEUbUnYBAKKGxfIrkLupDPeCmclz3bfQ+indJzcy
citSSftWnUboJuSEol3GhPZLAkXZAMCwMp443Z8/OHyYSlCdDZ2pqf5dvQMqrU10r61ivNtud9dN
j/kZ699tOrT5sdokMp1DmSU/77S1Ml3IKs3KAImoD4YwZEzutLotwycEakaUmIEUd50K9qKXntVX
5miTgGkanhdD+du0isuvxpgQJE8GlFIW7GTp6a46NZ97o7qdUzObrrmWii/f/1aSdl/AgKmLVy+O
YsgnYnjAGPTKQ6edLr84b5cosUbLH4pIbEHr1DiBntJ5qj3/EtT4PGfiXGXc+dqay9LUArRFFB7P
J9WTE1Rt5fioXeVhCEWSMWyfQaQyKglGsDbFizDqVbtXXhHqGzWgFdcCWEZKgd6MABVEZ+Z5LsZ4
/c32QqHK6P9Mno1kEX/AZdQHaR7S+x/qQ7cxCY1MWUIOB52QCrOiovg5qk93sZ7DB+gGJcEsmQbo
6k6mqJOiyfON+MHWjT5qyHXUPMmUE3jjG3aUyb9PiC7HgCsxTB11wW8zXAKKoNYy70ufV7cSbbVJ
9c8gyjvJnu1iedyFdcxm7tcM1MjEMsJSlIniimty6ajDIz4giTlGEhfvcIb4aUOmnFoOY7JKuz49
gjTtogWHOAz8xBfuiBc/fOYrzvvcJOsLxnQ5ifBSv+3DCUw16k/+0wNIv+wmIhWSBO7Aw8wO0S2c
A2V5LIscB/8s1zdaIAW3zSXizF7vfdPA6M/Pyl3U+BcOgoooSAR/Daml5tnFYCx521vnCqfXQs9K
fGKvZchOzdNnhz/KG4HA3RWfeV9+EOsi8627cxMqjur5Yj5CFaqm9Jc7xbFX1K+5Ufhzxyyx5//D
4vAYfCZGPwzs/xXW3DlsQCXe4kg/x/jO4EtSn4EBnVm3JzHpWXaiylJ3y65IWkZ3cY0OLRDd6Dyb
7xzNoU2JEzD9IAAFkwdI8cU/OcK3szi46Gc20BjRBsX/BRWCPsclrT6Qwo84K2UxQqQqGtOtvofc
mXcGeB/yfFwpikKXyZ6Dekn0+qmoso+od6dHhLbDJEvGkziwOXRIP8iDEvjM/qqyl1VGmHFjfeer
esG23Gl/8PibO9gc5F1uCv9T4uMDqalz0yt99cRUrLQzhQ7/nx8TkvIQdPtPFhkFN+ywea9LCBGW
yulEqdTb2MJydWca3jaaZfaC1CnsfitNowI1bFK43u5iF+n8vvjaa3sFS2HVjYNfIrIWaQg8dYji
OVewutAwsuyWJTMNey+aiWka1wHYGmZfwZRxkdWzjwFmqKa3EohMIGEYLckQeq890wxI55LGDl9z
C9LyOBVYAlbW23a1Qly850qsuKWpSezD/Sm682J1W3ENSNzjfNLmUZkQZML3y2UjaZXwfcpAezoC
cvSOkci4JvZ/WBEW3616QzRVtDughAQZyTVbwkpeNEerFnda6KkAFmXyckVqGGxBXec4VQROjOgl
aRWDdmdpn3nQormIu+ndmk43aKor8WNvON+aBzdRIoeg5GaxDgwOkdXzXXP+KBPBxTtPsnDLX3SC
Zi5LeTLPsgoTkPafhwATZLR5pFvFqT5+NNsYcT84twmJRavrK7Pesvcf3FsfSh0nx5xwceLTlGZW
g++lOrAHlpRBWOgKBeM+t+twP6AHy0o+p03A/ICLD/NGDIUn+P2/0G7SsCh5/D9SI/w6+fmTHAOd
1FWltai6tD5siJbvexboPLmWTuNEDaNpeSOWh2xFQY21QxY10tD3Rpu2rXf2SM9XdXrU4uIHi9EQ
y/+dGW1VY4nOkREbBFwlPFfHXfCSdIuKLNkEa9HHhROLdgLhVBNxXo3IWeAugZWPXAadgd6cU1IU
vsmX7xLW6qLDWZxUBhKkPq2m+w7smL1VPsE5zlU5BMYxnNOHv8a3+aCDgQUTxAfG2d7HvuYGNmg3
3quuAI2aYiDfwg18fG4dwVnXKLQXjvZqhsptLwAyGPk3LGm6S26sLaDSzu6VPXjtlfbTLSu1I4tI
XouEZ5rBgQQsXBbzBczeF8eLmxRUi0YribrjYHFYi4kGRuDnlRr40KDvvY0/tClbciuBhpJRrGRf
KnFhrzGc2IDsK4Z0doEeyU+f3oRPnI7AQRcXgvf8dv2P4Vvwmga7Q0egIvBZAYmZ9YJVgRBTzF3h
aphzZ+Yl8NihD9/94rXFwAPs0sprMEgLeNqPI2FZTg3SHkVuUyxZTsuZB1NqP04n823Z89WItlXn
Z/7V71T84KGk1dxIo5Alzz2/rr4rVqozT+O+/BkcsRQf9w26M3o2ec5Pkp8FZ+FNqqRLhPzR+Jdo
AOvbLVQyBpJ5nPtK+j1sSUnauqb7p/jnWBmloDJxipEC8HxTK+wkD/8gxXyzjn2t0TMBCxmhXmma
vm4QbdKWdhq3r1ngcrbA54ZAdVk/tku+S7Vl9nYD6ZJEBHk8PDDezk8mqpwk+8LCzpA9UP5SNvGQ
THCHhcNkhM+So+ITQewFvlZ0tdBf4WUdRqlAoQ1faodymXFFsvU7ztJQnhmytzWrvMLUc1Ghk2A/
FFEosUVEitC1dpX/3r4mXrATlY9tADBQk323+4SJwH0TOFddM4FP2fvxJCgRTYowPkQ8yUk6Oe9S
Iu2UFo8ijbYXUW3YhYEp3MDYy1e2kv3TtMlhLyOTmnds7mDx9wZCoVsnruRtBTSm1Ohz6PwhZhK3
dAQ2s2l9SGcj7XU04/3IE9Q14z48BpeuWzuhKO1WOMQWfyY5kLbtc0bO4mhZEmbN1QLbdbZysU8P
DOzY9fc/lEVMBkTbrX0O9bVvcsYxxwwIKRXSHDPEN31wSc/cl/mmi3jt+Jj7z6aJ5oVryR9TYMHL
R/OSP724bkHwHsd/plQAZ4TZ9+LbscUb+q2KWriCLxQLOKT+pWy4JTHEU755RryAymSN6NtweRS+
qqs4klNM9vVBLFicrlUpgar1IySCK2vuDuQuO8YA7SVRj2rGltCNnRIfsxeIrAnu3FwLoZDz4vXJ
p64U3OKoYgSfm5y/gXFEFhUizF9ma6gD4U+RG+gm5+4aEOQfnLODcB+k+gzNxwWA65izROa3pTJ0
1lL+T7xpaAZo5XxAegCVkwDzZqRi8mhhqZ3tWK4KYHj+euJ5WuBDz9RBWV0lRDGDd9bCdUTDBNyy
UQFL3Pns85+J53K+qPfAE6WnzX5nTQxf8DZ5ZoJX6fa6CEWG1rSG1v5NqSO63ed5mUslruaHuYQT
oeLTjKNJBfSPvp4hqHrxzX3G3PiJ4ULIMkvi33RzSLz9+/x5inTLp4EPbnqsLMIKmykEpJUkaT+G
SuR/jtdjQ74g94fHncjdVM4bh278V70VrlMPPlMYMWT30eWXn3dJ5KS+S4epBnJEpWnAKGwdnKtl
VNcHvo8qFvZWXldxrdbEvnVk+KLHeeUy2blEUgdkJLGYrYMMkzM/aSaYd7lFT0Plk8+6Z7mXTGIY
0UtI/gx0nrgOCKIe1Jeh9niCwkgkEmCfgXMINBIJh7yWzgsezzDZNG8p9eHXffaTDii1kpiAT81+
3YYr/5pCGhcxYJNjfzTSOfkoHW7ixOVIgp+3WcGMVkODERLlWY/k/7NX9GKN2/0RcYCZ9Qra0cm6
uZuGnoRPQPPT9he7TvikZqKmnIB48fGR8vjMedX0He6um3WY7FilyqQRN6oNPrS2JJ9VW8f8U+1g
KILB9iVsdX1ZeTNUuHMHKkdFPZKESImcJiCWG0fBn67aCe4ORe6gRv8jxiuFRxAAt+shoDuriBRJ
L6ID++F2BibAZwcO2/WKEtm8vWGXbXs0sPLthxy6ypLnGQPMGvJnHRWXNS+jnBPADa0IZjEt9xVJ
cpycwqiCYY2mGGDLJsX/oPABwNJmNtkjSNlX7Z5VjmENFV/ssGMiVn380NN9mhhS/v2uPzklW+Uk
5g08V2uLObLw6pn3KLbVOiSRB8LKl7X686cAAI7WlTdpFNGEfSt96C4ofvrPCI4mZSQBA3Z1zLdR
trRxkRr05UcB6xQ3UfoS7a9ohPHiAxuB0GkE8OsN4MklbN0a0xF5EiK+PLzLpMa2Z6SaN764lxCl
+lrePT/4HZ7mv4Gj/J3uaDFDbqrQhnMjccdnCOlZl91DYIIHEjlO69c0um7Pz6RwSJ7TmbiGy52q
a+MsyH1zc79AOuEuhjRXtTRwtQZUMMexHozM1K/Bf6wEwkBwYN+GD1QMznvfd7KWT+0I/ZLgfs2y
gHURR/F1aob4aIB4hNBgH0EKFbGt3//Ht1DFGYJKr2gIO9O09LQvT7WG/YWhJQuceYz7cWpaNSjf
Wp8z5WWXSCJ0YvXTL4+8xv4zhCbbtPjOwHVD/tRJzOLCYY28yo7nI1jkEFNxk2EsTeGkRkfO1uqT
Q2h4xvzFnIHJpFLQdo29h1MRSUnO/knpzQtOF3+IcQSY/iHZEMFZVB2nI/NPiFZ1CZvglTMj//8F
sLsObXrPfgK3OJ9R4d//3cwZ2BEwEuyex/AUKZVT8Qx0BuKorHyT29DN/SRIIYP6gtKA45qSqw9m
K5KJnNU1ija9JEcladJahVzy44RUEV3Sq0wntoASQIuEdvPMsKaMWVi25d5daEiVH86cMf26n2Nd
hI6OirAUjgKyfJ3OqbaCAQslF8gIeg00SBmVii7tgFiOpfhVuohPHqCDR07oFf9f40JjkE7GQrPT
8kYsJT+BOQ4hokuMy1xt0JF2iThZxsLkTRUKNyjQx6HJAtBor6LmCyS6xXmSKuI6CceG/YWGCV07
mx4J96IR/qLDYSQukYpiLPAgHNZgCLvmsIX0P3R1xznhJV27G3ZqTg3qFd8EXavZG5VufKKav1oO
JbKJiSljEDBldAlLuYJl+nR9IieeFmVtveh8BkYMkxMShCY8d/AR47X1mE4gR7aCuXk7M8ZDOzYs
Y4bgGyWRNKuLR2DsNLIjNvHrT9+kZzRBWXJezO6J0Qi77KKUBAZDMrppilSy1KgzSAK6Ac8zuXZY
FhWLHzkrajCNotWnRw//3Iswomkn5oMOtIJiV7cEpeiW3QpJajTtLwGaaLWChMFk07IOrm0CNDUj
lC9yylKa1qtblfWOoiNU+gWqNYX9nuXhPRC8FX3V/unX724yYMhdgbrmyPu7PBFEtWWYQ5XDPq1I
dZp9AQx+jACd0hfBsbFSSpDhMXA1v9oSnAbsAlfr0cYPQedHx8n4nkVIKg3ufIyYN9r31iCo4uac
DGr5Q/QKSMC/D/r85ecUyOidtrco5By1GoJyZcRvZnuEmwRKSsZVIDXyP0L0c2bK8NYCsURgte2Y
gyJDoAyZXAlIjG7Oc5KZZG/zGaLOdFfq9g88t00zkDRPCk8bHWMc+IDJI++agnKvkBOwRzuYhUAj
b17yFpCzREQenWoG3tWQhDgv7g9htBaO6Btw6mLcwGHhnqJt8rgMnYpHYYFEUM0F36udhXPbyTXc
ZgwhbOWotLUCI9wOrBv9IjuhTjMie9wC/J0ZqE1Jj8ITDJM5Ibt8c2RkUUbjRSZA58kwSwT+AXO1
k0zNLRY0cM9hpaTMbqhAkYJ2MiL+xc4pc/i772sxclR8huEprujCNZ7lrB3UjcyVXSMSldZrCqzr
MVH/H5I+ndR72ZD+jWoIN4RRe6UQlsnsqSETuNuQ5AsyFylENPd3Bvuqr+Te40f0tWJGdul21xHJ
1CtHzfDOLbhG3rk6f29/kswAGUULt0A5sX1vTzAoX9kxO5eZ6H/AGBRKsNsu6nLFrGmuFQRx0Ux6
79igdFQInYl369rTcsUUYzZIKMnlGDFuC4SNB9rrSMqDoeIBGi4tdvOW8ai8kDSiNIZjSk1sYnOI
a9XcRKZ1Cem1h8dOB0vdw27pFt4S2T97SBWqXpllF2sgMzwC7pJnErHt5aCD30tDUU29EqYrUClo
tg0DuQXKwgyxDFAgcMlGwy9DGeYvZ2mDaUEt195lONuEkdlJ09fsaSr7dERVLFymLfS/ehiY0Rqx
Ii2NwqlcB+5YYQtnLhj40QyisHQA36DtkXvAD7nNXP+qHLcg/Y1OJ66dZu9zU4gaT+ChNZ6ikCaF
hHBJaCHuW4b98MJvkPydbH7Uduv+gFkvXMXHgZqfbcfR6QUSXDU5ceL9U982lrQq4QCNrSvgWJsP
6LF3ANKFMUgi1gtpBOY/r+HVYFUUo3VDK8+vYZrDZOZUoPfgqz0oOiRb5jPGcVYtW0s1MtTwklcc
N5383UNjM6xtLP9dJrem4RmjFyyQX6bQ2hUakN4eT8cwWFcJL3gUpO2iiCk1hb9DJ+nDYfqCMsdE
cvfVVsyPoc7iGJJEFd/BY4WZ1WBsFcy638Cp0sFFXxdAtK1uB3ER/+R1/ls16CSZAK+hgOtD1tFY
FSjtNT/BvoDSK8cy67xot49YvLknycXwUs8TF0EJ7TmNUgdji5vjj/uZ81RO0Xr86/Dn6Ktfyw4P
LoHWiSQ/f42KAtbDjiSHgjeXFuy1BLR8ch7VXAGDjBSDjNZe2EFo6qZFixwI7aY4pOLTiAqwIb4c
ZHQuGGoFhsMaRm6/WOPwNeU/viOCbDfYVWeXbxw5+91fcsJLsiYysqGaQ4bzVXF+jL8I2xRqAsg0
J7f2wvMxuX+6GtIPKvhU3hVBdVImVKIa7KQ/WRka2EJboyzJEOfu9WJq0vOozyuOJ24Yv/DwG8ek
Akrl3BHVJwDAuZ7V+4dclqlzzyhzoLcPBskpI6idAwQ4WRTjRpijBY8fCXz3UIDrqK5Skw/qka3j
UePZzDi3lpcNvW4Hoesw1fI409bY5dRF3KGKM84qhBfxAIvVC7uMRqWD3MV8GZ+6DAXdNrprq/Fo
r+R/5/BaaCEia9fqB0CZK4Li2Zx/TTDBxAbBLGxSwBmZ9iCPUhuxB6WI4vRWMxYRcgKqwNv+oOGw
geSkSG52j7c6K0ULYMU+QlvO12r1wjgYgNPQ4iFd4yVWY7yIKOst4LHPaMeJDviu3mGosqHt/mF3
meTtx+ByN6cexYl0NN9WLkQjw9cY9OKZBQXNx7vSTj3tzCtdZiKGMPmJMpGJqwqsM+3ooVf2mMmC
oAeNs64FiMVQQP8yPWwuUZLTJK05QfwRLuerPbpJwT/qDdWNJwYp+7wmnItIpRrBur6wvYg9R/K9
hk1f807uAhSvfsJSLZbAtGiIhzrkgmPCtBDzF30w3ZkddlXkFVXV2YiLzCl5QpAki9ljeJwhSlK6
UsL9vQL5JGRiZx5kfwqwVfDaK1yW7AleEbrsVt//DTx9e6QCBK2MFFsyBmVNTX3qObDSYmagfDfp
kXa/4agvyw3EkvD14O6OI4u5k92wmodq1v9peVxsANySLumFfgXpaL4/QvynDK3A3Nm9Bi6mOMP5
Hqd7IynGLxAINbrGcsn81Cqyw5Pzj54nlZwT21ZTmzO60tLUz+XXc1jR0CwNDGxYoStF/nCNgfT4
lvrhRcN+rTIWOcGTfQbh7XBk3PEJo0WZwNQNb1NYLG9pJpwDVv4CXRzTV0VhPJJsn6hlDduYOJrU
1Bn4IJrOFN7mP9PTUMNdqS+xxGEVJ4g39BEazQAon0n8F/TY49sJ6t2tHXhzX6UG9kuunH2LzVjY
j+MtW+uEPu5dwA93F1/wvMeV3ZvPoLGRgKZ05ZZpOckL3os4MV+MDq5ngq2SpF3RPNsMcNwW2LjV
HQJE82B6QwKsWYIHLDqLIGDrQVIGOVJFP8+KeXHYtqV4MHqxoHBwtBNe0e3+bUmz57bGXWSSO2ql
UijkVaEfpQNJxLFm6URoLzMI+L6uVkZRtqeU3Q5kuVXZJN5rK5btCisNBI3aosVVZzh9JBKo9/y/
le964vzTXH4ydq8MQLf0CHR8+gBxEy/Cp5CC/GnqHo2WJune65+LNAFU/0inG8wYvC8u+S160why
4lO0sv9kgY1fX+EEzRcUkimdmvQ9Lo1YI+wmdZc2LjOGPdWtTVWvha4H0I7Fj8nFOWlRYb43Fx7J
NjsfYSe/sxc0SIX0aBe/+GnqP2u09RYFKJX0AkbEOUautR15alHt75s2aX5nLfInon6xtK0gZUDo
XlNUfwaGUZwkeSPtPpjvOleTIpsErK6TEvj3bvsMMe0jjBTbaPcjb6+e+7sJhuufEHBlMn3o0BME
10R1HF0A3dAeaAtXTtH/yv0ikO879lxk5F9xKgTt3uxpcJuVsgh8YiA8+JStYrukowbOEmrtxu6D
Dq6G2vHuv5kzJMvp9V3Dh44/rlaejIet+iZn07mcNVDUmb3Z2Jznxixd7VU2jyv9jtIDbHEWeCh9
b/MI53a1MkQGQ3Su5S0HxTdjMSrsywejgbzJgP+g2UOq919Fst7s+jTO8XT8nYzWlFmjyRdowv4Y
94ww63+kWLlGoac69homw/pQ+lD9rPMhmpBoiTRoR2FD17pFVNxtnkn/eyMS3thxeGUB/HweD/O4
DWaM3q0XOswL8UnZCekcYAxLrRUNmzCT7yEAf10CuaQgHdVnZQTKN7gtbn5khE+VJ6wwjf5Bn9s8
mfgU++9/OM27IXmaVIXH8V+uU6oZb9NZy1PDgBs0UfBt0xAL7UcVo4ubLkhpyNp1PQTx8GDtmo/D
7gWPE2DXcvI9J+WAmTrBxPsKeCuL9pYA+qJL+fHhGIUFv6i0R3zvh04VHmBoPsLWG58WehXlufnD
3capUhjOSz+wbNUqLQwj323L9vexm18ulsjoXxMkcIJNNNKh6BSuYYJJLN5WQGANHeD+7Bfi9XAq
YhBuLcWIX8pADvLlUFgpbL0FGxrzuzYgbt7Z4wOi/ZzDEVZbyLiupxEh4JbDGbUqkD52VMWRRykC
hwWRSAznd4R8aOjnKk+TM/Q5f1kadWGMU7ifGoLdPJCbbT5doFCPp0upC0XJGgp+aBZ0Jx3DG5pg
TzBHZCptnN+lbpmV2Weplk1f/4Us/P2M8XuScL1Uxh7mmhp3FLb6n36ad6AAR7yIaBfYYrBrfVJG
Tvd/B1vq/djoPmlODuZrMyNz2xSik4ZOBEGerIxvkWiSp+fD9i8ojcUTczkLq9PbBdD9wa5+fAzh
YAf6gIkTL6xcnAOqdSsYCUhYZhQvWOEyLsvACZo7KcF6Yp0qStL4cDTotazpEGWsJg3DIhFSPbeN
UUDFlYnAHCplugMwSd4u8XqRTrW22gW5GQMHMrXp5zZVcR/Et7uM9HripImYym7aCcVoQukzagWs
GE4hxXo8XhMs7yriJJpNh4Ljot2CI3qW8Xw8Rs3hjK3RyBc10lxjnW6wFwMFJ4UOHerhdpMgjNlF
Y1GRxIHCmNMpi9IdkrVFmiVEiq4vJDy1gQIQHU+dvNJ0uqubfGwE92pn85nfpSh0uvTSM7yuaqoZ
UMpWnrJhVaKifAm8D1DwzsI+luu2IvhZnj+vm1ptNkkdATPl8Dc36Ebzzcye7GByhYBQivdTtLod
PTR5kuQJwmygbzdIORODd9R8ucnGD/zTAYdBrXmXUSt8VNjfdzIQsI8WKDrc9Bf5QJyG94s6C/iC
IGScOYsmZuWL1q+iz0ZNMLIAFRBD5V/j3Kz6tSFmzDbrqelNUhWaU48F0u0eZ9c7hdrkFOOAugur
fUDFncvjBKimEkr6XXbbB8pl97nBtG2/dDhfpyIp4EKl65I4DroHqAXaixA/rQD2rAOXBZV5+Y7T
r/3z8l0w40ylwBa0YQUWllCJIo1LwYoHbQKhSmkAVb/FGBZCNaNQilLNeuFzJ34gnqTREuBydbrn
Y+SJU8ImmcvhzQ9EMVclYLSYAmcyu48WHHi9D7KVfvDuvmkYbXW/jbbKodv/Qd/9FkoZGCFBTtS1
Vxcej8lKxXOnW0UsW3UlaEPHvIqh7vjbXMl6jzlwWZSy0TzidtPMUNS7RhogPpHSb+fTTR0IegHY
yEkc+dcmrO9PjvlH3x9olh9aINXJaLLNYEKvtzNS6A5Lng0d9lsj5gt8Oq3CfauFuCziWlrTLNte
9pQLhTwJ5l4gKcYYcEkE0O+3dur3Fo8nqL9ltZcfxnnFU5k4LJI5470hllTgShv7I08XRqq3cbne
SjEjui3EDu+3Cw58zjCVNzjWmqmQl0gPaPXAxNfo03e8Sg0+xkP8myJxkhpOW+qVqiErkjvDHCqW
YqlBA12ihaGp3rHkp3YUPC91CfZnJCXhMH2WC6zc9drK7avF+kQfUIZZHeutOiykvzpOlu2MZOwN
gtH1tDdreESW/gmnt6uF7/+5ppUeyndB3KFC/eA4E801L/CC/84h3aEowBTXjjhZYjQK0BKjkK86
On86elp7HOT+aiJKh+Sh49bR09I0q9OcR1Zn6a5V3nSuE2n1BnWG+iUJNRCe9m/uBRDfcQ4rJP+y
mNPV6E3Yab8WziS6p7qL1Pf0niofDdE3VbOW4NedZIN5Aa4lHQeKGY0ZBLOEMyzJnZzkWDmDrNPG
XEFO986bAPKIHele2YflUoo3M/YbauPj5ep98YsOqxFZ8kYG/CtyhsCC/+d19I9LaJJZyGpJJIEF
l8xciyNznpyH5ytrmw7nG0t+Bukdk3EHg4PoEJ1URShtGGDHSQgeS3axav0O1IVRKEIvIK4Hnzn2
DIHV+ATrzbCQJ2OWxgDi9P8zMLgzcn9yb5OLmXFg2v87SVNAdTMXVvi2xha6240DvS2WsMfa3Aic
pKVxwNZXAgGS6qk5yDFj8DRoHUB/HFrnso/k5F0n4IG8WxP2a6/berWX/NofQNNmGBHv2I2VJXe+
N/f9t2+zF1v0J0rEDPF/1hkfJb2irXWF1N1Uag4j/5xsMZd4cGXdpNfAnl3kfzqtmyD8Ev1wYCP6
fEHJY2kmd1BmZKL7SqnGfQDBWOKYKVOphOdsSYHzNt14hgvc7MRVWj8kGoxVQ9kletmF3OznfsCH
jypgg8uWsBGZB8k5uxTWtE6KZRUSPnvawcFcpcZQb7BN1Wa9+gbINDlrS04bAea8WVDsU6D29fEO
FgxVP4Ig21YPB7Hlxe+P3bRByG0n86LBLhCn4RQ/3fb2jcPFd12d7/2TsX/zBSttAGVlFuKHPZ6R
Ett96toWlV36dw4H4PQ4OX3n+s5OQxowxYbyv010tCeFVpdAGnAETx+80eO7VhdK17cO6xfZQoGh
oN4vvdTSBWtFADpXJfXMrJOG0AUeDHukfOkpTALvcxZMOyV16FLBbZy1P6cf/ZH4+jdqOHKsHwk5
+lW2Rj5H4FIkZI+nFLJ2tL6w5vtpYpQ18c7cUVqojxQpRMZ+AgAF9J8VmxCmm/ofus/NHel8scjo
1sQJxt+L8easThtj+QbiLCmQNXIKAgmFf/ug3ebm58GvdR08YR5OhSYpxU7j42KdP1hfgx89rLOq
LSAK51S8z1S60JjPKA9EIGfJWDa4MyYEfUAhZvJ/duK2II6KTAeaEGsgfYh35//LyT8+owMaa2b8
kYf7GwYBk2oj1YBq9mEAhJW/s1AQu+G6605dcfW7+VDf1a9uOfaVInGNTAFXsYe5GdpHQFmEdX6O
zrbAsemfD55qgqg16n9APH/IKJADWKnycJdHCvEenz8WsecHstYsWzCRBz8dSWuT3M1vvEpDQFX/
fhJdtRHLfCdu2Ki+XNW4PYp99sIxrv9SlraHJ5TeT9A9cTiZwij16Gk/dDRVwRwxSKxCVBw56c6R
SaxrTefMB2qq3iwUjYLc3y5rjVe/ZBk9InppAOhNooQn3lrsesDivejX59hQSwtZH25cdsTuitR3
cDqqxQ2JE97wEaw/mf0jGeFNgYiwgivDc+4avLvZDkNYih0t14eVdFqeXe09pJF7FaA1SMQRlKGS
TM3+0X7x1fjuUcPK9zuinqIXNjpra5+kvns4JB+kDMIIuv0kMVrb0Dx+F+7YIfIOs0rlIUyxSAcF
p88iYHEM6CrM2c52O4koiOqc2SWppx6H5NksUvpiJvryOBjrJfxXc7gbNEPwqN7v9TM0rAzmwCTo
FgYeRD9ATYOylY0hDaUa69ELEodTeBGgALK8PfPsTaMz/o+XiFp9waHU4nO4i+7cdzi6zdhBEla/
HESCHTMqaNlKLZMZ19oSXMzYYYZ/8WR7T6fkdLKKE8ZRBCd8ro7gWQWoj6wnOmrkDBkrqFOsduID
EfwclNF2RzWgvv5MCoyXE9mCP1ayhD6cf6bx6JPtLdUALdIWUxz2U7/eE4awKGXH9Bi/iJetA0fz
wH0NslFxP1LbNNQRyKCMxFF9CV0eCY+yHtYmTZt7w8o2c25xy6EhQ3I5NfT3qTzM2NTAfdWC4y2Z
1GALPp3KQmvRSUUZDFgI7uQsc6xkRRAmNIjNLWzbHMK4p7uxgkJVIqlPkD7qBvu92z0K1DY3tpiu
gCSeP20sonw1XZx35yr2xjhpRcOyF+je0dN5mH/ILvCDlm7DbP/f+gFxHpZFHbJMRG4q2YwpaKw3
7TMyAve1rYal8/sxM4oWt4YDf0sUz3UesMzMCSyIczTFGkP0KXpxE4pidmLhTb7f4dXS+bwvxMlp
sUT4x27wPxXH4RkjCYd4VAPeZLGylQxFtCfRxSAQjHzLo4phpRnmFBBlKjS1IGlA2U23pc/JgruD
ctBnvp1VTk4WfXEO2Cu581P7Z0MGZGDjHYangdA2LVh5IN/100LGMKT3GjsPFbH8c30/qkEQiihV
Yg60fbYl903Sv5Wnia1124xV9bZ9+wjdX+eOgt+7CzHpvbZhLwqme/r8QTm8vs8TB5u1urHDIxTH
hs/+JNv3yrA0+azEgfmnWYcmI6uGUVwtEWbaAR62cUgdD6JeLy0kEYDOwio08eq7BGuJ7FoSTvPf
uUWihqmexKjz9CpcoYMPMeNhZjBaHNmDbLNWQjXCQ+7txCvTGxN4N2vm+SBZbuqG/ajRnVDNfzdW
FWwR3wYXdnlZlY78qx0XiExec1kexN/Q4X/Pt6lSDoJiFt41O3Xu7GMO7Wc0aNpfiHbgbpWyE7Rb
/Z//e8Txqkpnyc0oaWLtwP/QrqCu2g3WijG0gABsU1qFU2GgT4eQNKqvUA+7vzpA8HhgfK/7a5Gj
/2Hd1Ht9QCTtYor0lzz3Yi7Di3ekFrJ5Q292++P4io9EjAO6cU3onPShRm9bOS+/WDt40Pz0TPJP
i8aVKR5hr1s2viH2WvD2OyJbJ+zlELhTxzdaTrMJi6xfP0Zl8uXbkSSmPpTdaFr3UcUbYHXyxnqa
qvA3W6ApM6JRVeRTytFtrE22WDZ0jgJ8e1FZBlE5sSwS5L8qAXcMu1gegj4gbqnxAY3uLqSaDTcX
a9x4fp+BTmn/BMuAArkJtd8W7/46hNb0GkEMXobH7eG/81XPssaR+PzrBD0p2k36tUnU7D4D9TKK
JR2IIm6Yxzp/jGC/o/UgaDDW1Eg6ec1c6hfTdbqv9Fj6Jd+y9So23X6/qvqvc4hcGPl6rOJcXIIY
eFhu2Wl9Hr59REp4M9ttYEToSOwX96caEyo4AOYfQ8lWo5mKgD/+O3Z9oDWT3+r+pUNdfuqjwVsl
Dy8tnkGQCs4YxEbasUwRBvLVqbdxaDxDIofuUJXx2hbHj/40gnmqR7dhO9Wu8QBFmRRw/0ZdDjzt
toyG2EKPQGqHTsKUp9WOcsgsq0Y6A4XDdAKVupmQSF9k69sK4Snv/rktj7x46ztlFvRgYQ9zrKWX
sJhvCSL8rQUDyw8kOhmh9GEdQYiTLXKECZSDs00X3bZLmw7btZjNfcJMDvj6n8sFTIxrfwD72uVG
GYUZHJttQ4QGYHeIwpbyRBAJDJqqInWU/PkFvKeClHLBEVSyIXN3WGnnl2EsO0TRZaChAsu1Um5y
ouXx8Qvh6PrN9a2cNLWFcjHQUs5q+DkYarOwsJQDbF5B1SroiViutIj50ahoWLOmVUexL09uOSOm
H7W5FgmqIIeHA+L7HT6ahuw1qBjUODW3+513sAwKFH/b6RMvU9ruGVNNybWJt1NGWSzBxpBBz6dM
LFmf830Ja2SV8AzWZZarWNmHB0DMI5mrd4npjxjSIZXFE4mXokVsYaw5l64aHO4vFPmXwztELbWQ
86oe70nWUV1ChE1e6VCXizggxvLjn9rXGOTSFyCVe0iJd2tEP+cnVDebIfxmQYEQY+qtUUvziboc
Cteg66gfcSWYcxEU9UMOjZTP8f+IuuUIyhsK8EEqtz7gqVAFPSSTaFgg3L/x7Ez/aH6+0K1bUTyk
mKfrItMYkSoyQV13u3P6sjpSeLggk5V8YXh4NmLBAPNYk9AE8RiZkzqS6dEr6nuX5hu7WBJpVl/A
TfsC+8RW1humF5Hqqahi3rEhy1xBcpibPlDjSGWqsNvnlyTouODYNmoxnt8ArcFbfPhRrlnGu9kw
q9aKVmRGNhajwkn+IPiBgndlf6fjjUj5KNmSaYiFcKgbVj2KnXPlYEn3OLa2IHkXYuSoPTadf/ep
V0v0EbldLVGBQ400Ic8YMnrzs8kSyCAcBQglalTxZAXEnnS30fgcSKAZ+FAa7WV/+EmnOmUuXIoB
za2VxEUQzijfJEQdgdbr/6UZhe0xe0b/Qf4yCrcrG5XaSrZaTxEcLcrc1a6yRRhg5xUVgsE+tgKj
9oEjrkSIGAu07p4L5UoY//r+mtYng/ysR9166dVe102Usm4U5bqpHhw/M5ph5oEqkg1Zz9LkdBKV
Vb+c4FfETFR5ntep3clkti/qFPdgr7w9mS+LQ984Q2lB7izWtzGIhqXn4q6DQBM3W29Tc8Z97vWF
ybELddpF6d51SMKI780Q22+zxTu4JA4Y/apa0GvDJp77y3O0EMv3w4SEEV5gIXO+pkl6hTqSVsOU
mqW+x+C8KlvcsBnnVDIWkapXg+yb+w8dZIsKmCNXenSmcnuFtAUGrfoVI6T973v0NhY+DslWc3tr
Nyyx9funbR5bpsk0b2ytEPykr0WzNDqIplsXTdvXaNr+DwHln33TLpqX/DNbi37zMg/L9bSOeXUb
k+AzSYW27hcTXQpZ2WB50LwMmt1zWQqt+QkejtEll8MalXSL8Atj4+faam5oGNvS4w0NIpFmvfzw
utxiJOvoaWweomDqGF5TgqMfGbOSyJQhNGbVAPY8EEAA4Q22bt+pot6UxkRb7sdbm+lcaxS3y2w4
EIQzBZmhFU8EU9MzJ20etC+JqvdW26jNtX7IfwQUlXUc9GMAAAnBZsoG2CyT8WZL0FvifEB358nI
kEyySr9m2E8Pxy5bzEs/NwEHAJHfUtp8LKqPJ4Yy5qwQgQ2/nwkEMIcyKeOqlrBib7AcPM821V+S
khOBmkAx58IfaF9WaAc7/SkzEGy3K7+jE5O5C7ElcV5mZxJ3VLI2HULzm4iWAnNZnZjmMrpTdw3t
2zMcb/bHgB6ahNrtPOZz28eotX6NfqO4mKNgOpDVFyJFC/qu8pcBLKbcmmTnkuMi6aQ9OXXVMCGC
OtBMSvW72qfMdZypDta32h99l9AnBLnfuyYfCvZe0cMBhIB/M11esfr15VlGe7colng3bWpiQZZL
yVlUcbeWfbtyuTvM39Y32Youhijmk8Hr7tmCYfFfg6xKPrYkg8Xxx1iVmTSDDJFYCGu/V2Mu50x0
hjGRktzxRLrQ39Li29KIZBDKqD+NEhF4AbY7WDjxKhcPkmdwXNiNUbMNMzUcIveuP95tBEf/zhuR
2WF71zdzGPJZJciQGKnJQu39TTPJCNaFvXEJCJ/8CfZH2S74FYe8QxEEJwKr3sZZG+imCMQQj4EZ
N/HpT200B37V71Ef8elx53kC9rRKrYjFF2Z7DnhHDRabYeWyfJ/48/OE31u6+Ckuvjl0gnIPLTA9
gfPP2ifpdpktaSLvrxUrwjwSHl1oy5PhuxAhgNprhCN0ohi1OrrX5QhCoDb4TUQWnkpA2cko00WK
68nOTKfF1aYsR53LIG1v2a5SZZwX7rW12QmdGHudNP1nDdw+17bcMjL3l5londgc3hujjL0afHiO
E3r072W9h0b0fTIF9CBG+sILiYP+Dyzq2AKUV+9jpvvL2N4X96gocaZ0nkxdXy8W92KvdhuNNQWX
mQLHYhPeFZMu/CYZIzo0Ah/4kk82L80c1bv/GgjOJT6ioUCrDLSsG47uMDgT91x1tC9dJ7STR5Gd
Uhyb6xF/A7LsAE6FdywRRHYabvEBUS1+Ey+nfcxqNpc0k2yqYpe9V/rt6qpDbFqvZJ4CrvAraJ5n
O5Z21Egd2ZaIG3NrFgNyPqyKDOtOPkXuQLnPr/+QxVxmQqgcwzRpYkFqjGmaiIzb6K7H8KAw6R0b
EfVlNKK27b4lI65YCnTOcdPqhYEgJvgWBrdyPm/5ohwdOXsZWzzzuyo+BSjKFR6a7kRWEmt46tHC
gtoLzjcH/7Wgo901E6vRFmI2W2FRNjB36qBa4LaSH3leLhRQf6QizgFoIuDQ9JylUKNLMw2QdqRF
AYstrllZvmUQZgry1oA7qR73szWeGAE3Ui1eI2FHbDgwD/EpZDVzxpwTBnRtE0mqq05oFt+kArzH
DT4tlxoSerijes5m9/u9NTqe/w//9ob5kbD5xYCNTzlzmpv4/usTghzNBUGDsrK6SWzpHeCxy5HS
YEq4ZV2QG47EpPa+9m6RkhyKUCQ31h6kC6b7n7VTIBEC7FsJD2euX3BghzTVXhPMoS7IDF9Zh+WK
r/qL2m5Ba1HlY71wR1L7Bw5ACJS7I3Iv2GhF6DMG1WAxhe7LkWxgEmuH1u/8diDQ3AzRZ4HAtVoY
KASyVoP3srUTBBPGWIBHStBc8Kr2Iyh5LWrhVsPSLN35NOA5NaizOHNAf0wTfjJoFwM6Ce0TiuiY
Xshr8dGV+6PcKxcrgwsYgVauqTB29ULBqK+3ce4KjdK6fHuI3/8i6Npe1fMX/XUDFHJq+ox7lkFp
9fvcw0z9o+OLnO30er4kcCtHb7zNj5EuGV7PfaYNal0D46wZC3rtJvH9G2VmBFo2yiFoeHHjIiwb
Vo+MQwIKvLcG2vVUis747Bvd6L4kumqSa8IKWx+4oit1iMwVB6Arii3BcHdAY825oaB5e1M7LDwM
luHfe86SjP6ro57EzJu6wPHodE/dQAFZtmzJwgI8rCo33Gp6VXRRgmTkgqELFaGV2iiR86I/v7Ht
EQmi2TVEDwvgvzHmw6gkspsIoYsLC5YDIrUCpefbcLuxnMNEKd9tp515gqCmEfxsWXYzJZhrzMhh
6epT5xg4QN5PyOk4Capba0Ad0mqAFGK/sUqkDDGyV3FtrKoicfNmukgYLXgY8vHeQW5DPvzk3C0P
5LPb20ZPJifbK4NzKiaYpLfrU0XEXQBx0iyK+y5BkzfXRJ3sjtPKqU0aarkCvUJrQHkEWHz3RsJe
yx1+LXDghMs/Hf9BLHt/e2Sd6Ug7y+2lXN1ot4TrwvGCBBwnkq398HIiDv37CJ0/hdzHaBLqTEUv
j11OQSZ2EZfgNVTvOlkjYm1DKI+BQmLew8pKkoZfEyY8LkMwyovo7a1qb3FG8IP+Bd5XrW1IWlKZ
j4Rq/eqMDWXiyko6iY7Bd5S247UZ6wqGgd2le5LLefQycjCq9LFFxHsTQ4cVx4bJetX+i2GXXR0l
QH+TM1hpI/w3fTyGThubrEr7s0pZiPMQpA85ZJ29saXI15sD37wKLF8eILAZGObsV8kadb4Anz8g
np5ht5odn7QnOMiAdtMCu+dCRz97Tbf4QDGSDsQZHMJu4vIpNu/oWv1r+k+bFkaNaAZ6wQmOeoNc
NvSoSbhMpCKbLMVqeN/yaH/0QKdIIfpT2uxHeMw6CeAOu4I6VoZc8W3/+/d0ylWhdAkpZflJem4L
qvf3I0zzQ73I8+JIg6GnILEkrFWU6ySMDMf6EgrYU1c/wt5WZR/CI+acMKyIx2cFfBrjE1dp4vwl
zsmVwt1EA4HYQceOjjdeQIHHtrWWpbDx4xMNbrn2iBO4UgWnNO43vcTd+oZwBqDKlY+qubhpOL7N
sMW6ffzBJ+1dB6yBi+ZkxIZ4gt3M4HC7klWSdh9EJAwHrQOII1ENuJd/BjrLmFqjErGtcN4IU8AE
zhdyUkji4xWYkJ2kFE70/GCuC241wxK9ONqLYjbfXcDJhVSqpHkfZIgihp5g8vIiXeDV6J8Jv8wE
2wkvq3ZA4xa49Todr00YtCE6q+MuuyL4+tueTqpVty6wHSXw8gU0orpQFJUslHMDwE4bbUL+DXNY
tcUqytMHXgmRosMcXBHoSsR0R+kjUQeSZFFKw89q5csGxYiyJsKIQBwlqW8IPQ7fu1VZkC75FYY9
iHjG3kjkoJZayo+d1duW7Hi0+r/cRkUz9+amGCqkaQe9ItsiU+KGrrMeHpuKM08hwm5N4IDhz06d
r2SjFoxqPdTh1F7ngTQ6+GG0p3NSKeKz0vbAnis5i47RhTZvzKaQedQgB10SlA5eTCtReoaPBIi6
IhWvnVy+OparA/LniEXgug7aZh6FnPKW+2pKBzF6Z5Nh3ahtzC5xVYXG9BJXH0d10n3lA1FWs9Ox
qq2+rQFwEZFzLYiYFhGBlcx8HT9O6z8vWxeH26HH8EMhYG8RJFRQc79A6MfQXmEqepJ2E5SGX4pE
YgY03c9iircTT3pDQbVZ5JUAgz04DszVbt5mhgWQo3ftXcfGIi+VuILoxadHwphtNgVXeQ9x6Dvd
Vzz9Onl8t487rNo8PtYiwdIkGmNI0m7aUI9dVU+c/WMRCvnn+ed9Zfo7+yv3QgNteB8dy2oci6E/
3/78TtU/m+U/5cOYrEUkb+xZK7Tb8cm0JuOdoZm0fzsceN1qmGonIiSbkGL8zrgjAqwK4fC/vujL
HqAZW6qdMx4GWiEx9uTa8O7T4pWam501ZtmYEwxQcHL5kzlVPSGEgK0UZe1wWAOruX+XpcXzgQld
X1H8a1+ZOeBjzlR3VxEeIZRfhvgbpaG5zv840sbB33Un6adVNjLOPLzE1NSB5/c6lYIYNKIKqyia
zxvz8z9kuia+uCHyIPzQYtL0DtHbXG6/DTu5+PgMjN/Tg5MhHnpRzT1ouZYhCtYhQzKKVy/W1N15
GhWu6WFrVKHGmrqQI2n9q2hlmUxAA/Mzb5ExRCCRMd81mMWKKaEGGwxSmcBbCAgIxfThG3KlTIxl
HJDK+kldhGxeG+ewubEc5VWv0VQKZ7K6GR3PcLQPM9iKjAdR9sEf8S5i44jLHd3Y9EVI9QVB/UkI
1higiBu5sKBoAtvPyxrodbZAAL9/kHFOM0Ohk47V2fhVnWH7IZSnWttCc5c5MVWQ2KMXUBEss6P+
ZyEVg2LyZlnjpRKXl+7sJqe33L39kjMfvW44wArERC4JZW24LAx9w7B0L+ZlzSyzVdA7KZmnV/mO
vSEaX2ZCtakVW4Bt/osRPredGTQnduVk/XfDhcmuUGYf6VOBfEuuyILAsyc9teawqdx4Hej+Knnv
Mt4oAWN/n/HN+2Kt0AL7Ll5GLQWKTlRrs1kpl31EggpkcaL+mfQERt3yHtevtiSnIGztgb23sAs5
AtC3UwHM0w3jRTrAI9cFFjpe/k/PB/UtVz9i2m9YK3iemn/VvzMwIPVKU6oW2FxJF6pzpJrZKk7A
HBF5Z2B5CyLKHpolsq/Ycb3v9sLy/tJ/w6164ljj4SU6cnuYAtHfTnoqDgJidZhjMDFkt5H+IY2J
S4V2Te51zg6OXwbr5szsJsehdko8/GPk/L94rEZK/z+sBxXX4Q25rTlAVsFm9BXmp45fvZ1N3tna
Iu38BEIGtJvCISlHJQ4uveFWie77GR2C2Ofd/ipqVM14J8NLibY22O65x1N8ORLS36B9EhdHj6Rv
xk/MHKxx4McLkTI9h9b/zhPvb6Wm5qRgbIf1MVj+r3QK66ePZbrnzeFQ4GdtMhiL2iYcxXDBAJ9z
0PRkZVdAp2sLDeQk3HFeNA1bWYnfEzNdUs5APSM7UE/Iow28JzLGxPUi9o9feDoeKqatAVpgYFzV
BVwftudMkql8NEO+A5wRB40blWzWgzeNCO8jbW8qpvIwy+4NrABtHw5JMgYKMyQPXlyWlLj/T6Mn
nwzwiHcvsyswk9LMD7z2JpmPD/XZiCL3OJSHSki8moCY5xi5TDE1hNLBSjmKGWpwpApu6iDcTMTv
1fNMgBZeDke3m3i+pGlxeOyM4ktjcObSfuX5v5vOE1xdGUBdoPDh0TMkoZQqowbcdqRzeuhpsNB0
qe+ov2nbkQyQ4MJYRkKBRylwwNgwvJ8ED0Sw+SkwYhTVpTaJ9Gx8N5eOMZJHLsvBsgJ+4BZb2VBi
OyqdHl7SlD1AUYuSfdDEOPLVE34ae5yVyj/OVV7dtyjpEvRTnJi+SBW84Fb250QA9I494mD9EI6b
G81gUGJnCteGBFXxP3dihIGsXiI/Em0/N60DX0dzi7qmoNzbugDIuUmDak16drXx+lYo9L6VOKI5
STZHdzYh7zPoSfEsjPHlEsGyOapGeTxXkQKYRHtEHWXtrlGf/077RWPwSd6QW5m6nlhVxqgr7Zco
hHugP/NP5MjxkxyC0+sf18ZCYIOb9T9MR54ZRc6MCCHXW66jqnkXdamfxOn0zTMxJQOp1AmpI3lV
SdeOGiRmrpIZ6J+rnVNyLm5Zeuld9K0Rkg32Yxg68+4YPH+09njYRzsGC56bHdSjT9r/pUPSHD/I
WTKLP+ZlYU0n2i0VI3eIcdspbXlujUSLqPiq2ltxrGQMIDPJaZXwDLEUPZz2/CezLcTasLKBru/s
5DPQVxleuqHn8nTzfD1ODf28s9Hp9BTeJaezO9VxZdOvqdHqhw2nsYveWIBDlrP+shMW1qxHFMPs
+qRb4B8/m67/ZXuTW2+Ybo39RCh85EtSNvMAw5TsVb25qc1Vi20DMJzfsrR9tYiNNr4pOlxbypyz
WEtf3WzBFc4oLaDH3az+/4f1x+07hajZHlo5AHmw4xoUf+VyQqzRoPAH+Uwu+nqRf8CowPgzv7F7
WwOcylb/Leh4hF4An1zK8NTI2oXDim5hCmRU6heKOzmRT0UfU1EOInFn7gGAiT/t+wSWQ8Wcb+qo
45SdHzudoNOY4za8tRDbZLE2gahVJtM7gGkhlcvx34WIzlW6BBCiamrpW9k0KUcI4PRcaT89IUk7
3b/79VjACDOY2utkv9uz3ngpPPKS+xeH2fGTp+fvzYdFTYIacqzGgcaPsaJfCBylKG9/UGauoV8k
51himYKct7MPZmMDQ3zGic8XORYRA+NEj12iIS+zfzT5QSi3Pdwe26mozqby4OStbaW2M/FyCfxM
HCNZu1SZKqJtBIfEkgIfLtaoAMqvzRHfrjjXZXSeUNnoVaGwEQ2TqDmVwe2jISXs+GJUdxLZruVu
g2cl91dq55v6fJCm+6RZCNzcxd0U1bK0pU9nHOlCxDyuz/B+i4jR6dspzMKlrXd94NQOEF9fGO2m
LljxS8D9rm0tn1GmiFDdFTBCqL8O/pOTDKeFu841N/tfnqgUtBQIkOgLC3CkLn6HsjxfHQMog3Fv
1Moh5dAyycmtV39pAHCwhxaBQLKOZJFquxghvHz9r71LHDFq44f3+G9YgeO2NT0pCzw3FV+eQj+t
T1RGxiGMf8hPT5lYIXKb0aOsMWo21alCzefUoMZbOdQvRTBtU34huzZPmWdTPDOEpiHxlv9w1ZBh
rqlWmqEHMzobTLeuZb4KmV5rfPoeQ1V3m6SbYXkbCEkS3o5eh0IONJLZC+fNxP0NqwtIy3l0fDzr
ey/DhCOWicAR+ejeFKmDHqpFaJv6wPKZti6cnEAJTgjeYcGgyyeX9/XzlHPakHObWzP5xbMCq+Z3
h9LH79sjE85vkLP83J3+PDCHiTBz3SCyq2ry1g4fZWYjRkfgjauPP5Al/bxgoP95j6AL/mgyG9nw
QFZrd3Cu8a1N1QM8NqnbFo9pPNykFIKSfUa6qUJj/jXGAG6mMEN+xO536/W2Cacu3h489phHWhZE
142Vjo0f7fxYRJ8TLnEvu9HjJTbU6tPA/4rEFSHswGVcfEs4+c9Vw05LRAf5UiDTTFzDXzdQKoSp
Ugf5endypzvjbZqpg/c5dA9c4neeO4+Ty+XKn3X5K0KxI94J5dypHkMp8liEdxLwPCWpiCGexDXN
j/POOApioXHilKFeyrItI1O9HyQvfYjh7LQCI0TRtvl9ZWf7dIhhADuWGQp7FCDaH5/ZQSOqZSVf
NC4SxlVWDQ2P25X64uBEETsA3LPZPyhzfDHK0Sg4CMcaZK6ulirBCcG3cIbvCjppTRXrMzR3ijPq
YV7Q2IAyct593hU8bDVwx+73cIU+c3uXT9ek/j2VEWJFytXWP78yGv9ktMB1g0GGVCs2Uyanoj3P
v8M90cePb7n/cmL296DKbpStZVvunBVg0XsytYq4+bkzRwvKNj5aCIONy6Dq2kLX3hlHtXEdj4pz
iNw+Xx9nvht+oMN8Ky7oeVDVwpLeuLh7bQ/FEfXlULobcdQVEXoCN3E7g+3mF02IyReQMYfzq8mw
0Im0huMoWq9k2Cw/WMz7WnQ0/1jGyNwmAnySMVamAkW2GeO+Pnr495VtAJwOL/G8RiLtRb972LFN
mxlRdhmyPTRvi0Cm5tqYSGFR04+eME32iVN6Myz58TDDjtBIw0Pju3HFj+y5PygpZLGN6Zp6G4lS
yWDouxr8npsq9nkxYWG3ex52OsL9ZA/rs1fagQr3MdMJoNyOWe5n8cKLKTW8LPvYhRNa2qhXd5mC
GIzDzVsbYgdcFbzO2zFE9R7jl9bS8+qlm1dL7ITz30SgIZtD/JGelWkirp4NesCF/Oxy6QG+cadQ
9lT0gY62/j0ROdhSZ5QtiulBnsMBwTG0E8Su1SRTVBv4L+E8i2gn5g1wyekOZXXaDJGTaw/31gUV
GPVLf+65TUZ8hy18CcV+4hqecS2mKn5p0wNNkitCAINZSH3xskm3mcj8Ba9mUmBVyi+q8k6fg2RY
wRI8iLtjw+A82DMPwvlW3fgHGMQiSaBUnNRw5Ak4wMjEN2yVMeOdMaRvj+nP/Jo63JD8pCEw4t3m
sKQ/5rHB6oGP0VgqiT4foVfYNtP6iikqa2ay0TD4Q+9MTxQ7eYNzBSUI0B/Wbus4xym4ZQcdaKcC
cuX31uYURRXL6FgMo2oKnATdyRue6V5YQYkNuQpFjSYzjNFS6YAbtF2By4it4QjvauRZcwp6MVMr
fuWU86MqraRqW5aKhHnT4bfCwObpUpiC1c+MoOUjiIbDw+owIYVFizB1eFbXj1tM1kA0J5D24tM9
lB4F/PRwKu1YT5LlNxnLQn9Xjoe4/Td2lmriCCwlVYqWQJBm4DdRVtTCf1uXig3yClcse89XxeGo
Tl3Ru2UOGmLc7FApGPntK6toe8gZZqTZEuBeTrmbJgmK2RSbIaYPiFGsUJznWCL+8x3JkrEDpSg+
6WW5yq8fwGFPeHeiXRgRVHIrOyRTDmrVVJSgQBtZIUs0P3gxpV58FZIaf130lkBbiZlHIQqHsiIX
idsh+DJKouSkhMHD8JaZbWDS6JuxUBK0CF0O6dvB+iYqgzzBoY/LN830EbbPLDfTPhS+AJ+IRTxT
81Z6WbTyqKloq1FQW7Yk2/OxCMKJAVKxLQHXyELuW/O85LdQ10KudAl26Y1+K6OGNuu8mvPEp9nL
mz9cXQuiAAmgaH9G99WdI3vlg1y5ch/OReM7y5IBI1Ph8/O78UdETCVJsqbAunBqcH2CMsJ/vyXz
thAkBhXwLYZdEogDXXffkzw8bmTU4zJIMwVEUcr63mh6dcVU0/c6JkeMPxEwoiyd+FLzlXpORpX+
Yg2hnUx6GGEtmgur9yOrSkFAOcuh6fDOJ+l4nZWSmy+l5JjFvyoUC6qweGyHjcLgMhFRgf5Olylp
qfDwBUTzLphNazc+d4sCrBoqyQUejYdu3AVXVqRdCR6xYBZr31+4R55t9HEPO6sCnTGnz+VT2IEy
640XXlZUVl3NYJqcFAcpQaRkum1D/mc0KBx9W1DyMjCo6NlXloFG0IXAUy5TwS/x8pWzdvwFi6iX
lNDymcldaNpJrTpDM5yBQCH9YHmlX8LM6nE9tI96meeRgwEy+x3vzGb1RKkGmYzJtsdILqeA6XFk
1GEpFlX7eyGZH10nwQQGlJXEfDwx/qwPiLboi3XaOZD61Thf30czRes68WxHAr/rjZpkb7+zkUDM
3NX3W8ceSoJB+tqKezXgViOSuvbKTo9CXU3QwFSDSeAAsRSzX1Y83J2wg3qk/Lk49oEXA/7KwsKm
UUQj0aFeF0alJVArOy0ahW5GqDdxYGO78hwSMeecgnuzoJkz9LZHAl+Huoj2GSYzQRSF3/kOeE+d
54d/c1O2/htvww7gHGveK/QnDsJQFQHNYcJqJpntJba4nQdFDg6y0Z5Yr6jBhGsNe4wjCHgHL9w0
JNuR8tXPCGKWn/uT9FgDjNM9vgwbMam84tHkmkPMEs2CcbFwsWr1Ri5QSw3ksVx2Uq+Ag83WKvuV
O1C/eQMoaIKSWqhufFzsF2rSVGEGczzi+371CyT2gQzsw0+xwkbTxtrzGyqw7+pHH3nH29O2XVw/
/BnZe8ymac33pJdjDmRTGes88XRniyotRK8pqYzrnLPx/fr1Vuly5Zg/FZiA+1uZeeAMFPr58giG
pemH/WGQ6DA41xrn4XESm69qbPCZ+ql+JJ1DvJScYgyheVFA6C4TwTxa/KAvJJl08d6FQ46ESCkx
N+pONFsLYwMgmeC7PrN+oYr7eXaKiA6+0J32NhcQlOAVIaz45GwMGPv0Z7sM9dZlqoR8tKnzEcXi
f1HGQ58as/JX6q1wkWIi1YHExO8CKIqMWagmcENCXvI2E7+UGXeZz7MsnSm61wXeXv3tKh47hGbv
S8W5b3UXq0eZDxtCyCMhSsYlZehMrTqLDSYDE22csTmhWBJ+vN2WATk8J5j2V+R88yxpWRIPoe2c
cvZtS+mzAvDe1ld+VRMfkfVVUc0PeFut3Oi3sntsvWoFY8d2ZmsNkIrFnl0xqvO8WGhYSov4fbFX
Hzau+V0HEcux/WzwFOJj8gIWbc5CI09RlNn9OGARDGrK5xD7Ody+YyztjbCrp32KcCNT2uZBJChf
39Uc1BZLjq8pSMxZ+Pyg2fgUAN3Aqvwzss9bvQwwTnJUMNtTwF2TJKWArKRU9rQUeqq5Xwbi/bpW
g9WH+LFu0Ocnaqt1cr0/tn1R8Z6aqyEbJ69ijRj8iBKddNlnXnO47Q5ikMjCWHkhNu9eIhEm/Zr7
0CaX/msjRYXZeQZ5QjAJlBIru1szwMhj76vhb92ohIELAROB6qXTXzx5JOzxMoSda5+dz9YOzHyU
1B9dyJWYNVNP5v+lKO4ibGTxX4CDQifFqZgrWP5hIlJx0HtqAKPUYF374enuObrGM35iyIN4F1X1
faFdpxWGyzf5HoY4t/Hl8NkevJ5gHujPHPY/A69bbJVok2cGAjA0JCfT9UZTNs4kfJVqFXdvAPyv
BQoWt/HCHA15fUqojdZd0d3oKCUw5Gm6J1L+v9dVOnGD/lMqfFx59ZqkGLj5NZ1fj1hs/MC6MngI
NtSy/HvxwAB0ZTJs/Htd0/AlcDapUYeXVaDif2c4xHhpCnR1JFziuh60DxPpIxJmEUpagNn9nTyI
I+waO9cvqISKoIWXU/XuNs6aZ9KEzMbqx/LGTnt895NGXdaLVs0SPyxKabAXA51JR2uHZ8LtYIwP
qrIfH8GgB82JK9/QwGbTzJSTH1y7DcyOSYxqK0U/defdsNzEDXQbzCrlDJEklUQ/x2s3F7a1E1fv
MPnT0DQ09dYPC5PpD5O1B5cY6g/I7TszG2E1a/G2vLAAq1ddYAgoqIIrEJHrqgRob7I4zSA6FemJ
Aac0ofyAQSVZr/WOibDWbSiB3Agl7yDM3V0BsbkpY9omAI1PwgYjubWO5pQCcP0s/NJLaEtxtimF
Xe82RLZdq6ML0aUhtoID7PfRp/6hkrMQYJ2sVYhN7cGt4XVK1RTJTGS+/IeQBpNkEcp6OGpYc/ij
HuOSKWj+mVmQAQN4biJCF37DWL/QBdKposiP6kakqlItNPaqTceVqg5yDFPkKKOUAPuqsrJ1Ldn4
Lg2eHtmBdCTVWfYX8mGFggP8ld3KwuCDdIhnYcav+WvX2vDmMdr1+gvq2poboaRQHOHI24d6LqVD
S7sdjMaeWTobyAzOzCTKH24zgTbPGIPfwKRrcPcrR6RxcLoaq4STKbhFqnMZxm1p2FPSM4cGv76o
+oEyP5goEfE2WeACAbSi9CCNr5FEfAjSkoqeEsvxN2SWw2aPtYj5KkXAc1ty47OM0KHgYRJTYhj6
NnNhhvagoRrmLCz6p1SYt0Q+j+EfFFhuvUjnwLjF0rwB5asJ2f0oQxJKV2UTFBMG/ukwq/eek5os
JlFwkFUOJX1kb5F1JPmNP/R02VMIvjK2UTdgLf6o5GH3x3Hk7Td5psSJjHGrO4y8BmFHAHyv4+eN
7OjJySnY9t/lYFz6VDtKyiXF0+TSHJu+nSFrH3qw3dYJDSG/oOeKjYrob+1xu9mTeujijLhTOUET
eKGkitKGkdFyi7nOd1rsCJWS9TFKYUAp3WYJVh8MZP5nvGyHQueFFLltAB9rfY19KjxWc3VYAXjR
mkY3sJQcwrdKbzg9JbmXTNldwWaroXmxg+jlkbYrmyE+b6YxU9TivOdw9NKVwwP8UZfiGUuIavqb
LwxP7fi4R2Qt3+Um++ik98VHtTvDEQFSu32ZHgmWr7BKiYbuBBaWmsQZQ/8cmk+/Pd3RxFZ+JuAn
tQvWKnzKrnHo64loSRLAA+7994LMg+8iaxjNIcZ/30xLR6h8PjvuntLmayWrGAhXsx5+nqxv+Xud
dI5U2THNeTGr9R4HfHBHxGJ04UH5v/vIywutczaO0MPBajgToNYiP/CqRxVaYOIJB3QfzwXy+67n
HBSRYXSyW57fmfhM9GkdFt+We2KKy8lUBYyrBeOBbzS/Okfq3THjyZdYLt2ZS9z8Aq2Fr9muw7/P
H0jxrRCBU8oiWvcQ3CVkvn2hV+vum17SFBf165cWkxi3xgRsHf1GFEp2NFllbhRtw0N4X9LYihBe
aZDXwBAv++/NC5hpuFIryYOi78TNoEEK6JPlhE6hIWdVmcEDMi7FRPTVr/BSUr2W9G5I33h/EvOd
sJ4IeAZT2CXfNYHx9Anqr8bGWkdZPZC4R3xXOE8/dofNkTxqRbM2AshQ8a/HzPq7L1k2K42BzVjl
qXlFqhwv78bV1ARdfUbx+GXr+NMK4ZfSY0/6kfA/7XqPnyMwj9p5p5A1AOV5dFXf8DQcoDagqht1
2P7oQVlrRlqIDopuDnpF4N1LSWF8C6Ek0d4I4BAyJBLuJqnJwA2Fys/0Irnw31JZkjWdVVusxXpp
3Kp1my5afFeGpq89Eb3r1mjRUomjU/niz8J6GG5VPQZKyxAUGuUaPNGDaoIxsg+Pu4abXlQMqSLa
hkibEWLrhb+JMHirnt1yOl55ZvM9bcan5+fYMks9E6xLdIlyERQ4uXhbJCjmX/TtmEgGMhaPFpcZ
9TdP1KmBb1UYi7WIj+RbTaxdeiZyqHTl9lmzfkYnX3XoHBMpIga2/4UN2FZJlJIHtCddNJamqhFd
SjrS4DdcCUZar1FKhS3KVNK6FAjIlvx4Ej7EqZ6e1067RJ9laxqFZEfrN8fliBJBj14hfAgSkCeE
5kCW9H0XACHAOKcAUTX1Af2tXGLAvYGM8H1VPtOxdrvDzG/S422dCb7BoQ7bu6e3qYpuvAn5mjBj
x4c+Sn2vwVtqkOtwoXoUG0do1Um83L8t6iofVGvGRGKL8yu+RO6GeKeZ9+9sOMd9VZYKSw9SwiX/
Sz8qDXgEJ/OEUr8YlgHQZRlJ9SpWlni1cs/W/WEiBp+XmyE8+Ru3yZtae7BUWVEhN9QrE2+l80Fx
SIQQZjMhYiPEKa0wpcaZuEC9epYaqNYX9y7hLeLCEiKkvfM5Q82/S8JoJm9HFGDtcFsvs8TPMKCU
OHxT/Ggj6HXeIozXyBJCd5AxJor8zMIn2yVxqw9Pc95gexUAQ/BMuq9j9+wBBldbKNwT2XP+i+7A
enYAVy9yr6F4BHdq7AfSGzZ3HcNFAtyDmg4ZyJUI652CgpLK1SB3z5socktDwT+PR2OzICi3pD14
pTHD/EfHN1LnjtPx9uLY0XBRh/ZC8MNkdgV7NfUxLNL+1Kadk2uutIOVNyFdi7+mhCk8IXK/Vmbx
jMnx1ylQMewPTwTQtZH8u5EZnwv1ULmQUq28u5J5A249Z4E/NHeotqzNJP7n1M87/UGXXXEDQ9V9
GUUXAYqn0Br//fYYQygB0TTuT+4CdehiPXq8GveKWtPO+b/s67LHNO2crHOy/5QhKOehjSFRArd0
ivGoXrZ1AG3sHR/zTEZNOk4riGjtzSaZ+u90GeWsUmZbHI8iFvCdawN/rXpnqnDe1BkBtw59p+EI
0XfDSzjxbAjU02POoLVjjmk2vRfAJRBuoGQKQ97/Js89vsSjKwdUZ5O7qmrx0AnTTec1pzptwBVt
hzSG4XWhMuIGVrcnJLAtLO41EykkacSwn3l3Co5fRr3Io7tPYIN2edfwHJCy7C1oOrBDR+rvtCHA
uMqX8J32bT+m840owLrZHfb/de3P2dg/icPSfJJ0QFnoN9MWWzJXnv6WrXsEYXqbHxMDEHVN5nhB
wEL3jWEcwV4SmLQ7rBg+EVQ6NO8Ud0SrizLL+AH9OIq/a/4KH4J+Mu5jsj8nUcDmNtmSRtBAJ+Bg
baKH8p+tk1HUtVdLGiFw6MDuIoXB2c3gSebRvGTzVCRzBQCsQP05sctomCjjCrgihbmrHi939OIi
ZALYgVj27z1oLIAlc3+Xycs7SAKTjgNzOElMo3W3iJjX5IrG37/Gqopbw7Bt6nXV68Lj3e9hqXLd
cCA67jvTm7wmdVka+Kkx4CUq/dDfrh2mbxZagl34lQhhs1TdqENETkD+apQ7/2a11NdYKEX8atlw
xw7dg/mNn8LjUNZPwPddWHuk+jAT5taGST27Y3MMINoQKJVPjqfZLEHImxyviyYnJyGpK8Crn5v5
KjnK3OIyqYumniO0cP6Tntv7+DvTGzPn06ycPyMMzdLw0o/cg53nYSOyKak18msY1yHYr18aKKN6
Cdye74YaeIUPBKuv9mK0Fav/+dZ+E1AmpNVSgBvwc0I68qERH48qH+fpR5ulcH63Y0y3iAzl2jJL
fIl7ePhS3ZKEDc3C0ebZjQHzY+CPUx3zzIM9GNrab2DOV061fiM7ixPNnHZn+4AQl6egyKHGyAdR
hDf3EgaR3sErceaOs3bR4ZvX4dsVDMaQ+0X41zf22EZmF3brU8FHuwQ0elW97XcX86FTzGM+YR4F
Chc1PrTPwsjTG6LLjIYbBniNKKRKwA4ZcV9PZCu8UkmCmFSxq6Hrrthsmhs8keIALY8vbpGlGs4I
Xp9g1LvIQV3f4ulFw7tl5sf54V7Zjfr4XHEE1WYURX7S190UiZMqmgt3ltB0/sd/dPVcQLOFhiPC
4/HzNkCuwZzGdGpPkGSghsYYf+y1XKWiQJlZ3Y/zAsNgskC/d010Vgn8siC6MFxiC2jLqJxPSSGM
Cw39pX0wICXq0p+N9p5plnah1qCJBaG8JlL26CWO5snHh4jr1SIv9Owf4KQi8SvsxXuDfZv8wh5z
HD2+5edQ6g30nHnYAfJ6nxm6zYRfagzMYbRX4pVUazlC4opd/RIWl7c9CtsE+5xcTDhoVQ8Us9I2
/lJFqvnWqod49UwocYqeARX30hlwb1b0s0wlTrCEPWTVE0KbmAO28NUWzXV4SMgoBr4Argn+pnS5
yF1PKvGNCGCb3v8AVEI3k5uoGDcNlM25pqo2tEvGrMpupe6NoM4ZzpcO+680d6HHtSoocfewOGd2
iKoRsS/MWp5FzeO5ZRqc4o32PdvbAL/t9clUpjQjClHl0Ag5iAIO9YTe9uOWFApMHinsx5dse8KP
ElJwpgIDH4ly+5AAimf0ns8KQVRdtEzT7UWIBf92Y0yN94dtg+Henuz9k07KN2BoWFtn1wPauO9M
6k3sUjXXhvAGymT2zArfxFki6ewQZwykEwPXDtxRnygDKmtmiPLD6L7x8Zof8rzdzb9kd0vULhqZ
ugKW5LnCxmOMzsOAQImseuV3IPrcQQA4Yx224fVKpI8MqoJZ8LgD2mPjwbc7SuAYO8P1Y/okeoBe
2QKcGojNp9gVZ2+kHlcICnB79aUx+qf89YLLS8/n412Ok9b0F+dBpmUOszChXLUYQU2KKAwDzcTX
CbmUwXZyrcm2cUipQjfP9UNsGVdRjoRHy1UA6XYAw77hUQXN2+Omu1L9PYqe5pu8HSups+Lxy8cQ
zrK3/vsiIqK6nzltKPgGVGP7YgIcte480arYr/Ei10daIf3tT46mNUE1kViGYWLsy4mUsWk0mejf
JipaILknpUJXrMa4RqfFy3Uowm0f5jbKlUvGS5HQQ1Gmny05nWVjyX1+8XAKJWZzfkEbCD0YEQJP
ESGnjZkg86YIWlLGFDSqOq5wSLT2xoisJLyA8P3fRkf7BYf3UKegAQiSXeOBz2lU2ytEPAw0QugV
DNVPPAUHaxYjGSpqkZgx/10f2hPE/jALLwR6PxhpkoJA/d5Q6BwfHNX86pIXNFYUGUfQ7gYLQyqM
aTmpqH/Taw2rnVi7CJyJ2fhvGBNdYAMDws4nvtLJt5Q9r8810a505LKj7gcOdOSsYIYk2PWIv5VJ
a/sMvkYhOnQIU6szH6+4s+OcKaiysTQMpAA9s88nOgYHVNR2Ml30IiIkCoyPEBpX9qGBHnEwhKXD
AjKfj0lUkfWPCJrgGQZrHqFNvkXpzBia1Jr3MepItY7OZD3XtO1T6WU6b8UsQyGFxUDO7AktViys
yfdUXNivdvBFzGhvaRbLyQ4T3lVBNiZkczN7XxjnrbS3ytdsWHMjIR2kdjkzg2dSvFQuHlMWXmvS
FjCdSRHXlcysl1vNKdzZp7U/HiNTOqOSodO/cKUD8m1CDcs92zBlV1+6R3YU7+bloG/GXVKqBL8q
0SSXg3YAhFLi4iddVWYRls52ICrITzDAD0caEnQyiq0pptIgbhPFKAlMRuPwutq+eXhYMowpzXDl
8ezqQVaUYJVRrklWyGox2Pqb2XRB7HoA7hUCIscfdWTQUQ4k3NrPVPxzYfe/YC3zgqOSNZuyvPap
RuK0dL+h0EDdlL0IWppuq3ZJ/Pbg+6d5/5htDM0DRfF11NkGapaXAI/AH6mU5bMAIrnzIEq5oOh2
WIBgTrcs9o3VSn0/TitY+QBFTMC3K+BTKcI2NfnLuHnMGT1ALg9csgLbRj20o/b3TQXKI4mEDFG4
E4uUk9263po9l4x+cpvF8NGzikd2/mSpy1zZo74CKkR01wtYYoDNGFH9hYPjS9aca+A7a+I2xhbM
Au9aZFTpPcCHWVY+ABeyQ1B+BYnRMD1TFIPhhXj/2de2N+2OHeDnK6ucZIh6fd5yfC06MvLlsk92
5ye142n6N6GffmlI4mpTUDxzlamZfBY3ov87ps1VMwqMrH3Ie/CBYeB6g19DJiK5+GXCN8yNMvUA
ZQGUCmOk1scpZtvMUVlijBgli2sFwBPCAno1Rc1LGFI0fwOHPiXnmCaj7tmW0ulW77WRg6Y/bLOx
pO7cvkHrEbPrOlyXfDkmuZ/yN4zl3DkLPjiXRH2WFj7fLrvAcLWgppmGr4gX1WhePqyd/CH3ZxSD
vfhePmZ+rqmdM3rkZLbKQlFh70FYAytVPgtqVjjHHNKoHccIDF9mifFBFvRW9Wl7VaatBqf1dO2y
IJN+HNDhGjBV0L4s5woJCaXjmhK1PnPMFDit7WzMPiQvIAoyqSxlqpnNyBSJJmqgQcJLeASjJADk
ftSU/44MDhV0c+XmPWp9zJNdEaxU8J5B8/gtAM7fkT5Xm3+aBaCW6L6enFGugH+x3DRw+8G1iNd1
MrzMAWAMBAynlYimRGHQJpY6WxRsp99+UXVmBmj6oPf5+h+nGrSYRoKG87RpUikYDLIEstkS0IX2
OiIsSpGMjoqoheafPpjDD5ig/JuIhrVtb1VOeuibGRXyRdWzIe5/Fj1/aTJ3L6aunk7NhGrHMl9N
HCnkVA6J91Q3OVRQfVrxIBnLUnbRPdT6mZP47MOx3QroCnVstxDsjZTWkzTAzSNRqMjIKzG+6L05
2U6rVTtsV85sVj8Ym72O3rvspvu+VTf9UpTZcJFU2f1W4vSrVKF7OVcFxHpw6V4oSQYVLXoNJtJ2
uYp0vxB8xdya4vE9kebWDvKNqlbmiInTCI1LEESCZBCVi9fkirvT4Caf5ORvWolXNkFETmp7+7SG
rml4r5+Xr9wm7l2tLrnSvmM8jhMkY+ryHE+gcVC1QBQSgVfeX2O8ZC7jUSliq7C7Atxeei2qr1u3
87Dhup1+2b8ZTTWqYzzQdnMLYY/MwK34ju3P1thMAeDBa2MlmWszuHav1l9rYwfQs8zOq6kQMh1t
DLEgA/KBbDzVR+vAcTA+OzSqH145wkvRxyWL2riigl29cla5rbu6oF1CB+la+C8F1ZG+dfPE7tVm
VvimxZBm8tL9gR3WdXy6IQokZBUQRgsZ8H0/FzZaBhYPnX3gPzuJO0boaiCkBslClvV6IIC3WB0f
3LftMAwfvhshjGnEmJpSb/hAywyce+tvJBfTU6ojXzxkAeslotVA1PUjUJYnjxqFiRFOFVjRqhB7
BRRksHNw6q2Uyxj23jdUKJFyE92lao9DzhP4UEjvr1s7JStkVpLbZ0wfvE+eI9bxNRJ2yP0wstgv
xbhmyOYsI9s8nYlrbVNlBEsxn39lVL6IR5vVvZj6vrl5Olz14oKdq8o7fxf5CONcwnNB0/BB+/TW
hxnh+n9HlL+i4z/Q0gKKO4ONHkCJ++L5Nmjqy/Rie+owpW3/laSJRTuO9dETERZpxX5yTAjYx8EO
vzqQ8zrHoI9LVHH7iVVqzy4P3nOhH1xufSnbegstpgXw8qwA6PohHy6Z22S2ZJz305N4IlV7Lkd+
l7VZYPOa2hCPitxxwce07WpBXkefGDXJJgzRaQE7hiHkpuznzav9JlLdBBSCBuxnxe4RbDST1xQ7
8P5R6+576YodIRtCsMzikMsEr2rWzZBl/m+DdcvkDC2wstFSIGyprImnPPUDbpbbcEHH7YV4fAZD
PLxDvd9XzDe5BVqfP2pGnEin4uh2xD7SBGujtjFXNJSs96EfKKLdv3yc95MG1X5pnwB3O27urkvY
id7L/8yM4WkrF27PobGUfsXm6I9T8HH5jMNr7B3TR2FyoIbIldFDAeziL2e9lSy5pa4amFzyiT3K
8/LU1WEYcOO2RhJtfmd7c0A5cQ+HUWxMQ0WQzkrYadyaEbxxpRLMQTs62CINOFUdbe1fmSreKuUu
RCMkWMgmWa/X96vn44/l3Ty/sfQxsCM19GCVt34g+8stCFrsn84bTzLOq2CeespD2Y/eKXNYnTIc
/PTCBV+cu0RUHffSdKC2ewTo9eDjHOmi8NIhzARNAaCgwpsg0XVvHYoB/xxZ0pbwCg5raEKFjbGI
xU1J8R66/B6obud6Dsz35WqbpLFfl0Qb8guxtUBOZHGo2sm0hIgC656c0rTzFT0/YMbl0UWqb88L
WkUpLDJfnEAkoe0xTKU+keIr/BZHJFlRyQ7E0Fwk76VZGDuhyBvAS85P7y0jnAnq1Ib2u4S2MQ7u
XpD0G1N1ypsUPCZfK9Dd8fQG8bG3T31an6It/kpOYKwtDwUmdwxVoTN1h6YtHucGZ+NH5bYqJuU4
2noc9Zky2FmUGNlRKF0k/IBvgSluKNhTjevDBmgPRgAj6CJbnjjNru0AAK2MHsKIbr6S/v/Vd1WA
uN+ZbCJlEdNSJSLK4zoG9lv3Hti7azaL8X9ItK09cK7Rm69foVvuq2XZkAt1RUd7sHTadix2E0g4
rNmQ4b5WqAblPEFMO1YjeQLOJQ4LXtgsRzyJNavAJcduhV0yRP7OlvK9r8wr7rRkzUymG3dudSfn
XA8pfixd5fQ6mUA+n69lZ/NmV+jBA1zLroxK1x2KoYwikWrEnan2BzbXgbDUiApxz748P9t4HMBI
AvoEnhVc0ASLvRC42j7o+jnPx12sTxhU8y3JrwzDQm6ou0yIpaH6yIKMOQlB4hRJvqgaJg61vpbd
/mQgctgtjWi9/W4PvOlalhTRSrJEvfPBnwXCPUCeCKuhHxy3Xdd+jAQNucY0CG9E66rLjm2l46pT
c0++gWeO/1fvp34Vh4Ja92uRWf/Ge797VsACtGGfnOUX5PlAt7TptTrFoZGnwC+TJWXYc+t4lF0X
97fEUK/c1iZMy4bZryZKbHJp3T38L8P+mbJzR/QPKjdLw+nq/DbVuzr9dpbUbKuXGLIxVtscjBUs
7plftCFQM2//jOPmwpBdV736qABd+dRmtkc1ef398ykY/gxo/E3THYKX2wx41K+F+hJmFYo9YA27
AP+CSKCMyiltrPRSdrayCtS9He8y5TXU97i3auRn1X7mIaHcLyScJnA9sp751nDX9+WmLDy2r6Fs
7cmICreQelEeUXumI4fn3fYSsnUSNWyqvo6ffMsXBPfUAvQlza+hOtaY9vz6Ch1dmQ/B52GogG7n
ujZ/40QcBnRu8BU9EkEh9mLBdpP0CqIFFVw/yevhpqjzX2S3Waupn7QpAnh9ZvTmtzQ2yfHywuVS
CbZMkUw90rtx1fT+oa9hF4SvujioCswG+vHTB80/utKAy5nO/9JN6wZ7l/ZZU4OSBGGE+hIa1Xzc
2npxJBMG0LUYlrA6xah5tmFWseI0K1Sd4TH00wX02tLO6NMldpmztFRp7fYouip4Bn6zq0fB4d9g
ODM5xVVMhmraTXiXAb1ZIsct+QmzoCA19yEQhLjPJ1S34fsq1TYgZ+PovqxdS+w5NqG8Uq58zcaz
N/dv6OcEuoH1++JScVLAcR5a4hDnmh89hprKcNbfCBzGnt1IMEwo5+vR/3EwtVKhHOTbynXm3U2s
x9XQpvnj4/yBKefDQwDCInC0X2V5ZRPBdMVLv10E1e8T+rN0VMxlG09EftTx1dLQPWPvv7zWVDxR
c53GN+fbo5mTkEEQ4hdHVw/4wVpVCxdEYzfvIy9hLdOJBziAdhg6U1Loa0jt1QVNAMRtg+TkZ95q
s0KVU/d3806Eq4GCm8mbkZv9fjjX36Gf2DM2yNwJUK25WYCpQAxZCgqMvy+1umDdJpyg59OjngNj
/YdJv/yehvHi62aP3/mX93582sdj/m+bJql1PX+e1khHdna4ItA6VaEr9O+BKvbWfxoUZ+oGLQVA
MfnDpJNZMyBmwtqEiJDEkSd4T7jFFRmVrGnoQZNvbs0AsDpY25/LqzJkZnK+5PwpA5ZYLdXnDZkd
2k8ylugUurdO9aqKsRTdcCikwe88StDxfoBr/MznS5gHZ3XLIZuPmFpAbQw7zbaOlNFkH39yEF+r
Fu9myzmiJiVsifAmeOWOS/pjIrdWMbiAON4CckhNpo5Ux2Zo6l0J6+Ks4ZA3YyV9BH22ON5nWWbs
TDjBMvzbyJX0wGDT2msPChp79DdnHgKKzgalguvNwCC7BnjI/k1U9mB6Igy9+LktDofD1KtP+vJk
n0oe/jEU9LcDq8QYn90S9JNRIFDsHnT8se9RovpEm591AJqAtsSn0NT4R7lsqVC0NP4eOFge7DGN
VOCkU3aN133bEgoWrepifSL0XVLMkWInvNbginzqXmoNWLFLHB3La22ykxi/ypcKkm/EFqvID5kk
u6sGsWqG9NlH6lzo+sQv+0IOWK55FmV++xvKpFLirEJ7+GmLTY0iW/PAJ8Dgam4MFfiwZfk6II6K
5W/rjvIcmh1OkN4vJiz7oaYYuWjMfJToQoXvYWrI+WD/UHoS6fNSQmJEA6pbQ+drIaV8jw3uuy42
ZNwVSCCnhCuLWyYXZC2fNCn5WUOCTB8R01yHkOt/LfxQGcKmO5+Np1xkjZS7dkdXHf9+1KY4NLfz
3PBi8og3pVO/srjSxz9ybHLUO9KXfVru6PGNZXKqfnWcBBrl5dZ8pj9YO0ZmofCiPIeXfapffsvt
5Kmy33RRThRS7SMW6mmaYo+BvShejMIlQsVdviOsE7hw7ZVIQ9kkxCfjMlM3amhLky9mFRhJsHFf
hrhDg1tv1T9eDb5915Cc/veDd+hAy6lKRBsXfRwpN57PUWpIIGzB37w7P3pWlscjIazXymOIQ2dd
qn5Zw8UYdW7/SKTjmy/TtUxmKz2/c5nGa8ASj0EOOCILlhoaWSPcgVAOIQxx644Ib1IAMGfF9Vde
R+n/1/uU3qKgeddbPzt+VgIuyoJDRalv8Uuzgk8rPli8a9ANQ1dDj6h6KIOyhTx9Fw6R4T9d6eDB
ouKH59/9n9iPoiVPzruOoDZ/iKt4FBBlpCXI72DSGjige77Fi+2h+ufLoeh5EyaDE6B3DgsJOIJ3
irYOVNfT35zZRLAbrWK7ev4ou92skqOoJm4Vll94NPrQCPvsNS08PT1IA3jjPsIKNzh4eeFbYc1E
D395fJUpGi8K7vlwHEHZT1LXYIV6gPgIF4L7cixrRx11Bt8wAItKCrr+3XbAkHEk0MxzL3OTfJwr
9Uf48c4KG3EFV4iaN6nI4zxEv2VVsrW+my3/2i3TkzhspqACl29I82bDx71sxx0fjm6o1EcwLDD4
djY/zUHxopZhNPz0DfUo9LWtrxNVUs8rpb5nuNaEYMmkCR9WZ7RWuXAhFm0e9onHkQG/v7aoFXMl
s5uQjmUh6qwQnlloPrwZ+ul5lZZw6orMM8baeMZBp9vL4hL6SeuU6VSBwUpNW0bRYmz2YSKgRFTM
11qLPO49R94iBBHQR0nm06VEJIFLPSEYrarZuqilZ31UNJ0nrOB57s0Xr6qJYcL4CTqBmOsttkMC
HKaC0iYoUt4Hh68wgUKaBj6fJmjEc0rhTrdayFh7ht5/sAA+AHWaN/WTGHbEun5PEcR4GnjUcwPO
J4IOnUr7ctuDpVjVYKQQCl2ocY//uPIgdr1dCrtGfHGu42b4rKjGIu3EqP8STgMzhlWcNYeNoVu/
4iIPqzW7UWy7ZWrM2CZ23BLtMcOLpeq4ZoTwUNhKwlQHluqApWd9EMGBYD8mLUf5yjZ1kI6YSGFZ
vC3m1UiV00nvVIqP3/sic9EfI9gElyZqfONUsaidD3IHjLSVpGwiquhcvzjgsDG//dS/3PMbxkwc
OeGPY7vtYoKiF/ZYkZaLqaZsmtZESc88w3OlYxCMCDsBNKEOIo4WgHB3460yMNGuiGbKBylbfw8q
e8T3w5RwwA2Y9vIQWHtUQTFPLoCsmeltkuxKpfpUVxIAPxJK0o8xXVnsTffoCmPm9CccnzYM9odm
VqlVRZ742RkTMQya5GtBwUc8FLjkwndwzg6mfzGHArWJxP7rrsC6ravdFjdklLtwPPNZVFWlMnSM
PSGRvfaC7pEZ314oOH2K/bnTl2fKhw18v5ECmAnJ9ViAsYKEV0+Esz0uvICO+3MjxOkkuMkYj/lA
ZaChZPflAr/CiuVpHjFSgKxwFJrGEaFdxvrEbLNQ9kMG+Dc1aluwei2hengtAyt1drwqsoslJR6S
a+pepcWbLQFvgcz3+oGqq01FVHHqA1nmDjC4+bvV80GJv0TOiAa2r8OJrjbaZ01hlXhM1atxUGfz
iWgtOcV7CWCRRmXifR/feBbH7Y4YJ0ciN+lBvpWZ9RtwzidXxsRT55hheouzCgBE8LIuZRh7ZhyU
g6SDUhxaydFS7FrUD6vdqugRMhX0MfyJGvBN5Lq01QFUw0IjE5DyZ3q/5VvqWW+iB1xCDFrGEYHU
3Qlq2tBUoeeUJ9UZ/l51lG+J6Bti1xD8XiodtzoAuH02j1Da7xSAUi02vacTkELcBpbDCqQQvAUV
rgWfzzsHPRtILGcxF7+tZP5IBYefX9fhloEqQfLJi0ffHONW1heTN6zh6hHW2trMY24QRTCEbkxS
khzy3bNpN8wcohXnIVfMiAMbWMZXOpUmm5+rlmS2SmX5SeXmvJVH8DHtBbrfV8/CUuPxyH9P9axH
0ASDA6D5tcVMQPy8CzjBHucjc/vlTojuxxx/d+VhX0y/nNML4e6cxMzGSZWIQ04VcVGD6qxPVKxF
ldq6ZVo/DLR/9zmUrY/TvFY8PCSdvymPk0F3egz/nA099zyabOtmUAXiOs9pyNR9qY3hg9GT/naS
QL0erMOJ4Of/4yRKrpQr3N5v7WjeWLlIdy3luwemY5ZVceuj1Jj4Y1WjAr9QB2yInwhkNAJhET0s
Y8rMoYM+Bc80rbJU4WVPT7pBLfp9j6TZfspGyy2L1g+B/9kTHMZHLBI7PCi2BeRYsQb+fmeAib77
sieQq8oTS0ptBLF/HXTYFslRfNL0H9BcyB4MYox9QoumVBQ4BBnHcQ+r5Jit2ZOzTm5Y3JacGgpD
G0hzIUAkZB9sQrRopRaAytPpX0MajKFLSY7nN330+oB6AE/FxJdsgMPPlkGUhTs/2lpkkGJOe48h
UY5zCR6jwjBNq1x0uJT1aAeSOnDZI/hplFCgFjtM4XizYkWb+y2iY1l4maZOL/EKyq2MamyzkNqX
72lEt20wvMg7HrNE/V3VF/VA7pgj8jmK/8aquvR5eW6ktnOdqWXjjOqOxp8T3Svlg1a0tDStx+EG
cLk/UPard61TJt+UCBvCAUfVEVV2Y9+QVTzqSvbFbnKkLmhy3zcC79JWPcTt5hoDx4YXhLot+Gc8
2sOzHmEDCmIbKPwYaEoJoqNUjZqunrIQKDx9CqavkQzSN5Oy0lg2Nx2R3kJtc3WpWGC0gU8OYTKx
ORGew/Ct/RbvG+eDzOEzgQxcXOF4dMwI94zbRhUokqCR5jSdyiurBu4zMmrbEV5c2P5dm4I25MQf
Eofpt0iFQyErCwAM2Po/V5FjfhYFAlClISlHW7RzlI9JSsoq60xO0oqFawjrcmffr/gMfNMYDo1m
nREqjoRxzA9vDvZ6j82L6y9wFE/JePE7GS2urdWdMNXSXpgIyKnae0aaTHBXFdzqpUdeyiFgtKiI
t43+6cC3WeyhosJ4UUc5IACUueWV2QA9ZMgxBDe/U5dpBX6PnwJ/IALUKQjahE/XTKhtRTdG2PAx
ORb94S7N3MNuDuRficpDEwI4Ce3l+8T/kvrKBavluwyr5ruBp93XVMv8OfH+EvIhGrKlo+IB069I
ctNHv9U7Gf8V8iTWF0tBShp5MuZP8geXcok5NdmtG8rjPVrRv/wZNz2JAg6olF1MUWj2jkUR+U8X
Gcj4ndZP6WWL+V1MHBE2XnOr+7pQXqBp35yJVStdyPwW7lLPxaisAEc1xDGQL2y325fJW/8kc3YP
wYpmQw8lDJshTfB2MYwGsIBbOWwBJCerj0+g+F299KO7W1+P5T8d9b6yPoLy1ZQoJj/apajKb8Og
LenVnKtIsY2YoY6Oi3bcmv7KLWYK/+W1aPtbP/0jl0j7AXI1682mIvsAvCzXPuhOHmOoXS3RHdSq
cZ2bylsVwN7jqZO/mBdrmFanvB1KlDFQKECXgrMt/gibpdP7qsIpeYMU0GV93GCBKNAsXvIgTsbY
dhwqf67DfjPZDvVOXsjNhzXSXEbRE1y+MuHRkMum7x5FlsVAFz96aIjH1nOTAO++qZtD3iRQmaDS
eLu4NgcQLZHzVbe9xqsLQEZXAPHzTaYy7qW6OjoPnS4LMcriimoDL5uljpnrKu+nq6BHJf1bN9de
Lo92rnw9+2iJk1sLbqf5YG6KSHWC80hgSv7THhaqEwSXswOYsVp8UMOv/XOrxZGrP32HNt1WPeTc
ULwU5vaz+mB6Kwe8sEqqeAdFGG/FnYxC8y7cySsWTy0gZ6qSCfk91nE+Qe9XQ/n4KLjsT7J2P2cO
nB99s7UBcHQu0Vm09XUpzd7WauxUKZN6L3OXe2inpVyxAQTlQY4MssVJoTIbLoo9ffSrdLTE+46y
URSksOag5VBILx0PUJ1p0dnEyt4wZMSatn4r/7jHLiw/1d3Te3DwuNcEecRiCj80v6qOqdVwppTv
kHobhaw8uJexLhRGJQdOowJqrhV5jnWLoqmmU6ysZYSEkG02O+G/3PmqHtlnWXmqi94NK9Hw1qws
PrHby2WQNUK++2il9Zd1PPVX0pXYzn/AEmFO1E8Pb9nF59YN+xEycRXyL8AL/pNF6B5Orv1b1brl
48cvP66gA2WJIN53+k894mJ/C6FrxZhcVGdkaAtZJDrtO6ZR332pNqd5Ny69i8Tc4kQfQiFdzLY3
vSZTPQnzI406PQuMt7fwTvCwmp2PfuoDuMMQdAiMgH2gFUBBWj6FMbJa9S5Xcepk7vBbeTh235ep
YYENXpYN7k4dsxmrGQMv9TwVXRBHCVoY/VlkAVDmLcMfY7SJMbRmWXzi0fzFvSJjgg8/L+gUhmVK
VRy0ewyoQ00yn8HubwAGJao+8UdJQLkDW0lyKe3M9RlQDyr6UPW25a3S9APRznCFnc7c2oaGaoli
0R1X7kvD+r8GaKtGAMb4wE6P2MkcFr/u1HwEdnRAd6yJXBNDyvvywNtVp4v+0JZXkRmzmKfTI2Hw
XSsZw4HSC8sl6dxc0SWEnLgXZaDGLj7Lb42YOTiKihbSzNSXAKaw6/g0GwJOLc/vCcC7Jsa7aFna
6qucCQEMvBTmujMEv19mtWJW019JLWBWeoXJKM/qBMbIjS6UHtW0zbPD1+cVXY0dwlBdRAme7L++
603blzFeJPPo0WAp1f6Frwelzidosa92MekO4LCNtWnAUVyPQh1oqSp6VNFjqgg8htUGDaw6fKST
O3PV6xkBL/VFkPV2Ww+Rg+bcRvsc897Jf4r95JDvaM+9+HNyIEUudaDt6wJti4dbSE1Z71ftV71q
e59D74rFvGm4uTcg8yOnCnz6fSNOMIdlgJTI5gL1P77EdTxvYwJUhvIbOWWAHtd7ICVJRYJlo2le
A6iy69dwxHlRwvw0jaCf5E6JshOhItnpESSLlvsEOEPkfWGaSAkU/99XRMjRi9O65pvNhwqJq1Zg
nphVavsbKpc+k176h0kanIk/NNr/bXDmgEKO+hnKSYxYsvMlQgwtIEJMZ2EFDHuG7iQO5ZhhIJ96
H2LATMwWN6GoE8xpNOrymDu+2LNcjp2rCv0BxnL6ngq8AEcf3kDQtADVMWgW4CgXF7y3gQINijgq
uuFvEqedrCTrEC37+fiovA/l8I2L/Mi1+uV3fEBiKJuSm8yPc4QkArgghNU9pHFFELoB12p6jthx
+DLvgUiet3+T1O4r+xbRrz8YujTHpK1vcQp0jhHhL6Yhf5CkFRQIKwGmPEDGOVVanpRdJO4lPDiG
nIDl/z5amnRIWixQssgJjvHDzdzBaw0k2hmilqQ5Hnq7ypKt2dOmoCb3H0//wFXwI23UBZ9LaMgL
3R/d08XPolCvK/5Cl1f9EYCEA3vtwMlnmKNhZfkXdNiHvJcSW2oVRQCWYZaKag+aydfWK9F/DPwA
24Ufq8//L0q6j5FyRwOA+iSKroma4SCWC0qPHq57fmnn00VZOFrcMCxWItW9kLPGMyDeBzt6srn9
u1SV1Cgn6dJB2hBGRMoP82u1BMfSGxlxq/sp0EmUOboRHGO5XLzUJLvZ+02VRb0VYQ8Z6yptkykA
Dw2pIK4ZjJBSVHURnKt41EjYYlL24AZL5OJxJpySPBxgkRO3ZA0IweybAMdPxTFlA1G8uyzAzhUl
faqVM03t6+sHL90yAo1FH4Qs2w/c8fSCz5yT7KG1NKOYfsFrzZHV/ecYv+SmOva3U/eXe8NkJeog
ehl370Ed/TYTdUWjCDhCws3yTcg9CwS8GBK7zK5dYGxVyrmHjTmCXDwqss1sne0OXvmh2FwVHPrE
IbhAYTChSeSd7XE6KrAz16geacboPdnhiHEZF9NC7KlHRWB8JpDQrq9JjRhmUKLy9DhYf6WxJ1em
DqhePt7ROAGsZPU/ceBi1DcuLJHldS950Xzft/BlwiHa78dEEP/IlTIcCdH+Y/oz+mzW23v8TAFu
WF6Jx1b7rUY9toFAAR0iF3cf+N76qELus2li79KuVuEnB/d/toe1YQKO00jQJ5zvCuKok5mF7rea
gvQBNmpqu587AIe9t6Tf4ryIWGiGtpW0sJQeXgfQz/llNwlL/ZJzCkrHDe6MeoYhBl+x3dIjZVAP
SeNe4IlJiOml09fQK4OnQRcJJsIQeR5xPrDyC/6ER0KjAiJNf7bn32W0P2EtPbK2PsD0CA4I4hS6
qUMz9yV0oOq8y2XiJVFZrKzbpWAmEtHKFmbi7++R/AdpK2rRZ1Omb57O7IyNpQbzPyglHutsFNEY
pFjH2nWWcikgdyWO6Lcf8EwltosencrNwGmxb8v+0ridUrUcMF+7AAMYwat7Zi0khERL+L2iFqwJ
htGR9CmHNxzwsQxQpWqBDxPt3RUXx4ikr+JbG8x9TEdDUCzmvqQXV1J7NHknkO9oP6BTkiPFiGt0
CU9kgRIUpjcdrCRwbwLIQlcjSARV3JfpANWlkwcm/IAYxjipq1p8s5EUJhvg3praMWkgohnqcput
pePrEQufGmXYpj5JUkJRN6fL/ihz5D4MmKoMJqGp+I70VA1TKw4WTLPZZcy1B8RLQWuUPOnPsz/u
Zrj1LOoDDQhoiKRhT8UOZzyZmldHlh9bfMXk/Ue3NeVD+tE6y7OXmJZuXKDKHj01fooVXURCv0CC
hlRAGRJQ1ydZOGLvIjWdvPX0EZFHjghBVSgvn2hPWpPhe97s3bp8aDtIkEIQbuo76QTMs/9OfHM3
l1DRa9fHdq3RIiuajPnLpiDn+6WkUrEwJ2dIEv5dBE64MMxD+fYiFiwMlaq5upEeik0vjsS1QqlN
k3Vpx7jnFC1if+iSyeUWbWgdHDAQmjWaQU3abzI5zBV+N41/vAQx8yLwi3EaEpdaBNdcFQlplEQo
fRQ/6kCUrXieX+os4yjsmTln+9EaOWeXcL5G8/UGHpunANclkAOTEUT0uxjozazZ6FqJrWEkWhDX
hW0J/KKWoEOEE1AplG6+a6YXnUO37feelG1XqKut3cnvKoVKpI3zgcELXrVj+tlWmc2/dX5/RXwz
gHGIXaKJrs09RrXB91YA7y047RgVAii/KzDFm4I7xkcqap6n9Qh/wy0Q2TPeA6kkCy2VjMCsK2Rq
WwhIiirxF08EMLlpvjHFg1Kp+UAKeb25nOa6VkVMz59R5fBfXbazOGMOb3Ixoer/ylbbuamla52+
6mvROVcjTqIR/3kyLkGLpUKnWNiDZ5uVemh7hZCOh/kWCvLB2H9kU1hbtaqc8NG8cB9nlSWfQ2/w
qDyQbNyyGB7n9gcA7lubcweagTSVh+BZX1ShSA/gh8RLnD5UqKV3qUumw0VaLMtb44vujPGMCDso
qZXXFWQx3ngRzFTiQ9pevu1+vnNIiPG/z+YObN324alnncFODjYoVP9aY3QX+ERLESs3Px+nfE14
cCRwzXLufSpAbCA11l7TswgUx5UnqRwQEpKnM8LGfKZ5ev5qzaxvFShXjGdM94pNC2eOHWYQkz7k
5L/P38nXiPEkJhcGPVj+s+MYqHBaQ9uolFBsSs6rDG8j777HgWSzhRL+Sv5LburdKE1+SUAKJzO3
d16weiqR5GGhjo2ncsJNfSWGeHJI5bWNbc7DaD1cRGUabUMeSG8/sWhfZqUEDCsW9Vz3qe3KnOMA
aZJEvAo+2So9+vXu4wJjw53fXZfSAsWsEBtzrV7p7I7osOkJJBov6qOGS832ixzy9vhA8n5N4GNz
f4T2ieQjuMZ7i782cmcgNjy1+5D1FHZvwtmMssxFRoUSpvUYDPgfgvuz7hmCAJnvm/2L5QpTJX9c
N9fGhdKHUbnbqf0EXe33SCkSt/NAUEVqIHl/yB5a5h7TrdTDkqFRsnEstfFhoqzB0SnAOTn+4Vx2
o8IaT4ILE6OiXKoEeGpFgKAyKOqpkEFuSuzJxVIZ3/yNoAOh5zy8rPOLQK8XsnCsppVy491aRzah
MO0ZcU+GuLsZ4fJ6gs/fJ8waNVKrlOR7sOQ2ktAR64GmP0BV/CAdnejI9pLAIzLAcmuJbUNVcuGP
GyKfDuDole9WzQ+QU+Z7yxeVLmBKkoldIHQi4k7Yjig8YfLlkXdbdJpLVRJooCQOjMIKaUgbq++p
H+IeyHwNduu5B0h1eEftrnHQc6QfbLVtT5K7qmfzgS33bSEuf2gY/EMH2iEuFC84huZnahsxzhZz
03vRhTBccJfgKFKC8loUzT3iA0tB4+jXg1Cr1bhqVHleDyYeHvT4ZvE9y/O9XLJNM0BD5Fkrh5fw
cos4DoWccPIDjd5pP2TZ1t/5o3tuY4LDyx6zStqd3al5bnq6MDfKSYfpF39h8+7YFrlx2G/kSpIu
YP4fmXjcmc2YXRXbBWPbR16/yda+316SMQTxr5X0Xgc3B5sm/STaW2xLD4pSm+7cXtmsRjApkMOn
HWPsvmPhTA1YguQkEZM/t/LiD4ImjimkEVyJ+blYnOTxVY/sPKZ5LxFxZ5XJvzuH8klx4R1dA3lT
dvj3ZURHmncKM4rpTK+pGZXELurNt8KaZdchE3TKHAMjRvXSWrnVnhJMF+cOX3bq1IDnJOGnoIAU
fr41JzlMswIoJDMLDNEqh4EyIxC+/awTJUIR8p42pX2vbXONXr0TeZFRC3aDM+oLlqAaRKaRrGdh
SknZy/odGrcaxU6Livw3fIdoofnfEpXQDaJxjXDOqWrKYW0ruPxRYXK558IRojTtLpUbUJHHXkRz
sGBY7rWtCY+cJbAcLRAOW2qtKA9c/TJn4V7V5y1pdlIzc1anLVvfg5cQ3krF54Xlaxynko6nXZMT
Pp4ZB+0IDIRFmfuYbuYnUJeuOBcNFEXEqQF320dJQ0l512cRldHLvPtHJ/NpcShlpkV8vwLYl5La
fgkt5llnoC+ACG7w5Cg2GQ1a3l277OKRfJ0Y6tPAcr7uTs/iLv1zlmXOW8fjUMJzZpRKXgLOMDcw
2L/4MGseQyl3kj+sk2RAZAMh9aUMNbjlVGFje5ImGt/uY5L32i7yUbsAD2Hhv1hGllPHJpUa1gP7
P1c42D0u7oKcfi5O5s6mGBLryLta6q4g5J8muYsnPazpxnY7HcBEjo0nxC9oMv+pVmSRaBIF8y5d
2doagFhNhvik+gGGrAOKEU0Vv76mREiZT3VPLhHwy3d5hJ2jtbFAAKPKI/uT94APANCo5tSNTNZE
vtDGVcVUBsppnvlpcDuvuFXI7X5Beo3DLrfVS1OuBN8G9Jbg8CBG4vuqKFGPtm8A6qngdemnej0O
ttocPRxtJVlfWhVWQiUkCLj9GORlt9Rab4PsK88wDvHKT/s81ObDwlJDutbG2wF5dS6hA9f5WFGq
zADlvJAGCrpPFrd8EfePACGbd7lA3qeMbxvFaku6Q/sNaQq+jTsF3scCgG0vCcgqak0Re+5goXdb
FW1/WCDiCNqChdDrVHF3h9f7wk1xTTG2BGWuGtE8RMckGYefKtqMHDkOKd9XUIjrnMTJ96+xWKXU
pMyCWZqnP3qGQK34/OotLp47nS/jFQfmnD1j1Upk0F0ur/CP8efGG/tb+WZXt1dnB/wXk+CTCXm/
lERqVSzT+h2TDbm9UYkRlMaoeVUi9bb6dqi18TM3EGMpx4+6PQsghni4bMScthOQjz5hlQvrpO2r
69lcI3u3O65EOhxwvPWff4pjOEE/UPi4mSo5hOzsyEcguv9QMI/xfl4XLi0Ji6+r0FB/0iYqWPF+
rrg0tqZ3nMnPp0vyFTmgdkIl+D5sQaUgS6Jsr7kgaGcgAvlY7nNSGsOOOzrOzJrv7iYi+C1IJeOv
6nJu2lM7Eka1mqI6K9zRScmSr+kloum0zdUO3bNY1w4+i+aM2EtmVhBB9Y4L81H7CjEh1mFvqDt2
VmxJPXKu6L+hNYLpGEfwB1+NUQvBuI2gPFxoHtDwkURUzISpectaJEpjrUSqrfHoCjSNXZ79xwg4
cz4CcROV/58XqK3BLk4fHno15aIdm4nFpOgRTU/Ja0nwVjWP/xvQzYCZLhoa33EZTQWZSZ/mgAAu
/12NdUVOs+6Q/QDI1K9JmEOHFuaZsyx2O3KphorplsxHymc9S5YRjWyR8g2CYk+3KTj+o8yfEdn/
61gg62O9qYCZDemad6f8oTtNmakbf+ifS2goYmCPbwzlP5mD7kLGTzMBsqYsCG9NTlcF3SCb3lvj
P4y5fCXHSuXaI7cH+fsfJxQxoijn0nAbB136m6Qgw/EGyA7Mc8TFL0itdeii/FeHMbZUYkhjxUnp
WYwu3t3n7mawxkY6Av4UW0n3dXrX0vlok3yUJaTR1z1Q38xABdU/Z4OZSKD3lXGepodOrGxuKalm
0KFecZZQT6HR8CdURu/U7Sl3CZQrrTnwtuw6MxXlphNkzwvDNcap/+rPPrt799YPJn5Rds3duOT/
QcZI/JnQhqxkXhhRhV2h9xxn46ogkaJnPgk5Ptw8Ha+XGpOIaUATbqnA1W+aDDBFIBV6RB5FV7t4
EpwEopT9OCGO3GpJlBViQvlSXuQ0JSsmVUIzbF2GV8rtgsz0VzvlH9bnPeEMN7i+b/AB+oEIWz61
WEZWAxwvaAvoWtCssb07u0lwmB/ylKA9OValz+HlPXN284D5j895+EXz9nF8dpNf1glSa0ye43fZ
+x2Ibi/pwbXHQCTiVTD0mZvMhhwQMli6sQk2BvvzfFnN3ug01bigAXQJN3us+AH1Y0i8fmJkYbnl
tPZ3Njzcw6H3Y3f8Iv2eWpoC9d9qi4pLz9HyfdIeBB9xChBgY1XRm4EK4gmVMVbhQxM66X5dP5aF
W6hwMlQ7HdS7pIXx5IShaykDETSR7PT92IYDVi1MBp1Pb4Sh+xcUCCWzDdwcUIUVRhOOqXLf4I+F
cZqgkeim2eHqG9Ci491XIOksHcALwTvAiJLrFOh10ZozAFCepzLINEAR1jXNUxF+z1vOEvA5JR5I
u15Rtfunm0QyEGJul2RFufPi29tWr3SuSSirwN30Quze1XB2i/DVqa2eqZg5z5xEGYc868kReMdr
M1b61/Mrt0e/3Mg8J8Y54BWFEtv9XZkVluZdTTrzJIU6M38plzv+nVDF21nOEddCfxNefj2Xwsve
F+jWPOdh0cvoWtJ2rXAzrP+Y2zoBtXp+UeHR+OYyYBWH/9k7I414805kIoGKOucS8/6WKHrzG3Ez
AMBJRfaBlzrpPLriXisVaTnxF7X2OYvwdAoiR6WMchbxQ26GeWCv8epLv4Kg5Jmeh7vbqiKO6KLX
4kNdMZIf3cKE6+fglxi/LcxP1aQarRV98EcNa7FI+6288bTPOnYJKS8kKfy9neJoUxKEk4trzBPQ
DC/Cqp7+amj78CqurlbLY5QRuqItKo6W6hcYjZeItx/nxaUDsqybEJjllDFfwR6TG8L/Bz5WVBwl
9r7RXOwfC5pYXPGJ8ooRVaaYNMV22nJbvF8akOWBNognIS+uVfVfzfIEw/3HTJrrfcWvaeGtZdfk
GeGbQmsy5vNNJt0p+VdAVYZz2h/WXyNXZxHcY7U0wGCB91i7tA970JSjwjQ1DCGpHeAeT0U+Ed1G
zvyguiQ3QtJG2bV9WAadxzdD65ItzeLwX20qvGo3LgNGL2+4Hznj7NB9/phK8zUNQXEaBsbW9ZyD
8vdOPbgXhi8cI2oZpChO08w7T5equ9ouV7UtpAe+4oUMANIVuPLqZfyB/cwKhgWCgnw+BPHp1qSx
U0AG5jTKeX8d3N65a/KETdpwCbS2vAQ8nkNNHES/Avp6ej+HfvZet+OVAlQP4mo29oXwhIKuWqRI
nVju2o4FiZOEsZD8liL/Qq9s9tOBRTtCxpPcUSB9jjGBvuLUtdEXhOkV7nRoqCb/0yQoZH1e534Z
MSEB1nleYTz/5xDog5070xJmT3pX+4oStXOKHpvWmspDO1g3Gnj8KzL9qicqBdoTVktCeIs25eGh
TQLXHsNfTgVb6W8osxeSjuqni6NkxuJPoUvJPQt9z7uJe0PYkbBkWjf1H+dDNfysYE/ZlQFumpIP
AMaWQh1lPKa2ee8AWccOfb1GDrSyllF1sE0el5FcNs0buTWVLjDf4WGdxscrns7bj5wDZOPuqZMv
9+QvO3c4wpt35ORIzTps37PGiTK7s0vTThx6rRZ44frBQ0INkZRakVSmiVYK2tw1509/L/HW1++b
Y5xLQa2aAgLRdw+LTG3p4vu+ibjqfLoDG+wlmjsdM8eTIi7g7rF47HnNIlksTTzNqTAdh7pI0o4A
FSd+JuxviRHYPDbHkj6NSP4vMaT83m/Rp3RK93ZBlCNGVywXp53VlQVgjW4hHF/Ih+bPVObtJZMR
RXvhpx3uZ43v2Qc4Oitr5KOqyNIMawhnk8f0OdXcbqTkWYJkkSSwDugr+asRHbFB2hSkC6rfDIcX
3GddcEYaDYe2Lna18NBA0nm7dPz3XeJAtsNuC+ogNZdw7TOl8/7vC6Y2MY9MCC5AyMBHSsZQOqa8
33NWaDfYDNcFXkMIHlA9XXoBJXmHjCcXwjoKMX4Gm2iEx3zQw3zfl7Aswl3GFcNLUJPnlpgJaIkE
1WRYk6nasLhh0Oh52KVA3zU2+evFYBU/vaV2R6FuDU1WNSShteDS1hE63vdVd7hUqB87jKlJo2Nq
HWYkGXiGvugkGg+3N+p4i6mCkHv/grChtjB+QK0KwbRyM8cL25Dkv4W6r55d+xloNXTLoliM2f4H
rHufZyZBA2tle6hmHtWiYE24DGxM0kpqtKWe86QEv0rC8uIOAvy+QoBGrW3ndEYtvHtybpksRDDs
8U5GtTFALMuwytv7sBwOsumzo9lDRE/GUzSLC0VLLg5FFw7PgjbALgUP4BtqNFbBkuiNNCaMRaej
euubB4/n3Maf6GhyzswIo2EfzpCkgfIfRol5wVfafObbfWN/3VpNplfViAZ6afwnULrwXRnpEGgw
376/3PTTy9yYkm1xVz6/UtSj1j+Rb9jYxCVQtvtKK1vsECrJeU6/H/wB84bnXKqAEbTSzF2OmfyS
HUhD4RI+yiubzjWwYv7WBDODB0pyZEWEvF8A1tMV7HHVs2HK4FJDZY6k2OQt9bec6+rttVlGxFe/
XtK8pOkVeHk9YeKuO+p5qtsEAxWA5mEJjmEcIPfl/ryMhvVE25FiZ3LUL8uD8QAqVtEK/tId+jKM
dgTx0AyWqUCLatyyaGMbc6EeKw/8FsMMOEz2VfbfLcAfM0ZH458b5lVwg6pYMKuOw/Qld7nPh7/J
R+bz8ZtCyzY01iccf5O+VzGDrdgmB4xcAGM5Uk+XfIBxUylnvTn6q/A2JPcprh4QYMEYOlp/vXfk
tw2/+s63HUgMGiG/nW3LhO24q8HJYVVzBrwI+bewSNYXary2q2hyJ4dFsH1SCAVtrECZHIiFOuun
4Ts/ehf42zxGAFcIJww3xIKWTArKrBkq2t7CQYJtLRsAY0q3AqN/HvNC3+PI4D8fgWteaPor7aIC
vyhvJhdNKaYqA9wSVdq084i3iLRmvmFKBhTTOejaxqk/buxjhR0MJUgWyeFl2BHndJULp1FIt8Vx
V94+dKiSvP19bQaySpT+L+Iu5LZ+QUCJUJMK7PF0xm4PujDAuh3fpiPkcYc8SS0UKM7kdVgk25HR
toJOBnqtrH1lpFzgj6Fb8JWuiWtOMolLInTLMDDn7OOXLNgRbWZeG5+Bg6LYa1GJhKNHxZ3UN0pX
QkXGecodW+xvrZymRDzGTCQMIU2cVRpz96e/GyIln2piXeuUKQYAWDDfJgySzYmRIjLK9jzeCQ6K
uX2WCwuXQUL9ZzBlgEr1klts5qYj3cplfwz41AhuyVtNIil6ujML4TgTlM3VqLztoC4maHB4kEj4
6+Z5WVhpk1gpb3J6jjLf+BFaYYSz/Qf9BKpik86TAiC2fFQQMclm4752keJxArrpFwnPeB3PrCjH
JtywY+Cds8mI99hfd1FANfidp5zWmu9426WfOjcrShPsVsofxZNwsM3Ijbia7/rkvuvfpOh6J7TK
UQalynuZk8Z8OI7Bzd1n45Ui2UjQ6rJSyJDjmpi9kE6cF2cYiLinbnJebu+8QEl9T4luN3qBA7Ww
VeX/NlYSu0Gzk9ufx9rlKaWzk0728F9x3S3g5oibucFRS0gJFzocYuT7ti17iCgJBsz9J8RgD+Mo
EUNdQ1KpibqIFX3o50AIIstb3sbQ5bQsJEZ4VfYyaptFZN9RnMTPwdoVKaw1xwaBewG6IvTprPSy
UR9HzYdQYqA/oKZ/zn+dxaZSSwMGPKbKS0VHi2capCSWgYZvUrVLQh903mgMV/D7/Y4dVuT14Mqf
ihKFIC7SecdJczY6iXgkbzeT8rbdaKpHiHIDYRuh++AdsKBh0rmZ3VpV9Z9Khwenyo6XsASAfYyr
jz8QbEgjSmvZ53uWYwYTCdoM5SkzdXpZPyQx1otbDnPnShgwkhDPIAMaXCFqJRpJAiKbVdfa4UkP
cjhGGjyc/B3Us0aPDt1bXxsy3V/cIza5sNxTHQW2Ek26BjVC/0YntJt0heS9MkNaUWUgm46L+yv7
be93uY5wVG959n4ABzbmvnLiAh32XQ6mgDQ2xVTiJMG6gYm6+BxH58nBPPmporoyfec9UsJRfQgR
D0lXzyNDRjLwxbAUptMz9zjlk6Iv6V33mIrkPMxk1Y+VtsWL1zb7WtYU6rlvp2e1bI69nRYcZXdp
7x1haznSYEepXGYW6bFHAkhPN18Fgv4JxlsyVpjI+x4eQPEAWKYVzLNRnLYfMOGczgaycPWaHscu
JoDLh3RAb/zxOLDQ9a3hmY8z/xWX/3iQCuW7SKj3goAvC86XoVWFSFx4kmrLZmcH2SqTgRZj4aPb
kMGAD8zMhK6wA9tAHvhwCNF6KL64HgV7MF/e03ZvgP2W14jSh9j9PiSg6jABYUwNpS+7y+N/i5sh
IbkjwQYj4Y69pTvvDGK7KKKz/Q1p1DGElEyv5/zBS1PR769PXa0eVcckrOOixEL99hO3FZZEFUKP
yQlULo0yh2WIfAzcIN9Gvb5QvsMy7ruAldrXy42yo7UipfSry1Ub9SZkJMt9atcsgaQuA9ORSgZm
U2njRC8adHwEEmvjEQetQE7HqCyAFvLwyAipyNU5cA87r4GgjQstYNBbfBBLgcC50+mgYxT5nLPB
4Y1cpZh492+8PGoqO1r84P5TNC93InvdShTM6L1BsNZjY48XSFXZmbCTmV5MEtIBKtsgrHcLBxBI
SyItimm6BcrFTQU5WNJIB5GgQJ5RpTsOfEoajWfAk3BhaBAFkCBKXw5CN0ceMutLXGOGZ1DvGQhI
kb+VRx8VWgZCt3mgq1vMjZicakYM9jRpzbec5JJNyQPKXZsNZLGulkqZ7TjO4Uxx26O5zxe5N6vw
i7Xkx494UhoFYig6oP/pizAxSAEeb0L+h+3CJ/nBoUub5BgeWLjBiLXsrdEU86UjKt5Y8K1miwG+
5dvS3x42InqRiCqV1my4EyDpEjJ3yBuZl8gr3y6FRfO0ejz4TN6OyccP6o19oYtJbZwaBE2WcXiV
y0TGdFBhONWS+DfqvKcmT97QbNclcn+JVqtODBBIVFcWJMcmwEt6SgwBBsSOcwXkMwbCLToyHMGu
cP4OW4+xaSJjwAvlX3VJPSgK/094yU//9ahmDqY+8LFdV4491DaEsRNksOnlxZfb6vk9Ag999Ruz
Mr3wB7cnV+xiPJoUtx2EevmSr7RAB1XMuN2fKXS6zBdwMbJARxPAemZYY2l8ODFfDDqfC7Lc2Pad
d+cSEYZS0Y/53CutrQ1sdprxVPvVOcnpgzE0NmAgzklUuoW9RoZ/edZI8wsrR/7i40ciIN65+S9S
huPC/5dBossiFqI38wFJm0NzDe/dCpwY4tVtDqgcyx2FiVvfe9Ggoz9cbOoR42vWO7clhNO/8j5h
GMexPQvq26gRcP2QhHUdBwu38+VGV9IgGJOIN08JtsFVGNCD+kKRMaw6xD8puTKmnkylB97J2+5n
RxPKlA8Aqn0SvWQLi9Mc3MzY3jFdzF7lUFBRasgYOo/4OM2Fn3h2hikM4CLYvH9TAcfsXvdqdfU/
HIR8lRo826tH9tsMKel8SFqVjXf+N0utcAuWWeIGdMXA9wnNdpS636EMgnePbqWHwx1cSdjiScjm
x9SDxbNbwcdZlGnqC+cvFxWWVsTqRTYdZrrUPWpT6DTE8takq9DAvpNenEe9wZ9IbYauUpPm/SAM
mpgiGuPRvvtSdoYE5DZ4gPa4q62onfuN3mE1NX82A16NBFqr4imJUdXWOBuS8AoxXXWs/FNgCZC0
f/p1ah+Bdq5ug28jF318M46IRKbwq1iwnKtyYdq/ZLIi97RXqTL2UoKwO/fKZ+eASijswTPgRC4D
96dbr5X6sKzHklD9qPoNkhQ8MQZgrjAlawocmwM+k4Yia+jFfsfAim6gQ+l1YM3QYSs0Kl+8sntj
X187vNGoHY0q3RY4/nqJyVTqYZczsR2ttyvcrtq23O7nqaM8bAuvslhhO8KFi0PeFP++vBC1CFK7
6I4IWk8UMXWIdBns0dZzOalkXH8DQ33s2T26zyVf4E2VxL9u2jYCOt3SEWSmGlJqAgR4qqEuPtlu
7DXo9sE5vMDY+gAbiy1exo9vE0fMUMiUMuHtt4AiAQCB1lilp+K6eKDUaix03AWcOP7cCA8xbil+
Cl6qW/pB3Y7qKCLek0vSgT5XjFW1l+EKYxy71rHejmcRI1wjd+v5Ytuqri3c1b019nQT96/cq3xZ
zI8nC6QvS1B8Kul1hmpllnWKi25kabiGniBdwPiB26FM926U5lK39J7ge3IHICZ/IjLgH1Sni/i+
aE9+mrPfab6u/3Ett9HhR8qkPOp/XXvP9hyahaDnlq/PVrSBdt/nsmskphZfzwVxJ8J93rS0KIRx
mgRQOJAzHujRQLgWj/d6m9V2cT3FPO3ry+Bgc+S2BYEPNxKSxm3ea6fL7SjLnrXUHZ6KbBZMJeT9
YwPKbMaVSb6XTLah0fUsp4rrCeB5y/dwFlxMwPEvBzoBxeqq7GAQQcKfu/2ZudmSoUURYuKmLjlN
npvXuynBLLQX4hftwNgr9EUiq0IcVbjuCWpY37oN7ttPNr8EVy+f4Eq1JkW5vpIm+Aiu2dukWLXA
EjMc7mcm+v7o/IMKi8jTIAKanqSrtmPuwgNpQ4sPfLI1aHfiIQKVKES7XgS/PXE8VL3S4V0Ag0Vr
vsv5RQPm66ecqrYHHH1LvcXFwIGA1qOmyImQFFU+zJM1hldAjmSNzHLQXxInlFvnmcOcWNqU1m+A
JotkIit6SQ+/ov3nK8tS4b/owoL5WDN7oN5wW3jg+440hf5/I2b5pAEfGUuZ//tL87sb+gqou+f5
MoWOLuNmSfPcgJG6OL9Q3hRKzfGNWEuiTBDv7tpXnT33Boko0/t6P8go6m+AWrYjNpKUHrlDWo6h
lr//EIwd7VNlxA/q2EIvNE856xrGUiMJeF8dpFvAtius8h2TIbwrHRgiJ8tdRVp2rOPf34w+sJyC
qogBvY2bx0KVOm/Q+vxd8NtDPlz9HKvVFLUBI/vx/hnjh9SZK4r9RF/d34sgXbzKlzgsLyuvMpN/
E3nVnBx8fmGJo+5BCMY96p+iK6d2qRXrPcHXLTu4fZcFnXD6mIdQNxpb8PjO7FlY4FmLfGtvB7yT
cZO443TplTBvKp76t0+HSYhCrj7g9KqnNMHX0S/xcEs4uPeSAO/b7ji1k5lyh9Ki2NB8b4LA6zrm
7YnxYsLbN94N7+ZQgq2/HcZ5RLEubv0wRUo3S7yQEfyx7k4Z/C3US1soG+9tRVLnajzdUrR99owJ
+ztdekYSTTT0bcBR8nau+g1MEeatffKzi+M7ydv0PBIO9lzc2CL32/x4eH2ybCyKX+uvTJf3dqXW
ZtQXrri3sqmbGItpdHqzTbN6QnxAHszKrjuxdBRG/BQqAppdaCl+YgSOqXOk4tG2OLecLSVPZA6c
+KijzqiO76G4vPMbzHE3uGF6gcr50OpzRtA//AY1i7Mz2qfsDPy5BumEffwZ/z9SbQhUAS8Sb56d
nwHCR8C6NdsAgBjXcsLqz2tptzrubAwxAoxTcpjuq5MfqgOF/kG8/X9V6pJdNXXF4HxTf2pFF+bl
Wb4MJdr6SKCVDmuzYpCrhFsA6Ykfjd0jQUkYHVa1A72ZqzI9TjaX3UCYS6mFi+Jb2ZTrCNOkdLJ6
jC07Lkwevrv0RYH+FDEdUm6fkHBLtx/x04t3dIm778omSxpi0Cn4EUeQHUTF8ym9H76e0dvOR1bA
8EPsA1bHAAAmDfQpQZ5LG/rT5Omzq2tH1BrHsQf445fnz6p9e5WogTqziS9Vr7Kbqg71SiYADjo1
1VJcjMjz0Bbb3zCxz6YlgSinvMkQz9IMQeR+4LOFxIs1g5zuyrdWYD7fZR9J9VVHaLL5TLdjgRpP
tkwinEXYhWhuE4nnSklw8MHYPM8v2wvf4a5c2WCIjCX5OMpfsuxsRDAwh5+aXOtyJISHCLqaYaCG
+21IedkB/utcRisWt9k2oHQFkq4KUSS113fZC9d/IrF4mipw2vwcdtmwXfUIURDKz9Ni2RUvRWQu
0YE39LF14rrR9Rgwxgnfy3/hswgWmYoifZNz9JI3BUWZiZsR7+LzzwEyxTnVn+PNYVuu2r3YPwmm
pQdbzy/NMkriGmnJiqifoHbOgye8CbH0shEieDPCMxL7yDZp/JoyraFuGLNy+56MhkB4GZd9UFHm
k2FitfPkLPY5l5sJwptc+V2D2m0KDyMevCHYtHx1RnymdDPicPZQjPij/+NL4Ps/0ePTf3daT2+O
3msgNoYhAmH0hWdFroU/EJEz02gdAHJfqfvANaoh9Wg3H7+OaWkGbU6HhdMmCM6SwW9+b85PknLm
FeiNoY8AEOXJnPcrMT/UQzgmTfMBEesmsuKQtpo1Id4kGWV/Vwv0M8tCgJIcIBqB9zxzB2p/4DwP
0CCSQxEOCprIZsrdoOFXkqZCraClNDGGE8piFShEtkEqL0vGkjc5YrqyKF/WSKFxz6uqagWQcBRt
tY1oRsBAPV7ysjl3jdpnn156XnDKOYut+CtKHtSaJkxjyOxFg6jy4Ras3hCOkoQ/wvfneajSnPuK
w6Xc87bFvnLJ/6I17l4EY5oE3Tzv0pXsyHXUvpSncoRLOoguRX8p9SgCTDyhXyTQnYKAjvkiVhUT
WyyTw9fhg6a9LtA1CN7xsDs/Axq+wJ2vEtU+uiBZlURlSOvn9q1gIOm1iqU+fT8TmGXz38Gg0OUQ
5soobMg/Z71bdVrR6+fYEQvA/CTbKKbNINrbLav2IT5HOPe3HVXOZ6m2sgsr2t4c3ryOOu7xHEe8
IflrAPfsK4h+0Ota6051rltsi+ek0Q4G3vWLG0Rx7beVD9cAwgkUPiaG8dlyGZZPusuIegWfOkSt
psXemasXUT8Zms0rDIv8n8FCGoem45edNC36g7/1NdBTaLUFWSxS3JJ+BN3vTh5rnTeRGwZQKRf4
KfAxgc92UkEdy2weCJG9K5wEl3YUMJqf8H078lLrwKoAojkZCC4skPx8Sznb3WxD//ZFw7FQDyyH
WHG5A9losam1Z9F9f7YQB6P90fg+JmuyR85BSYZfJrx5aym5JSYodzHHWEZv9xsVYXVk5FT1MBgA
ud3jG2kdppPvddwjma1p7FbxuGf7NQMEIBzWeay+jT3wq4pn13pIhgHlHBqq64bZXbKGwQ8FQyjz
AjHkfn8uUOv1KMG3eGjhRT+tJs/sPqq4Ri9NOol12XhT/KeSWoXJfa/WdYf7QV3BfGPwuI44PG5X
tWnTmSwrm90E5e7g7fu0eoXujjDnx31hFIaeO31c56TleKKE5x4csXOnT05v9UuYvdyULb0Il1DJ
4QLwoT0keCatCV5Fs+9FLYHErG26Af4XFUnnNL/jskK4QvXCn9QpSKEcheQFS3tbNMp1G/B/9SJV
sW0/RIw6fC9NWYheVw7TsbeqzCCvjCe1AXTkNiUvYRW0Fc3SO1PKqAnr6vvFB96QxIITBd/O2tdE
UKqVcvqYk3uLgWNqZkKHiqAh1YHQmpe5zwON4b3JPRmW7GWk87uXoWqNM2hTPXv9iJ/f2U8Vb9L6
xbFX57LrHXeIyo/06uKPsKvW6LSzcnvZXeG3GO5Muz1QKv4P6CbtIAoIyfoECAdA/0M6D1cCBJYn
eXw4ugZ8wejPZx9i20hwDmMziEhBPrHi10Tvrp4xuwC9oH0391ohlnNavDnFCwxSq9P6iUSH27AF
7beNJFvsUrAqfzIQ9EUyOznZLQMMQ7/cLShUQbd3TaKZXOzSQO/COho4eI+7sfS0TDduhqNNPtLT
OBG5Y9woPtIpbv4HmKjBVmzqfZxSFdM4ZlYDVQikhSm+v0/a409BDlOfg5aEU3LNmk0WKb1kq0bo
kWzrnpoNMfZSTNatnRHcDudHPaEI3YElnE/YqfIKt8ea0VW8XRJKHXrRfzqAn+DVM3S9z3FrejVw
d2NMN/UrOJJafuQSswBBbzkFQ6V6Tgj4zx0nvk00VepJrh9GUzBRQGahxfvAebqv7Si8U6npJFJO
3z3a/86I1PGlt/q9eyN8WNCPFq1N+LiYK6Nq3/ZWilBQhTPP5GzRttnK6ViPwSjlbpqJwmNX3Huc
khziYF8ERgRptvipA+K8TVZJ9KbmuXaXiXocy/giyGJNhEddAvVbBluyVaFndQQ6z9hpLKF22D+3
XBO38QYlOc7J1psuRWDhYl6MWrkKHQVQePI++fZVKyUKiyAKFLuNmiENKJIp8BvAMWmSyz4g5kui
PzENdewMb7tBGJWWMOEcQiUsAEdMK77MKXIEkd1hiNGwJVodCzK2xMtZDj8OYmToeHLaNs3hOVsk
FCS1c+jmdwZnYYCtzrNQAO7sWcTxsnP3J5KAU/ff1nkjCrm6TamGatVnNjH4qBxtjX8vZX3+IclB
F+0zhYEchJ6iMLH++Qb6Ar2F/lfmczqOftRT+Q/VMwtqY8XPDO4UlP5l5bK0auIoTQxZRbEEFaLP
vPlNI5Bm7IoTp0xQFiK9SS0HFKIqv9URUqfTZJCGdCPa+IzncRqGKaZPt8ob5PcKeINHKeylgnSr
i5CFfM1fUo/kJxz3zW67i/gwzkzmtAwdcRq/xyuKY30RL5ChvzfqaChr9W/yWif75LBxTvmHdPag
t2RP4+o8MaABJfXIlj7EU1i4HALTu+adAar7xGxFqbsPPZ0E0v0ET7on2cbmfx5kq0ZOW1COpCTY
qy8xnaovzZ3WPlqDEoTAYao9heIjVIychkCUE6d5YDqCjTvv1SpQLnpwhSG10PDZom63luiceP5X
z02jAzJ9xJEsV+HVnMO8jRMmouW0akmUajtl9dsOeDQgs4GcX+0utesbQvt4A9Aokws8rDbRr7q3
ZYEpI2aVXaMYRu+0jNvRA1Sk+Lqe5JTiGJf0zRNvHQZJP6W5ojwdqfw3rdQXkg/bLJOLc+hYe5kS
Pui3/thEI5wHgJpiFhwfrqYSzMalYBtQk3dyM8RVxzumXlyyVB5aBhI1P4Vr6l3FzWLgIPbNbQq8
hU5V3Dry6lX/4HOOKvgwBr/7YQDP37ZfcInsb865bEcL+7VvTCqbykTr01eavuMm9HQRujUBrpbC
KKzd5MRk0sTrWKGUvlyidHACtDH4Zg6wjdEYsxJQkV13lxxS/9dqfJIVWn5aTOEUfG9yu+QPY38e
e+l9P5O8Dg4bJduIerbkSddrimDrOcoezvQ2Z68heZrte6LrwMMJauxZvZHDZfD4j12i/VF3Jc9w
NXrtN6BNR0SqYxPYt4zj+sotpO8wNfrWMl9hw5v6SDcPZP442ZEynemRkU4PIx87D+HoOcf4ETDD
SsKU+cMWOX/hnhF1h8VcYF2Nz+uULAPWVhekzSB9YaVZXRduUvkYNmcwOrJmPsZcozOHB/BYKus7
M6Vd28JX4iyA72/CqZuQFKakDvuTrXQV9P7p71fZQayPQyDwmCzCCg63xnFrZ/XPy8gAO/L6w0Ti
+hYefRj9N30w0Ll8Lmn8WIxFdhnR+Gg/X3jyRfwQriL/gpwM1RhXRkA2fY6NixwhzM74Ft5yHQ6w
h0LeVCd4KwjT6UJiJWdlnLmcBETo+BRyoc+5KAD5wBNLl0KfXt8IoatrmHqx2kxXvmyoT3VMDjl2
C1yCCWf11b2XNR8xwIsyqIBlrByEwVWITy4jn3n1clxFojUoOAngC3/6LxDOfLleLKuOquAA6iQv
R1jE1RcRvPD3a21UJj/CQsIWEdE+XG2HBlz6n6QIC9rpsv/n7mCZ+OdmsQ8+JNbR9pSGdbhr1b2G
y0V6v2z2jKbyI9uGBOc1Bgibtbd0xbeQYn9JrYKQb7bSBmm9uJVyAnIk4YhVp4nekLqQQPK7He5P
j07vm0N1cWJRP2QPDSAToRU051scpS3qZM1hIcRlhSrPd1emBeyt7rO62Xpw7y8F/a6KVs70D15o
ZSZ3xMxVbB9pLEflVxOI7oI4hCLJdAHdz7Jkb/yWXMDmzgGw7I/i/P3pJ/7XzH192q0FU1CgjDJH
DRrLZZemRopcG2hFj55YfJMi62+Fftaxqoz/BaB4WRCBGcsixCTzDtf+9VPhUJp7H//FsGO293mr
Eq9jBGFcxAZnakeydRyCDyQsTml9DMStLn6tMG+NDiq++zYEOoXgsC9VOv+EPhbPzFlnsl8/zU5O
uNTXv2mofIUxxYMI47wSh9qvc03+XAPpWxK+feUiNLc4ElMlc3hNlMRwGfCIxiUL8WpXRyrrJAzY
FggavO1886lM1JUuYTqayPabPZx5Edka4GaRNBV6HV8DSF1iNhel2R5CsakVXjDL52ySZbM7TPJ7
0S1v3kzS7AL9NuLRFoFqeZOGJ2X53+ETgfG/yeTcRelkyzgbWGBGiiroXGCymLodccyJQcGBljBz
kBXBbaH3AsJvUWnZWt65Y0U7Wp5+9b2XpXwv5EivWMXu1rGjgfQweKlGh8JBQJqi5X/ybPZuHkAs
pmJwRJ7NNikcXx5DpECoYPpbM2FXiPoGWNmuigtFOj57l4EoX1FY6ac66gTacyD9Ym8lz6GDy+GA
Wz8adY8aTf40BPuA6i6BUGpGGac/JEydmzc2sS2iaDwxFm5OThZGMU4td7Sr9fYxnQnuxsS3WKpC
M9GJthT+RtIacdYhJJpKIsVtU2//akxWQe9Yf460T8ymVFJxnDAuA0hdStJmNSnJSJsj4w5hcg/B
cP12gvBkw0yDt4U3nQC27dQQcA3BIOpPBj0kXZgFwYEjdyWHoqX4tbWfy/aHJvEQCu6OVWrHsDjg
xKiQ2xeGbQeumZxxRQ0NFviUqyPxg4de6vr/1exa6JpB52kk97dCVFJWNBY5CGzj17PMk0pbthBQ
l4pDyS5fla6mbIcVxRfuzn924k24McvO4OUkSrL1FMa99KCB5eEF1XVlzu2Hz15NT+P32xhce26K
Imba9+azY1qgxznyLUr5+DZjZ2zKFCN35mJwJiE+Kpm+xwvnRDCgHRFlj2Peuf5PIo83zMZ0ZWTQ
GTQgrBxNBuWpD+NfrBnGMJUbhHyV2OtZgXkMelhPyHd6J836GTnj9zR53tWHKapLHox0FcP0vSWt
PCMEdnjhb30hU3BxkbcHquZ+rGeBk8QX/LdPj8Rt+6Uh0p7j+tFjZHSKS/qi3JjuLHuzW0VNk7pB
+bPMg5czytohq5apFjDWkSad3Mzj3JELDvhCshcKq0d50OshuULD9eT+o1qukHGbdSU0jGLU34V8
gxvzLZp18gbDuNSU38fpeuv/C81lKLcyemWIGYQgiDY9oNgR6E5FE5Zo+r+ItFjZlDA+4Igh8zb8
+5w8D4f5GY1kL4Csy/gamrOyYtVxJVloSK1Pv9tVCZmTRZIVyiSL4YW+5lAiPB8oXUsph0sqZL5s
HF9vSD897bnDRIi5eCgy2vRiic9Vbeg/PO4xzMrKZ686sCgWfQtyEBNgPxrEgU+I3YUxWbNf4E7b
4CZ9PUMVrgjjhGmZ+B5xI/3ve+5+pFpr/0p6eIsMU+gUNo9xONj7yIn9TrVkZhYcP8XEhMZf5f2g
9PmyABEAMepUBRGFgsjKbCLf6B5AwquReAk2G2xU1s0GzmZOMocmPwc335mSeJQjQsLcDo4Lp2hi
ZV2fZmM1UTqy7f0g9WOv+p1emo6/rFsyaayZEX8awAw2+zyE/Ve82LiWbMtB64yyCk+5y6vV48H4
jBJEgC4yqC+I/VTkM/9lwt4lqy8LDlWL+lEkifV2kLMLae0POqQducfNo7kSLbsL+LmtF8xWTPO1
zHl1PJSgDXA4hPAqVl7etGfWFxrObeE818AaOf9hff+y7HxjEb51zHDoLRTwnKpRrhfLp/ckslkk
06uHIeIX7RTRJnbFhLAu1F7+ukntTG/AK54GPmd1NS5BhQDotxgFKjjxIlBz5ZPIrJBG6mIjFKAa
QoNBRR6JIUrKA3KS70Oz7Fl0xyMff3vhiudOEmabolJCqf6gg5BHmlIcZ+hSBelx+ct8yp/RYudA
Ugrc2pr/5KKMUcvtokbwX+dUUjAcr3JkPx/niqcuZ+ydz7vWQRVYEiT09aLUCCpcEEZVSQ5Abve/
hcZ/lHDg5mXvgkkay2vOw3sNfQXH+9yNWFO/u31bQN+DBMCF2ihkT1EBKfAiNpsk2ixE2vrP9jD2
bha+xf7fBmJQaZ9gJ+wiPji0NAMtWT8C6ypfx0eSyul26D1AeYrRL3pUc6Kbkl0arUHjJhG10BJK
V4v4pq60Qm9JjMBcDLFGqHEHU7bogdEdUO5qqpigNick5oPgwAoBD3sRAsT+PeFdkwcRvCqjFLcO
9ABDkcr06NvW6XHR8KLphBXNX5Vqf5Cryqvte4Q9fZhjDGZ6cqAtvpI1Gx+JhNXcjHS00CntbRUM
fZhtfmPQ2Ngeq0BSUH4+lqtodBQQXpLu8eMvPADUud1FL28BDR01QJ6q7K3T3B0AdTCXGCni9Bs+
IiIQtXmmRZx8LZq2F5R1CIGcfBn9ZJ8v+AyqCZmH9j2CB3jEMcWU1atz8wJY9d+4X0atTJv7kLCO
MVMdZniz6YvbAXXYAARGb4aQVN0teUjqQDyoPPOvd7kTmBIPJKR9/uU1T4+3G+8XLgYuqiLgEawB
iMXfOiecEeMi9XyWN9Wa4TsKI+QIkIC/bqR5npvq1fZShA1wj+hrej53EaPXtwoWiUCVmVCSXdnI
14i4WZbJvA/ZcwODLujyRE3DDUqtcztBBrZKJdehppxBYN7AZKCZD/+JnncAVNqAjg+kwQpjs47H
dWulup1I+EwwG4SWzYxFmz1SsbBE1Dd3kxe/pQOZ3gScu27tDrSztSb8YBRYKASuZALxt+0O0ypY
3j8meiRJQ7jHoGdSmK6vc2ZXxeQBgajYZJgUA33nZLQ/Lpr3I4cOoG1XvnPLD1r4xmoqeOaQKYpK
Y7e/3s3pE7nFYtR5m5IAb5dJvvIjGv99nB3eFqbRnWdoBM2thxQmhvLK6Ftz1AEz7N5KdzcSuhlp
XwiXcuFxvQXME13Nj8dqGdpL2vgbD07b0a/TXPe4hzMS1rSAD/WA8zievMENg/nOawc7zkYZfccC
JFYeAiqMUQfa9e9N37uGTSg3q2eFpDFuejWq4wBAptAPYPot5EXJRYrpiKa7vyDfz067iwFMiaFB
7W00S1NOOnrxmLTY7N/wNKWK8HBcgTZ96kUov+7/hRceAre0rwm7kxnb7u6rJyodJ29tUCxeBD8X
0lOu6jOGFWXPKwtsu+Aw6B7zn4sUckxG9A9fEqQKtZ6GUUmrQlM3zvmJ/+A302S1QQGGmYtvil9H
bVi2Kp2VocMLlq1bfp3yEvVEq9fVu6AU65PBiLw32OCZe47axLyNen8ygXpX21QRkZJ9dxnCuoZ5
aDRehJJ1yVFuWBNV0Tm0YMYssMX3ECjgEpr266FJKQq9N33wh+LL6jSpoee93yC8FAdoqUE9o2w6
RvQKvysPzvhLMWGmq4kJ/KP9N4QGutVV4osvqFZ1x15ZgOy9wRj3uYRj1NuttTQQT4w1sPhJ7b66
UlU7oIrfzx+WdifGcRhpYNGcn3/jDKrLq04Abm41VPTJ+ZZIle3pkSAiPrVDWZ7MfZ0RiWJYSWhC
gB5OO++mhHDdlpgDKMWKwiTiql64kBVth/m5tNV3G+1wIpnJ1JkbmN+I31v63dUbJbHovOnuIc3+
WXyU+FT5BNK54X/R6FyEm7th9hRbpsLmCD2kKnce63Syqa28Iz1TfnrjHaUOVod94KB/EbfF9dPa
dpZ30YvjB9IXuovewOKcjPj3yXVm/aaOgL4dI4r389L4ORXhavvGqFjK2nYsuiHJaDBCL48M1GNS
lrIrwttNRl0SKmvpYfEiXVzNYDS9QUUZCFIF3AsIS5Bl3Dek2qY+fgehbMO7HZ9hCne4ea/KlZjB
1Hc4f8zNBuZj/P6N908Pu3KDIYeuFwoI5ErZPB9YUiBd/jNyAT1U++R54pjKSu3L6UdSd1zLHQJx
9dIHq03I1qEAsJ5sM/eDL+Kf1nizGwABwdyPAUGUqVBFdC+kvxuPznK1aJUxjbtAhylS5AM27YKL
ZipY1VyzASP4npkjQZegMiXhrDEr71LbUE/gPysAHPQaEZItCVagFzZcXdYL7YDwzMF7+NtznpLZ
bfTf/Q0yj51Kk40MLcWbCGptaJc28FoA+Zz4EpVU6uKtTj3iTHjVwxsFuRvm0Btli1l/Oz4p2o2t
jbZdS4Txz0Boqk7j/iliiXxQYlQRUrOzqRN8cDKSH5KzpQ/forw9eXHHcaknytgiVQAU/Gm/l5x7
2f7n8q17ijEfkA0PF59P8KV72Yc73uFeC5KgaWMleTnTRtzNNg88psBjs16cQ2gBqhxg2br/C7Rv
wj+KVNfbhdWQh2tuJod0L+LZFG9dH+xyo51RU0P5P7aDcbEq4aC0aZU6wFElDJHo86ibsKpR9hgH
0UK4Yihk1YsLMcLXGjEi8vNHkndtpXL8nWSNa1z4R4AMpPd1dyHgSkJHByREGPSAVL3rypRBQ/fT
FeTk8P6VFsPTZnO4mvNjHogvHhHRKp46nL/52iaUFLTF6LarykNfppnEYhKvDnvqYHCmRJRwWaxN
K81ESpyl8vfC/6pS6g3oyhdUBsWmFsBr/wTKz5zi1Qg+HFS28Ebx99nK7O4Uhr8YbQYE9p6KN7UP
F3EWBrDKOlNWaUulRN+A80vbIVyyaIMykvxoLyDwhWlwLBZw0ax/B3AGlZ3wbGS+IHIJ5pbn/E2u
nawtwjbBD5JYQ7DB4iYmuts56+OFwQ8PzINmyC3+lMnaM65uCDYsmXdnPMmCNNYPLDilzlbcqEW1
F41UJfXZ2uJbMKDZphGYc/0WE4wOGJBN51lAsXFidLXdJYxo4KvEV+U1/ul7cXP/rNwBAEHPHB9Y
qLWToYSQXQuOWtAo6H5r2M2MSUnankScZIVAZheaCgbUY0NGw+EWUfWfQXoapGM3x/q7KVgQShgY
pALC6GpFQT5z7WHIQTA22EXy6/+tEvvjZ7V2xg8LbX6Ot4YU57DshSjjc2+/zPX/YyXQlq810pQ9
6MaSUpCH/TZJFX7qBrljIHD2WJ+PIQIuXuHVArBDnTAUWTnvsZNTIBkyaipu8/rHSDvFmBX3pE7C
wnfGxKaNZu6ThaASM4M05C7+biAau7nCUx5Jn6sMprc4C8f88r7IwQo44/GcuV0FpB9uj+yjw6oj
icmKbE7g7vVga9h9t3b8DOeWBPO713/yCp0KWzfJP/jAB8hx8WuymLTlhxMNWUnEEwrP5GptOmk9
r8qzlSpQSBcfu8rE5uKHoIsM83jsKgsgVZFnQaf1zspIDd7Cg3am2raR8jj7WuYKh7FWcuoPdSIg
9zaZqqDonCFJQBu/bJGFvsIRoJ3EBdv+iJDi9HSBBuyQZwzEuGvNKOePLy9Lt5EvfYWjPPbyyVhy
2O9I6raBKF4D/H5vuvR5FWBbVLBxetsnThh8K5zNsUsMyEDax0Qg/2ZGSGPBb8WRNxJWd2snor95
bS4iIB8STEBDjJkVr2Z7817hE4PIIcc2Dau7QIi4zQzAIX1Dr9gJJSHGimfLl0vkphjcqzjE9oOH
wC7M7neCNbDdtvWWTlxwhsl7mGv/gKxMEnxnwYy1G5TEo7C8NP1UucnXlofj236EqXHBCkENfVjk
dkIvwVjfN7VtFwrDjDeu40lqrzOOmI5d0wICJ2tcipYuB4KXiLFIBrgnbhPOilHulEPGz5zN9xEU
u7gku5f0HkUZNoRaTJESJ1xSsLile9BFx8vxE+ZjkpbHN3EDh6ClzV4vV/oP3Nl8rpTXNjKC7UIm
IWSsLshikzbnhwNutAMQU3iD/qax0qOG8XzvQp8OnIunDHXqLwerkbys1UmEatJBCGGP2xaxCzV9
ee4Zw/t+kxriqXKQus2rDxEZuoJUioGwqwJN9K0ssXGplIvDIJSPHJk+hz25wwjCNvlHEjy+E85B
eZJPHC1TQJ7FwAmDmkQdb+nIR2au0wIZDY4cRKdzCTNqIZwK3T42PZauOy5c+Cv0uJEXSlURKn24
Pz9zrVwmvA6VUyxOcgWbO7l8D6T8COpe5vedSkJOZD4WrM04RdTZiWJN3tUzDqMFoAjjNG2YQEqy
f/ocHFW3FSSFDf8ukTrBIAnrAo3iZJ3SIpqdXMKiaQie04GsO65p5oStaOo2rT+eDCoRMA5oyzdT
HJVrrDUHA+fMx1qm2Obmq0w48tUu4R1rcY+x+YFtYd7ptGRrLePZfAvBbIJRiIWfIqgEnjTVbtCt
0VRNwkMFCAY46Q20JHYtxqkN/oDPybnUZ+LxEyrc6VemGbsWsML/h9JWLBg/gBG1f+OFvjjw37Uv
H4FjjfT2OfJr+Mc3sQbnqkYPjdm1zmY8fnd6x0Epbh1wNndNo7AYdCUOVBv+kmoNu6H2IXy9Njm3
h06pRKV1zpTF7i8AdpFhK2bRYeLUcKbmnL3NG3tfq1PtSRbmY469HlttDVANXeGKm1+/xjTMkWio
IvD8HKXCMDsLamCT1zC2rdi7+YAIxgJCyHA5mxMRR+1Uw8sCEfR05dh3nViBLRbAPhIPfDL7+qkj
ko/LtE/WVgWdO6ZH3BYcxCVpDRoVN+JRu0bpbgd+gUiJnbGLz+wdYQjt5xf98VvoKfvddsp3ZHa9
CAdSkTi9Lxk3HbwTv7ePyWxph0VCbRpII9jBf2V4qFTvByK+xptAWnsaRuoPQrog8kDdBvtcITRv
Y1LwrIM/rPbP/cQzRO4KHM5VzeY+CQVDzs06liEuqqXMEPVss22ir/NVNiug3ZaZaJ8WTvRxOiaz
MGh2uIkDssY2Wz2hjlt8nFQyQ1/5ALVk3PTmWM+mBMZUE7Ts+8/XlV0K2k+XhYh9AmmQg7fZhfwy
L5wgA3HZH2eMke2wqDUugUMiduIdocm2iWMlb9FSl8W3vMRPgHOQiADLYVSkmzZBolNsnwP6RUfG
xlj38GOt3vspnnp7xe3hlAIiQHQsYNdeEE+FDSxYoeGEcMGq4k/9LhzCh7JhHoQLXY/b4UzqMhw1
oD5Ana8MkBJu7j1kAdJRsH+5nlBjjQn0xtp7afvZ1meqBGkacOn+P0laJg2cBJmv1hrBIg6kEWKH
gY2ncx1XrH1OpWtsIXUrZNNO6lZJjmaqgYQqcqJ8ZqkyoG8RnECS2rzAtjdw2Dobjfuhx+K7cwDj
sSgDHf4YTc2Jfx0shhXR4isRiQMvdwz042sjWgqFxveK5KCpaG3egMTD0wybxsTErZ7Mefi+HNo2
WyfV+ej/xhhoiqoEv7gX+OiPIRdVemSqCx0uylYOAUYqPi0YF7MKbUzd/K1w05+R8AUHu0zignjx
6moWawhqRMCYEM8g6J8eoowWj2u2dA/GTnYedAuVSqS+xW1IfIvYUvDx1eLC1l7sXqi+zYgl0ux+
eBwgfa8BoVdP99JGA+1YhD6/SO2NVdydyuUjUZGj4WL/cpWaKq+mmtlQJ8GbSEhmN9IRp1seBAu8
Zk/Wm6e/pH3gMnnuiTuvWDDkpj2ks3Sa+k1gMgMFWMbkH1xVF1TqJFK9LsNWqBeRqpkcXF1gskF7
tGGdkRmTI7LvE3l+jk7DqtQ7XfcXuYMMwU/1hbv9Gp7Yp95qWfh0F2TKLHS9h7b430tQF+bdQ3qI
g+R5e3BSVMOM32t8hqaj3FPMHEOJJDTzxGZKjD0rKgyZ25xwM9Ic+BtFVP0k521YjcwuIEJNQz/m
g3XmpIqaoFGXz6m2pyQQSIoviPJOhoPemIs4ZhxxXtldHuXvozy3Zbs0ByPbzB/tdufcmpVHTdOT
RF3LtFa3Z8VOtiQnseW1ESZ4c0/pAf4CiA5idZ9AxuQtLW9xN+M+oDzoBWurswInS7RmneFL66Cy
6CSZMmfTB2CKoDCVEt4m/ye0njQojKWfBRta+THQ2vikoTPe5mE2TRQPXvyaIbikA5/qPvqzb5r1
fdxidbu7d+ZrcrL03Euy+JLWiPJmfMCP5N0GcARjeH+sB7oTRlQAXhNUji7ENjG/z69UTCDWAYuC
12vynlGlt8+PGKHe/6RjMTe9ncqtX4+Nbr+VCfZJjXenbzKL2aZtC+vULNeF23dBBtOJa6rrhSEU
LZil8MAS4W/j42mzpzAyHyUqHdyzuaLgonSMKDfx67A97NT/nbA1WJE+hu1j/ian4e6SyGRRgDzu
QKXjXJoySaezu9yToXWRJ9F+HiZbTWxkfNGJWoehuwwXL+5xM4ecFj729MLfskwrhv9lVmqk8zrc
zDO8gAmDZz6YTBF9LH7UrFaz+bYKO85jdvTFPUn/IaGM/5wzL0u42FiDQ+Q/i86r1iWRbaTjEnxg
81wAPbz9LwqbYBoHAQtRbnK4+Mw2w46S9jUUH39aq9zlLbECjgRF+LKMK/yhfUBsJH1sL+eD+7ab
UfUAKWzi9WbgwVvkAGKMNeBpLbnX573aob+DTFH4BXEtPIJTH4eKxOXVydADMt/awUi5DGmQCQUk
QggZyMcIhKN+st6If3WYzE12JQEdxkDNxG3Nbwoj3s1+25MSQpi0BF/eOnrb3zBjvgw1pOxg5tdk
fAwtEklCyrn/7sWZgTwId08Lbfzqoa5ZJX6AzWo4wt3FWYdbYsV+KeCbD23KQVxbAg77cLgvPqX1
zFvoap98A6/SmL4Bw/d8F9gpufQoJpOogfwN+WPL4LuhHmO8BKLme5N9JT6VIz75kpFA/THLViVW
hCowQcgXTQK1ina5nNEfZy8BY1m2fsrqzgcGZ7ATYZYjbualE29qtp+GffnOznyBs7rMw5Q4IjXM
dK2PhRQpL+JoWGoL+N+ZCmU2k0Dx5CcUYAVgho4aDnjiFr4bV4gaoEnSyrZ1Zf1e3e7bECOGHmT9
pWptBFu0lNnNwuxJ/c9muT1RF9UOicDKyedlb6tPCwDh6zWdY04zq8ZUU1JVz72Qrzq7BimvuXf+
6aFgXIwxHKEtAPfo2GEQown9tGLoDTrvL8/hMgJLGRDj4k+kl31NR6q0mlme2F+ICJVpvXIdM4Ny
73NWLlIjpEpmb7oSxa5MwwF/6jfOlQ1VTGe29nuwzEx0QCTX3muvQad21mpnIG1j9lRFF75oDL85
RH6DqjkNp2MQXtT58RmukdEpR/Ne0FwVKw+cVvCIsMbAXm7UNE8TKNqMhw6dgUa6PmA8sOt3y9mi
sVBCOiB/2mitasZ8jtpTQg0yv3pRpqwohppNP93sUcTySgDN5aSc2flYbUHJhXynQwNDXh9Db6vA
8a9yTpqx/bpZfugmXIgGmnCswERly4zdkAIuBKlxoI1FUyOKI6ADFZIuIyuTbSXTxbqwRjmD4Ouw
n3rq6V2DLUcSqYevB4obpKWr3KbHvqJPtavEvMOoHZgW2ZeoZtnqKeZtmkP4a6bgPBDTL/KbonDQ
o/1btCQvu7d3lvl5roDJRKEisCw88cjMMkQMgz1jpm7sgBrb8os9Mf3IF6abwT/6mD2I8reydR25
A1AeYZprofphfc/EwCw+Vmy9fDUPOfr/IHymyRnRrGjXSvuzF2azgJ/lYGgXaxuBQteJBCLBa7ma
rYeJ7N33VI+DtmaJxbK4KFDwInWgV2SI0AZTZaNF5L+CPIzjq8vSC5KMTh53rMyybyR6wfiYez8F
ZEkIuFyBVlteDuX8uHWqygUD/OSk6uB8miq4yYMsvBb2/m5obWUfDU2W7Oy4pWK/IdYFFuXaGksX
Dq3+InamHFrVteoHTncvTZ+FifPASPAxk4eBPsLLfdH3wn0NJbuO36YbWU5QkDIrxYmbAbVicNQ2
oAU08Gx68V7BYpFO0doS8J2o/k/cBv1d1PKSxsu4j4x72TxW3mMIZLnZ1ilhudz7GS7f5JAALMVU
6y4WeRYDk0JZNnL6AWA58I/SFQRhodCpiaeP1crs1LFJBDgDxhaQd+hmOYDkRVYJVwyaZON+jghL
XeLmQHhpq0hq1N/dr1TVe8Oe6a464/RUuZcyMBymOrRf9khT5ogfs4acgC7dSRorVLK0DNvDuoZ6
+g5Zrhz+Q8y3Eu4AvYYpUWD7U3+fDK6wHF3pcemCKg0Ck3IG1jfaAeiQhLhy/IZ1gFN+P8VF0OSk
JKdUM4ITWxfKYDO0nPeWSrHoBuW10JSBKQjMF8/vtUTgN2TaYd2IaQxSiD75jkDXdFF6Mn27Q3ap
k1IrxEa/BR++rugqCDgIe0Y1HhmOFvKl0ia9xoECrQrLzVF8//lr3NALOuYIsNd83Fak/HyQd/73
mx3IOZ45oExiWFcpd9Z8oVM71um0qAw88xgWcEAM/8zROa9wopCIfx+bC4cJJAlQ1cTUqQaq8pNp
htnI+aJz8rzUO1AiE3vnw0bGX3Fu3qZgwWUUaLH/Xk+B0OriswKzSeP2Z0SiurkqCDZ+9unpDusC
IJvXrtb3Mo+hDMgkKGZGIX/DbnUY+OYyi4AsKYWDui3s20S6p4Ocq+xX/Pe8bCDwBt4J/BFYzLEw
dAqBimaNS3vfOQWGgq76yomxpRWXbsv2Jk8WjYyMCavdEa16HYLeCip7Axf0ZOB+eYzICn5o4L1V
h9RX2TzckqML4WCp0pxB9o2t11g9jNTeCLOe0bIZw23P0yOKh2pLUksOLGdDjE0HtbU3/qc7s2mh
QTHaRJQsXHCX3+Sj4tjx5xD5kqfbyCGCiOwPWQV1G/bCZMnEKoN+23Ycs/VgUfryp9tCsMxXAaru
Yy+By3V5omEmjcwJXZn6DDcPEZ2v2QwLdYfq+U2LL7gDM60hYZLlQHEnOKPytViODvq1DjsuFRBX
KSMQwTZACnCR2xnDv2CXnbQCcI0LFMGfiTqjIa/ofyJu/qoCuPUrcj7eQT5Tjl/yHb11glAW5xRJ
rjuX985igYfS4yH8GDK1wtEOLsDTTOM/rnAQcjQkpOHa51QwVytzm0oZ20yf22A+R97xUUvBU37j
verZWaTW4gvdemyeJVbvDImQtJgXtosvtDWs1wZ12bTXvOYi6ixLVlz82JwFsdk1xxq3aeRVuLf9
vPTi1vFpnTbK4kosjI2NkkpjVbRNdXSOmDosp6zFhKmA7HOwtyxEtJEdAGL2czjPgbSDjZEKebZe
2VxJSWI+odTjGUnK10PdU6U+sKaLrA5b8l8W2AOUbUTPD43zDsHvVOOw3O29Iv7zHU2+dOdYAWoc
0Y0xBAO2se5y1W+TU3VakB2ajDw5R2Li1bCkDrD1O6w5st3tx4CtoH5Si4p9WfWoLR7RzRESJRmi
uZR74+xRSfXeBSzqSTBVKw8fpxUkOHb6lzyHAWhAlzYo5ajcfqJ6F57StPcy2R4WD1l6wROAg7+H
9DEFcrg/YQ7JdlVl/yHTvjx5wICy/1S3U21s4ztVJXh2PrA8WEiYdV7sokJYWqilnK9UMlrF9IJH
Le8hgpQAO0IfgnefUF/Oz5EZPBacTfWt+o0UZp7QpksSVEPC5Be0Biqwan4imoyLi/I/ysDstSt8
dNag+bMGFvmKwbtKWuh/2iysxZ+OCQT7TB0FC786mKT92H2qRSOgEP/FK4IbsZG2xthKhPl0PSX7
XWgf7bFmVdivoHfixQfeCgDMb8IFXCDaHSwneqLT4bzlI4d+xGCqCOuRY22HDywRtuaZGmHgBHO/
j6rQxDI65cQHSpOcxyfcMVRHMcdoYRFEpxVW4z9tavqmMTpQUd9simYqfc3+RTZutw2GJyyrozDd
K6Wjd5N0IfQCszfWnzQKKAcLE0NmoWL5oAFMMjBOPIBiCg/LHUVDOkY3KlrLpSGsD7cTVh4XfbCV
wnHcJkdTHK86dSdfP544jHwsQGlJAF0BaFDSQJAyzyHbzUmaSCLSGOBsJgsHAgZPzteM+Pp06xxD
ThjA6HVouOdpSfNY7YBROXUhBghgPzXplBp0oCCI2nvAuKajPSt09Q0ZrD9RBGhb/5k93u0RX/vS
A/LPOXWdRwSrOgHp1mySfoBzsgNeYaatvyQtvQc0KxdZkw2vRbN/BQJBlXwPG9AR87dATOMCEyZ2
PQCSMCWO64zySMbWbBSnvBJgckxB9Sq7mqHnuNGlCgoU8M4Lx3EB5wD/FaOEsLeDd4Yz1hldsLaR
kLRXulHoF8vMv3SU4dgnVfY80tZYT0Qol3Fgs95l4QBhMkKfuUHrSuy4Ni1XSrS+pJEcGpCtAnWz
XUCaoVgCoFqGPaVgGQsYfR+f+y/7P+njnypFAPRgZrKqxYPuMAGtknMyXgDjNCUCgp1E9WWO+R1t
I8zq8CfkvjjKjyRC3ANpJBX8cnn4G7qi/2Soeublcx1/7yLhev11eOMfGGOYKWBdVHDqV0HVB75y
0HhhlsL8VRb8+bOLjHHiLNmBD2Jq1SAys65KJE9H139cwFODmgssydWQ3g7qAMVNvYWK5eMx8Ego
49yr8PsuhdBjDJhJJRzeEYzYT7moEZSyJWTAD0ZooFvhuNis7n9LWQOC6UWbv/Jea2PhfBV8ns7/
SmEmclrnLLVh6SuetpQkKe4RMFtGoRaBph15Y/64XPO5jTy9/qnIbH20EBVA0/q4tRFz2S0+CHrc
k9JRovY5U/lh9R2ijmq/SSSNX5sSLwcInGh5R6gQ0ymbmYNMV1JPoZtIzvhuXXJ9KdQtZF6wnJhH
jIH0wxIlDRwulJjhOhjnYoaVlBF+CuXBfgko7NsEwaCzCaOKGgPlnrcEoRG3bU/HgWAa6JfxQbhE
WjhjZD0cT6MwiCKOUMbAFYWwxdhgbhvQrjXG99CqJnaBPlXsyp3lnkuMho4GNocOHpL1SItZ0dqY
KkM45vW9oogHwt/tkLUHMPF6ESvw1fuTG3erHsJmUOaTKCrsi4dICGNbzlaxafPgeAt2jRPA6bGO
+tnxMrcCUdpGiiWYrYdbwufD3GMnCWU8GxjwXmN6H2MP+95T5W0u0/crJJRcO8AtDLThmGukSrX+
U77BoFr76j+O+b+AQ4oY0XXAJGqGgol4oiVwhEGSUq6uf9IWRJJ9y9uUhcx3ILtFWtDPWtZn8bbi
adDDx5I34I49pUghzJLjevM7GTM0cueW6sVXG7KTqL/jc4RAm+YYmWt5m1lFND5EVDRlRtGwqCYE
y4fVWuVSI8g44Y++va7QXtTflUImJil0B7R9VdSNN5y8QfbUs6eWsS3lG4qyhnXutW1peTGdEGBQ
MLVrusZS1NsYpryfSZTVzvxyowgC9gTArBdP6CdBoTpKQyD1Qt7/9CElM8ifdpTVVPF9xnnYKSch
/hAiw9GoCI1DfnHTSAptKTQbzPQ2wdzzzsjbzvG6eLhavrKyH9eW+4nWli6yNI0E48Z6hVK1Xceb
RQR9dcIZ+0+m3zHoi31MpTsNyXCZgFFwOPOhKWVbvnsr1MbaeorXCojQLkGa2ywAuDCysiZg6oo9
shjf5sANaE0g5N04u5Qe1anV9DMqbpfH0iSRf+9KjYkLDbOQQYcA0LaGl2OZx8HdawuTuG0pm/f8
rvGsGW37jEG6GwiCVhK1I/5InZcNWUJoY/XC/CrMx1tT1pqYsOFek11P7oLH6W5SMf0N6VARwKb0
1VXDx8bUl5GBz5BoFQrYWbkLgkmZcsnMxyh1BPfd0eBt31Mmh09Yl2oNtY2Bm+tymHRHiKzxmHMX
1dqcOChQ1inkxiLd4VsUpPL8yS12blAhuVzhG0Be5yCntMp2YSa6cngP7ki2T892kkC1jdiXtfKb
AWk25sAyUWedjc73j6bzFJSFFuOhNIzFCkMl+uoVAML8404ayBv70fTVkqZu97m4zAKHmBfz0S5S
d0VoIx8Mly6AMF2bZimZ9BImk+6LlS4n6ixTt3n27XB+fyZeULb1yS837A1Ifj9Cpp71/Ff/IvDU
tCQu5HFYQROnTKzMzETYH2xPQDMZcMY7+I5sGPQX+rAn3aPC3HoOQFFXz1SfUWKIP3Il1AONJbtR
sM6p+Ksk8aKzeG4bJOZ6G6126hVDw88BXrVR1eBNIKDgxMPdT35DdITPEFuXGg1pBCpHYmA+iWtN
Z2WWQfaFsXGWn/FtuzRSw3gcp+01dC+hzTj5SWlakWYB2Tp4uv4fwBSqc+bPXlSvsllox2sxdXID
UM4SExhWSEqcSjcUMEau2kZcuQARaRp2Z9gveGO84mtfZAL76FDOEjmtGiCmTOfG0IB7/SGeIZWg
jlpEGoImANFh2uqHbftOfeKJCRtzKshaSS0FpOKypBumGJBcBar3bAqoOFLAiOKqgHm8x/m6xzrG
NV+2l1wklBLqoG8UvZYw18EZZqZZQvenp2SGV/Z978MPgU1DC5BlLJR8tnv6BThD4/sdE8hEmaz+
chyejNs/2EQ0x8uPu49DiN6mefciyt4hyYyB4JXXlj8uZpSAR3h7EkHA53T7A76O+wGJ/7x1b/Rc
WWadXbcKllfFBcGJ4IxHbMqc+H0Rew+Qqd+HHQHo0cpI/8q2XA3OrSX73qsn7dUIUuBcwrJhd0TG
AmZ5rIoeCzvGfQgdQYk3y6KWTI1Dv9TGrJfdzcntHxVTJLIL44BFEokdvGu9QgFQlni3OO6fjBhn
IFPIc1bZ//gVB9AnT3tTZzb23KSW6LXAq9GJJHDLgUYPjlUo9HSbFIM2pthlOt5oYQopu67K+oDp
q6xLRfnIexhAQJuFYuMkN22hxS48cYKEnwgu9Utn+I/acX3zpergIYDKoe1DZJY2SjzgdTVyH5nQ
IJQ0WqXxTGeCIiji9pM/wO4/6XYA62XnFFRUsYtEykJvj+f3bk+kDUkTHrDE3t7O3EQ8UsSZqusd
yEzr4PuEXg1F6MrcWaLyksNtPB5Or7CvwjIVjgb6kjApkh/sVnIjfIU3/5IpzyUj1Zz3Nn+s4dI3
NPPyTTyLY4RLrK1CNpynTD5KG5k5UsdylUcdkqTscoL5BKBpLSFdapWFk7K1FEJtYGnNm5hBJvBK
SMYbaKEY9PzKp79MiD6u0nMU0eBJOyDagAxKFKJO+gf0XQJIeZebtJPAWz0M8h33QMtmzPxv4cpk
w5n5i5CuUCgT6k9Nsk7oe8tInCrLpDIN/CAQr8pBTjHRsysGxQe0zgeBoA86VHBvUxk+w3Ju2vgB
4CA2DZXRp3pe+9pCwxZ63ecd3emRRAPeSx0d/rAXhzlNItDTnWl1jHwqSWOtOCudkZfw5rT2FzHr
Qo3L+0ZGVrquUYy+QMURwHimYvZfreZ4UPRHMxWtjbI7FUbpY2pIDP1n2PxTkcTA/MUR111B5CE3
sQXw8fihtikmIKdT6pkFbp9dutZm/qC3xxhHdP961u0OIfZnVlO1V+G+5pxnIcXro42rf40vEs/W
zv9YjSDZ6HbWsQIVa2D7LEq64ENsrAqC0LfvPXKQ/49wa++puXy0BDPE+pdJDOyPwe+lD9A3hwh+
SCLwTHdfSHxaQ9N2TWBbDMfi3Cv+/f6Yvm/SZEW8F0AELkOXw1NGJgeNKmxO5f5djZzyniOXx2EZ
gWMRYVkpdxhiNzmEcxWdfIYsvHMb5QKAu0YNR61Sq+zE3pdunSfcOcPlhySyjywC0s1C7ydD2XbG
PLK9EHyax6nt4bw+WjdyCImvqJnb/umrkc3D4VFvud8SRN5AzFZFfLFvtji3ugHv1B5oMQNONCgx
tNtV2GX6hN1r03fcie5hCEJ5gDCSonZrRZIp8yVGps1rHviNr3dus0RSA//XCHWDLQEBx1BEg8aH
0RUzPa/7Kq1g5g23FNDWEE0JaiR1nawBeEitw4SyFTP9Q/DuUzmRkI4UKni4s9SqBLKBmJ5pJaoQ
1X0b1sf2XWTqDX8rs1FPcdZ03vX8Rt6J5pm9wJDDBArm+jQ707IwvErn1TQqq7D5/Ah4rGIp3lVv
Z53+FGcPtkxguZDHQW46k13wnEzxWBzix64mhjpefinOESu31IVjzf6rEUEe356g78P11lR0UsZO
P487Gyg0zpYijWrLt7VBmi3xvKWRaUfcpsYl7YFuUdm76pjiJmxLTCiWsJEcW1m6N7QdbbNkgZt0
CNNHn9NKfcDsVLw7s2r8NQwi6PLkz86LZqdDMwDf/OfPRcXSRP2f9qzBb0P1K1wX7Vv+Zu/yD0f7
xRybdmKlEXW8ZEaRpX/vFJTw1hkQc8rYrF+til1i3FbYD4z5+yHcKLKzXkqgnkbsZjQLseeIXASS
F9eF4PxjU5+RqMSf0zRdTYuV0bf+qE2ewvTsmnLWDKx/E/7xu5arftlP105ZQCcCascphuFWbMKa
3RtNurTPs7PUE5hW+cl96YICsPcOAb1MuFEJ0gUj2rKM4Gcb8hWytqj8aZLwelFH24njkIjhhLYH
rmBkrAbHgI1DhbJ7ipyC1Ky1QLXPrNhkkwo7Bq5UxT6M098/0S0BYs7vwNJ/p8YoHoDQ57n6T9mu
gVF3fNJieHIcKTQg7pEpLQNxfxFmu5tuTW7EMqAAjqCpmffjretxQlgzOl2NkcPtH3L1otlSHKzA
rcAYllgqMlF0/NM+1FXCIl86hHrXB7OdPxzfWyTel140ukXq1TIk2AFvvuTx1D+OzDKdr6ZxBp/X
nohZ+fLnUKxpi2JwzRBtlDZhvv8oitn+LhY/tQXLNQ0LajNFOAxGBbcQ8aJGOO6MRoC722jVh5WM
IwnhoW0qznZgHJLgL9V+EBikYnXSmqH8QubhU8fLCXByEabCPYz8A9STmmoYt/ESCxTprLmEF7Y7
wDzS1DTLfIcz5iiTjIeeoQ8TPqYnWLYEnPf6rGmWBJquA2PJWPxgqL42p5fTdJS4k6P/v3kscvGI
2eBIW100Ab3DJ9M6cfKHb7suzN3JlJdNy6wiLNsr5kKfp0ADzGUgQmzio/MUAkFAa0raE/WQAZew
06pOPTFtfUUNMtFucI2fyidZXzJtGAAlndoMsoOKwHXpsq0k0WaI2volEVmV8yimwgQ2Qhkb4/Js
kQ675+zs0RpG5L+y0VNbuazS35wbTxUBZsxaTZYGanCH9m/8JqCLUq2RJKeQ5sH7E3WtHi6qKO0M
gg2gTowK1nPExK8JJ8d/IpdS1DOdw64jtzA18EGQwF+SPC/hKR0OmIKTzs0O/gCwgV8TDwNr7Mxi
PAnavtnsakPxF+295tL7889cYe4IXa1inYbUcmWaj2moe1Ok52EBKjyTTcb7huLZTbiCOKh3zdFu
mXpHavK2m+Qo7rPP2SER59bsOQxGf/hT02Z+oXOqFzUChT2bghRnd4fX1iSKy0tHb2zR3seT/ihn
sbuDU8VLmeOny61VfTQHEdsEwrk3+1jSpjSJ53TeeAP6lsulloGDj8s1FZZ0C9ifL12zOo/e5WO7
MvdHN1t9pf/6O42mbVfX7k3XS6KWaB8lWR0hUk3RboHQMORAr2Hye5/VJi/4i/JHd8JyAbczeu3Q
I/5QmmcmDowZgNOlAtO12LmhAXgQjZlmMRRBQhum8FxhL1uSPo/NDGkbarDLC3a7bSRYKCCy4GaQ
0RzAhefO3KT8N4XGZuHmyIo62Qz3dHluP9dgVWU1bdC1XMpkNz+8ufjIYhFugKwFjOzC6ZM1dGKD
rrhx/ne8BFs3eiEuOpwu+ZbgIqEGPtcaw5frbLzCK27IgoVAoPR3bixjFXNWAw1Gftzv1i86eB4q
K1DyzwojWkujQsxqpynLpERL6Rp8itA/n4Xmtw+NLrhPQK/dbi/Q8p6oVla96FQEAHW1iOiR8qi6
PK3pYK+ZFHveDHQqjSLXXRbG+odgSld6NHMzrXyY0yioGQgNqvY57Z/0rcxWJmKqE8YooqySnv+8
bg8Y+ie9TWaI79Sm2g4zOKOOgtsu9hEple7a08wdXYXt4cMPwjyuZYp2OE1SP5t8cJQ7y49SlwDh
ON1OLpZ+CplBD0Uy5ggtqFWpwXs4yWCywt9P3ilVt+9DgPMAmVYvaqr3GhasVwHPXSgGW4syU9It
htS94sj5jWbg86rAgOAWNQJY8njjBRmPWleC7nBnFLCqq9/BjglRxouci/QtpMllkTBE9LnVBDZc
kINppbmxJuEkzpGR6TErIDaT68PyWhUK74i85dUH1Osi+tCRRuqV2oO2mtv1XLYsd3rx2PT9pGjg
uDklYeSxH073JcX+/jxXDUgDq03hYLjO0/jh9ZE7ecsUVNAld2/gfe/RgWe0mhxOq6onZ8ZNUXft
SU2fKyp/aEacEzrA4hsUDLEfnwJmD6q/cCsz38vaDr3xfiw/CPXRxJ4I6oqvO+FZGaj0xcVVpFRg
JXDq8bHn+SOhJt/gTvmeeM/CHoK+Qre7o+lwm4OTtWTcYmEh25Bu+4Vl/8e87kqOTK46elDdTZjN
/NWnitllEB/MI8YSSw+dSYvslJvS2jaxp5psyiWuOmIyU5IbBIhzY8a6tqTVNLFkw/PFtvmxnVp9
vAJCVW1L80g3iiU2MOvb5iF76DWzsDAUsK4SJlYEuJ9i7jL43SBN1IS88AygboKqrXEeelMCY35z
sSjegirySOTU6/qtORVSSsuq723eVlQuxaJq63zcUEAh5PTAlLjueEOgxKaVrASteNdVqW4Jkwtw
CMu0jH0iTASrsv1BMFB8QV3LHgyGzYTZkbO+2o772M9iUeuBj0GCIDuQxJDmZUaCnR0TekC3Fbd7
jn3BQn9Mm7LGuTGxeffMG20VP+ES9sstus3MXH574I3ZuW1DyC4KNKurQakrajSwSuQ1g2mDCZ4s
Hz2UBlTXlpnG4LRPA1BBsNeXBK11WcrRE0580tI/fc07u6uP6Ua5rHG6l4BgZ/iwh63mT9TS0e0l
ne7SkyKUlr8mRoNRVri+7rf7Q+ARBv0KVuVdJg1djzEv8RBdinXvx2O78Q0C84A2P17Z1OGuLzam
H3Bl6ih08pU9qppjLADSw4enw6qapcBSxL44pUVVL7O4MTcbT5jGnTAoUTxUX03cWj367e8doRnS
mEY9XdSZtUc1ylDEj2U3VKJ8dIyRmhZ2ZaPdgDRh+7OMMC3MQus8TMSUUmuNPMUVoEzVSO2kmsQ4
pBPaC9KasFyA6lqvLn9XFzjqB4SaI7eLZj7YUHfHF+agQqrR0xeUnWUMMKcKQPWbhh8dRnHzTcFV
/Kl5adaQe5G8mNWB0gxQKdE2tHf/Z6OQbbU3Ncx8PSOFZ7/TaQ/a08jwbq79QOCyPAfKjSolpy0L
IufCekvEr+fzNa3ak+lQBxae/055rIkMNBtSyTMk0gF9mwBaWe48UL83w4sV8YT/oXd3JrO+YZfF
m7GE2HSWJ63AbBCOgMlOGPVDqdzctDw30m92a4Pp4aqpvHksa7OtQY1/H8pCVhUNSoE3WWYxjifJ
vXGpCLSmkKn3fcL7GWTeh+tnYTbaeQEFvIhOeeu9J6bzGZ0Hyd6UA5bvVKXfMzoK6AFat6XxUsW2
MjiYNXMfkWKDDZZx3xYEbRboJt8ZI822Cx66iPbBRm6hLr8V7FYBuPKzgHt3oETvKBmESgH7/hej
wo+u4a1PV77yAx3b0pzfniPBFM4hITQ/RlkQEflenX3RBgu3kgwZGeswiva9XPq2qPsabltZnODK
1Gm55TqcO0tz5Hj5Vdu92d2eSxS6YGg8tQAl5IbFOtJ0mTVn3GkivfPoiuTVU4pOpqHWMJaTIxXJ
rbsy5/hapFVR197FcooX5YvNubJ5YJ/EhrdX2TOYwZx42HS3yLijZ1NfMDGkH/q7kJhNLfBcGXVJ
wsqSLvsFiWUpt+XoV1z1Q5SQ76/WmALONmC0bkZOWRVKUoiMTCvleWcdamyVTRY6FV9npnGg0Gva
sIqMcXoXXN/KQ6sQJupm6xu4K4GQbFK5AXFBnHrhNybBWXVOJQKJBdbgXKTCJ3WVOGOuA3CBliXg
wdtSCO/361cr/X+xd62H3mMh11zomX/omrlDuX4X13ix5olwRn721RdWLKrx86LSDa/I7jfWErEm
1pTUaFCWR8wxvMECPsyfnqINN6mI/BvOBL3LudqHoTjpEu6uDYRcLWElrerJv25NQlKHeDDVxf/F
ebeFAXP/c5V6PBUlQDjzOExy/aHbr1H63RJaA08eeQ5kDiY03HbvSPQOIrEq1WuOZtcPYuTDFV/G
ReqIsnxQU4KDnhBUqoH3OC5rdX1H5OzvPlDmzWslUR5X6Oaf4mjetUIn1E2XSumicpNFkAft06A1
kdnZKqQaOMjFA/+hniknQxNW5D2r0c2vH7Wtaw1wGY9Dibh0QNg7TAw3jmfKHq0h/+GipXcexTU5
KI0QS8dwBmwosrUGDYMIsGgaxZ/mf48+QqiaW6KqaIDec7yio1nkllbt0L1aHi9LeoJTVhe/f1nB
Sq0gkxNHGCnKotAiLzSF6zkIsrRb6Fr+WfBaLyMaeNU7tV02k6KUxf5ZYWp1+kkI9zZ2tm+e7WbO
1z821iIoy9ruVxOXBV5G0XRKINc8HAfxrtDRrBJrUeri4H+yMiGNfio0BHRG3n+aRnGqj0HHDIgS
7kiNMbQEq+naMI/bDBY5KOsAFDdH5YNbj3lKSpWwxpC0EZS9ZNpoP1EohNt+U+gIItSee/YA2hxy
Ca2Jz1sQWK/2omXclecUlUImtoJCWmZz7TTo5csuYw6m7uyBAGqrAMGx8DiptcFpEMLm297VGoat
ygUyq8wRTyXEaquGe35aHxVKkn9uViOTMjuYpk4s8IWcGhBOJ37Foa41ZNMvsSQ1DxI90j9VSFWF
R0x45FLUeKWT9EJFtDcGxnKF/0hxkcLp2eAdt7RQb1cqlln9fnOa6VXKcTRGY9+jhQqhHH7br4He
RuWy/sEdAdowcYL+rxJlo+URYAzdZE+FHofTlHpy4Dkl+AVk6Z+0AiKdMP07I9Qx8NMopeNgurGd
Mzb+78JzLqmbtNWFVIQTw0Wq13bGv/6owa6PDCcJIoadCHZMxddf9rxpwEcJy0oMhUKGRfWTJB+o
dnhbHuHAImJ6s+LIiPvFgJ1pjbfH0Pq4w6ClU1pI4hsmyZnn09QQH0cpZDFPAEq/R1MpuG1a++om
vAZdEdyq6wwLMeXMEvAQMl4TMAEWUn/qpHPAxLgtj96+Ght26eWvnjII4f3UN3p+7Fk53FrVhbwG
FkXOPOIyMWD904aHgSahlUVGWg7Ze8FyDDJozPewaDT7tZKC7Ww/MsfKvf572UksPzUOLbxz95Pa
RtHxqzVLzdzx8gvG5uIUgWshFha8HlT8DBvs2Kws9dq0LRAoNAP9Q0wPyyy09KIxTmNsLYhNMO3m
4UBk3RNOk+PNBwOCqL0Up5fmQdG53MFHmNHB4GCs6ViL5hiU6XFZ0QNZ50INm7PwfAyrx0/r6qwX
3mQIxpYDEIdTNDIbBB+LJ0FBbnnOfHwO730r9hm9S9TPNJXoXRVolCWF8sfDnt9HyUwF5u3KH0cd
cWoMVtwRjhh741kqwIQuyyBFbA+PdskyAs+AYFgoEM6/mYq4hFBz5bSC6Ghsr1r5E2M+6/8jWd5n
PExC+WcyaEHyCsRVe3PbWQn53JKvqfvsIWSUWYWSeVdqGllxPoEgz/GEWC/JiRzBpFlqlNxe7/FO
j3nZFlnYBw8fnCk3zoGi+41rxhlNCO/LGJwX7t3yPmLAV75v4dO/WmjaGdlTRNfS/Zw6iWwTpvsC
WZffSiy4SbVQiiiylTWAh2eYBbIwBWUT6xxIkNAtaLWXDRFcy+s+w0ovhuTz0PBwovbMZcXKBl+J
XU92hHm7kMny8pDu7fWhYR+5k1UkE/BXWCoj0K4ETJgBqUphsrfwbo7w1W5/5QRhxT1TbM+kTnnP
rNqux1gL3BzZUjV+lB8r9vhd+xi648NPjsGd43gWVwAJccXhE3nB3pGLxBP1eqBIzKG+oLkWjUvP
sdU0y4yEJMnIJAQsaojTg0MIqWU85400zBYznfMOJAH0cVKUWztPbEqhf5MQG3YLHUSXRgu2Ozod
AFggAAQwvCNXfRBh0MXErEenB+U8xCc4bHdjnmNtTnlAXiI3wAD7GtlOwJSvB8+qLjSssu6Vl2O1
El27/ys407fyU6W/TYRvOh+uIyHkxZdjDcXEWfC5HU1Fi6ec4GzX5FhZGoLsgzU/EBqEjBJuHxv4
pChAeI3UHYNf7M1kuNFhPSAPL+xNZCZtep6Ps+CdMjBSqDZxDjMJq7OeEtAlGYZ+Em6iag2GSttj
zXfJfkmInbcED4N9pf2DhtmEbWGDrbk/W8TLxFBjk6z20ferql+xPsXe0TkojK+/8Mw+xd9bhwX7
K4upQsUO85XA4rHgO3ilacXwLumwQfKxUizBBdlMDs9P5DvfMOrhoNf3NzCmLNvSLYVQ1nB2s8qr
oeCAR4IM4XlW6oyr1FHvtz8dJnH2BxvSopb21gso6Lxlt9PmcX1qfym07NKPQscq/AgWy7ip+WAB
VJLVYwC9ijjjxNAQmCot4apfy5x4FE5HVDrsMJFYLrtNFW+mu7dRWO6dEXSKW7m52m410QZrXBQj
ffGjP14NMUf5uMIydacY0BVXBXwQqqy7cD5JOvWpVIRwxwtRXVbvcKQ4ctUFieq7RckPds1sKRVr
OKS3QTcZLrMMBkmIb0JRar+1VCyJlbinBDXd7Wf3kasbE+SHZvBSMgveizgUW025o/B8oNIgCWcg
rLHYyvnAGbn2VBKiIV2zbTHMNRMNddnMLZCxPgs+FH3AEDNQ8TwAGLKLTlHn4Qp+q/UFe77y4lTF
U6/Opc/SR++pdcTGaEd85wrDThzNpzOQS1pv/1dmQdTN2irG9NAUhypnj0eYnZm12mAOwesbCjVN
+YuIE6/zo6oU7GjwdghvWZsaOkRMoBFjqFAoLAxvaISOW80C1eoweqj+H98OIm3ka5WqO2A78isQ
b19LHuvWhoJA3h/KhrEKJhb01Q3whqverLQLDFWXdManuKkmQlbJSc5pX2/qtqxhfB/qGiUKe1Td
kMA8aaVVOxs7IR9t4dzcPV+PS+o8kolDzLyNdKzbAnLdj//s5n0LwnIoTfLWu3/TFI62Ts7zzxH4
Pu+0ow7XHDtUv/7/uqaDS5Do7V2v/LJgJCLi0gJLDHagG8P8eaJEC+Wl6GcWVpY9WUrKsUkHN9x4
RDUTq8ePIu6ISeV3sMt8BafY8CGJbwDEmBWRFuWObJoKy25ECtO+NCfpCt/8D2jRsmO9/YD0zjP/
eZJGtk7yKbpzuL8MrTUiAbj4Iiw8c79aRoxpY+VaLhK7rcGEU2WIRHZSKkT+BUEVIImo6j42qXXv
2M0t5iGwq5ovhMvaq85TyuYyckvT1eAHh0wVAQ2MZHQ3jHCpeBF7KmtNrUZ//64DEUVGRrt8y+4Z
dru7uL9M5nrHnPW4Mcd1f7nK3zaj4VfaPkgHkjBI8jUp8mq0YAABxOAjn7CA6mDZOx/pV/dzJnvZ
LiV/qFQUw/x6ni2nR2+yj0QJd2tZnQrxJKbx8PwJLcjKs4xBBTRKk61kddG0+W843O+iluXzXJsD
HJrwnrKHQFoMCEzUb/hKLgrJ58NEXHq3QJQw2VuMmRvrdOQUCnf5Wd1q+TyInxgKJK2x2M99J0JP
/JvitlBJrQpailfwIUtCLLASXbIkgGF30CNVxfuhNOEILx39M7Nl+kDDs1OhSlnwkTLWpdQ67qI0
7yLRpGTXdBs7SJFrxm1QlWmbwKgoCzOArCwvdyVExdHs31xBv8XqmCZhUfidqABk59fu2FyGH/u+
aTAQMdw4SWx5JnOLNyJstmdH8PnjUtD3mFhQMf/mvCzPCYeSXTkKE14k36kq2khkBjm2DjN9Ucg/
ahiFHJkFjys4O5+RY386/Bsi2dQLy7F2uplaw/PpUKfJbsbvfSVEeeYFhR2NwFm1XTDHp/y+YBZe
K8NbC5PT5TPXn1ar1GAnjnzduUeaGoPTp4ShR/jIGHnWZZ9xORYs6y5HGWkEqb5fWjdn6JUt3G2N
QyJgiLv+54pGRZNWlgohK7SnxiVfHzxNhacczT1ukyBxqRmaXvCcqDrznPzd5+Krb8MfSBctu8py
cDPiBxRIjDicQ3ae5rsHAj01LVNgLgbiUQjVo3pvaKzIl25DquTxAtV/ltL5tcLg6PUiwFXLIzlA
VBSpQWaK0HGv11c2c+E4Tp6SFc8oqHC6n3IPdoN4As1OahiDCrJjDhH7Y0m48F2Jdjm0rmkhXKxP
HbFa9HOjEATTocAQi/Kurid8/FVUJWVeF1kQpZwp7f3xI84H+FQxWIjmPJiX7/sfXhBXPFhqeu+D
bFD2h7jKsSjVcWbRSJXdnNVsHuYWNiash26PinYViPUngPSTiDY4GHj15ZZEUfcpZ3sy7CnEF3oA
xfBrxLNawWSMybBtZJqhtezK9FZ+4dztM5X0+WLl8RitsAALKOPNpTCTict9wqoQ9kooM0loONY5
rn4Hs2bZaXsAF+mMDxm/6t1572ptpb9JUTFgTx26OC4L+qOmToKIs7pFQZHm4MnsXxFiMOhaDlse
lYgM+3vE6vqL0dlAKLz7ez2MZil7bigx2wee5+qcYTF1loKPviZ2AmZj7nhGdLvQanuhw2DrKrf3
E12vD1/htqVtRSJ3pvE44krfhQSLYAXBRLnAOEoCO94d5L8V20fo6Oho45WmzorbdlMSpKOB3+it
q6rl6FR/HTan9KCssChod+8BvsST2FiJGvEXTxlmPupWeTATSw6j9I5hceHD2f6s94/f+APOx5bM
Ax4+BsPpcqvmZVLWapHQy/z0zljrhmHHtCBMfjhhN8OZkIbso8HLaqAQR6Y1p3xQgu+KetCbpg/N
Luq3aV+Nd/w1eSl5JXNPUyivKq54MgDRYfky4s9E2CnuN51d0X9R+hhSe3xD8SpuUfnqvptjEAem
7oZjTgvbVxcXH6U0k4dxDyjQFXFgiILoBAnF9buPWKu2b8w8NKCqrbvVVRj4IIxjygoNs9nAg2Lb
OSJPGCwOwARMgv1cYHPYd9IL1gievM0ZtNBSqm2v0XR/o8oRckwz3dD72tNUa2F8FWWEI0cJRXVO
PtLgNcL3fj7Qe8NWCqbXD07V7hmslpa5NW1gj/Q76K3VTO3MHDlyAs3H7hZzHsDDTSzyUGJ8hywH
K1Jk0eL8c5e/QQlB/8tK2ebI2P77nOqJKbHCt/NA5/1DUlmUk59cyu3VUmrwAqUJbWU0FkJGlAer
1hbqtumF1c5aYyGYdS7GB/vSxNjCAf4yuv48ahg5/qXxS6pf2us0PqUBpPjuSk9zCaFk8Jb12i4k
PgTUHWTAc/c//nsQjAUbPIgj64G7MUlVtskiQFY2a7HyDI62fat0ve/egJYYZTjG8CJ2zKfKFMWY
mo+OzVwUSDlC6gQND++0KoqsDzHTsG9ZHXnc2VMsoxN/6Pnxogi/rgAn5V9leVzs+SYdw7fH/5K9
+paQ4PbMkuxiFSZ4kjeLWiKza96RpSSgb+Nu4mX3dCmfWkd1Rjg9mesJXmTe//bkiHG9XyD0ZgRM
bx40UI13JJ19C33AZJYiNMpzLGIgouGlwJtj+EwXN2yZmCDHKTZrE7Rzm9bazM8HJ1f9qE4iykYg
gAjTSr0Z8MC+qfBhyxkEWsTDBxn/s3pHyqxBjdztiUhWlhzIG84O8Cbf02wxZbkyFf3AizuUBrjd
7nLy/XE0mLp6C+p9OPhoyKK68v/C5R7wgJKHs0QmxjMVnhQOxFvkwrRVnOX9QpWN5bz8MWYnAgt6
KRDy/Of2P75kOpsRaRliqGm4BrYE45Mi8587UUfHIAJkk0qWEoBT2cfWYBNk0WIE66XRBzia9yXK
qa6MVnDJsJ6eSSjZIcuLnApgTgP62fZ3TdoDvUEcg2AUqUifoUysa3mIFAb/ZaC4OZbozBrBulpu
1jKk+S3V1h6r05gOARxveXt3v4IWtbNnWTzLr0A/KhsW+JI2QcTdh1Wj/xJNxvHGfs8WiOs+EuzE
MVMVHh7ZVbtcF5sHq44ZJf5zqpjygGcDnwXT8R7k9vv7dcXzYjpdolEF4F+s1adMtGawGfPnWbbT
KVQGJNNLaSgQ1lgT1tIm1mlgZIuVTh34IUi5wBKsKrU3YxpDfq/ICZw4ylP2c9ihUyhzyK9wCga5
SqGfb87YR6VnzdUctGU/u+WArTnF4rs6BE3L3vRZbSGQ+0Ctp1Lu6Rfn3RevCug6gL1dfoDLumBF
GELM9l+7saWkDG4p58e4k+40ATiHIaYjiFBzD8rVN0aFDCGhXaXYOZU1+LhHfHGxLlj+chIf71V9
htDN8rtpeF9czQ38d1MsGsoAOaH+f/NTZKJnBZF5ONvB/UgxFJtoLurKk0RBgSG1h59XJ8A8wcJk
3I6qnuKCxsU5ClHsvcmdATMdEz+VmDzRPWGIEyYQ+YmzCF65XT/eIABFkRhRMajKg9eYlQgGRxKa
6Op61Apw0qV9rM0UIG3qpHRMfk5tyL+OiIa8Ykmh/JqudobjIkQjKfwGDw0Oul7JoNUIoOtXruB4
4iaJcxUjU3VdeucUiSnkpsOFk82uZTaD3zKWh8OxMEyCKudtIOw8gnfLDvmO51FlzBTGNDj0ovN2
mRVeDEBd6BXCit/GeirkkxsLM5dC7zN3blUkTmfppohYC7T/BF6rVKFvTuaFHFFsSuPmJYKhYd/w
qwOQwD6CvNcWt0WzxzBc6aPk5RqHOX4WhC40MBbfzKZylbuiA11QEvimrSu0H+9G9/9s/fZPKJQf
GTTNkrArS8upfSEkxF2N57zo43BjX1jmD8FiEJyPTWPK3Ww5emBtpl/eXivTs4m8goPZUHdjOW4e
9DQdH2XGFkAxFGwKb9i6NdBfAEPDSU2z5Zmt/DRz9W1o2/j6mZttZxEc4FmHKSL72xKnAkNlopNm
Li3I3Aveh4KWC2rnh3w1cH2t8vvtXvqwCemGtoqbRLXbvEdkZIQKayrpKuSME1urfvUbXqOiJKd5
uKIwrh7gBLMF7h/FtI+cp3zS+Ql4SsUjiJWUTaZT8ciMnf1mKppGF2wLbrjuQVRBHx9xVwK1/Uei
ecOAv9kfodyu9Ls8kKVmZKrl1W5cnJcZwmMKwSFYm50aQ8M5GTLK+OqLNfCRBWp3O9I21gKyFAvD
gB1zrYixbuJyZkKJ3eClFaiRUdxDLDT59g/P7sbp0uvmpGBy09qSsuIw7+1m3x2rzzX7eQFyoi4f
T2sbB4YlnFkSTFTHj1qlCbKhoyo4Ko7FYCKCXdpl6XB1Algx2IZGhTWX3D8VhdfD1d9OxUPd7LrB
ck8+xNceo0i64fSDuqiBOultyVAlEXf9IQ3SkmHDseClXdw2ZcqFl7umYvKL5o8ZsHayocdiRn1g
+iXYjQWmG62DrPZDIOZEnACgsrY5Er5kNxn9h6Q6cC+9K1WZBOYRxuuAJMIwNwwwveBDyaWq9xuf
dg7S0SN7tzYFstIJpVhrIThH5xmYEGFFeA7GHfx2nbeVm0CdkljeZ0XCOyETWVHlFp9OdRHQUBPv
W5EzlxAMxvvAH4FRLfPHmUSV0j12N+UAjm516SIcRRyx0GA7LkP6Lb5htL9A6r9KUe/EOOZLxnVp
JG0nV7fwGaGHx2WTv1hJ5y9T7feBWXzhyOjaYTFF37oN7dRpjPjymtYAIG0YaChgKknF6AI4RPMi
80KkihoZbMEDUAc9D4rmM4Nu73PqzYn+4FZbS9L8VJ8+/Qj2n76ux3j4c/OdUp+k/vI0Y6m4Rex/
QzIsBNgU5wk7z6BQBqLktHCMJVYzHT8KuW7n0VOCoA4DPJ9igzhdP2wIkH3jd50QTl30mkzNUMI0
07IXMh/W6NMgayoabQiuFTPh58IL0zNZ77uo8JzDCDMoXgFQ5Uu/JGb2xsJNopFgVFo42AjxPxoZ
aH9e1X1XGxrnkMRT7f5sqtL8ytOYj/XXiRPbn3SEBVIBIn3PLRfsIqpQvuybbK+CJVMIdHA8E0o/
f+A1Py1fKXNepDwDKNWCwb9eLgYURkhYpK2SDQHIjNwOU8EsAVBnh9lr3Pfr1Nl4NF2780fpURAM
q2IGB/E/CSwiRCm3TQ2WSkPCT88Nv60vz02RWxkzd1uGr6PCTN3cm5EZ/e3j2k8apqu77HAC/8R3
i+XtDh2dM/cSF2C+R1h3vAQmabgBXCGiN37XESz8mjzG6nv2i68dctY7fCIbBhev2w6xVd21p6Kr
t6kvJHijVBbIY+RT9Oyb26CaTuHK8W9u2jGI03Bc7YLyOsTCJzgL5TWqDrrtXfbpGsPZPP9PgCz0
eh3skeUQ5PkVsdvIzXscsiGPHDHDibNS3TW8OcfwbLqlDdA2FxF5nmJ+EUPJu1zW2jyrkod7an69
3ms50eF6EtArsZKpiHBMfv2TxocJhC7IvO/+rqaaaYvDWc8TE1ASTlw0qNcNYDcZkALZCuOWLu7k
SjO1Wv3Xt0Y3uRc/Ui7myap5D32Wn+LLL/PBTSwo9EJCFS+cw2gXMN8baZJ03rQsnGUEhHKpice0
g0yk2OZEqpOXTjk+1TdG2G0PYVOny3nSGO+RR1YPNcoku0BKFedE90YzSb+SzoNm3sRnbydl1kgz
xl7wjZbx2fTAPnZXWl5NojRXwDmQtlFBpbRqMPfd3hT7qBCPKfeE2XqdLZpv8MCgqwnFdZRzj9LB
v4+9K7zmUUeGFOMBGkNxTsvr0tUomOuA1cG3n3VI9SakKYSAvYUS79UkfjM7ETq+ewlQSyhAnZNj
pfzwGdb4KiQhnzl3Nz3MUkgG63/XWuof0fVTSPYolwEpb0KjPrq16lrL4d58mHNvu3rdo/UBOpIk
704/If2htAWJ2U61CIvpLQFTpJ66HmO5O+kKulg6W0RGDERskVWhefn6BHpUVKGT3VrUuFdi8Rnk
YmeXZDDyo62XT9xsaEH+L5WttlBPtt/Es67IfOMm6QicaxNS2CXNdQvyZtJbVF6dOuysZxdIq0GX
4TL9nFvZVNiRH1iBDeyqxFK5Z70YRv7i6Lo8iO8L5NIf9VxODCqYyB4P3JwD94I27rwbJEFM0Qag
wB4LZ8jaSN16npq6IuDhAevNQ5UH1BhMCaGHsD3w0PYGfK0P0XlRUmQxycbdDBQxolpjwmgLkaQN
TCKFVGxKaTWhgSaMPVjqNQOaf/mwmj0KqHAMDrUwvfyz2gBMz0YjMF0ElG6TMFl971BBEIuun4Pc
0vXwXI5wuxk3W3kXNvKy9t2M2CjSdJOH4eWe6Mh/G+KLVNBYDC4GKaHSuSOySVu9v02eGdjyBETO
kvy+1iegRk9R2Zisz1lo8zC671+NL60lQeux5U2F7cZeoI6HCwX8wBNcY1XdB4Sng26e5PHaIPTt
Jf9ar/YKJAFyjPQe9+UFogylizoE5yUPcJqsS1meZheHENKXWxW8WMWJImtiRPY6iBT1rMa8QAHa
CK9JKoaENCevrl8stbY6MGIISvkknOZwKF9c2KEbbx/nnkiKR+Mi2Ri3bIhetT0rWIFy0JXQ79Se
0fdjytqJFz1O/yLjAIjCia5FtjowMbAt436fApGFX1qu5diA3SU0Q2+GLKz2EisxDT0hIMehtjz6
qC6XE+BIPyORJpWTr0NX174lWyY2JigfZb6je+tUQxmlESEYVp/0/PDZGsYVQ2wbr2sfLZHpIRPF
riErdTsHHdH83ZNupSKEW+bghpSdU7QyHbmFIJib6EZcayVnuaAeNsRGYG3iGvA4ZVU+OzrdmDod
nQJ7+BPrpsIm4eBDEXhAXb7j/+nz2xlk74xORIDwjBJSykfvo0Bd6uXmONYfIJYHGEbi121nCcEE
2gF69aehTLMfBceUIctj+bHbt95Rt79d1AKHMrrZfewXkAVfQZ0DN4D36Zg5U/w3jGvnA3yDMBDW
9nvU9A1e9VxYiCjzShyVwBF+ZaJovzdEdOeNuskap2bbv0uxrdIQHvcu5r0sJdyleESEv2TM89vL
0kupgtpyuNZktK0kU3bB0sE6R8KKrZUgSeQglcVQvUaJVn14p1REEkoDsFy/dUImqHMFjQmMs5E4
EF7SY7QAK8feGMCildPTZ5Bo5LDXOJaIVgTqyNFsB5jJvNh92kVO8pvW2QlQnY51ly5xwr3vXVw4
pvhlpStC2dD/fkRDp7GmuqN1QCLOI8iJowOu8XEodM9PZsOagceP7FhDx5KjFSQrRnTpZ9uIFr7f
5h2d3utrbzXURmsVxYFUkicZrmFGl+3jJ6yjnuKZHgmow8BhVZOZf3aNBwL9e2MF3TxQ2TBwHw3z
OW8B5mQFm3PmJbUPGPu7td3zb2ERUnQyUTGpB/dhdMKX++/FvOhAZbN+Ep7uiWrBI6n3hoAKHZeT
g/efGLfMKjLn4H7BNd92juLmv51fnKlFQ+A1tqvS42PdUVVAS8WpWhhYE6bpWogqqH1cxzvIbE/7
yk6tzSKuuhfTVAdeagvNWUaoxMz2F7n4Bsb+xLbcVSEy7lW2UKStLmNaTSanasH58fc1G3MAngSM
9xtMw2JWngEcZTrdBEwBOAgTzRY6OuFSylTgr0GzvKJ6rDx2GDkitOWlmnx0OoMtvdO6Qw7H0MXa
P/iPTPyiYeZpmAMNK4Ly/PQeFh+3a1jKX45h2CyQAF0C5FtzD5dVivdTcdm/YOscM6maNT2510/j
k7c0+JC0OEhaDgJ+ull1UQQo2OxIPzs5rTBIM2Gp8kmidTq/FqO27ZARWei1DuX//5IJvzAOtFX2
wYi6TenxZ4WZiLGm4lMpdJCpvSuLNDFIx0pG+eSeA7lgcd/oTSiiyIhIGIeed1CiKExHaYOveQOq
OdJ9aqVTvArIw9VlTlYOiqpVXGwwYev1MshtcmkvLKs0XA4Hyppwd/qUjhkrtowhRv9rD4pf5Zyu
BbHiIsct+o/hNRTfhw5BklVwKi4oKuMk7vlsN0x/ENpDX3IFNUTUYB5VLNTJRxEGbdWF6JG4cV1O
Y4mI1kgxod10iNSMrUVEooJRJfm9J6NSDe2p1ovI0NlHQXrg/i2el61wH5YBF8T7ePp8dGghKc+N
XlhXMsJXQl9jJo63cX8G73MnAb3KzrlNk1cBRwjLBjiyhd0gq7wBDIeutfDV0VUPafdmzGEy71e6
8pmiQrpsbqlYtTMg3MJrlUqbPsYwmKvgw1QbtEj/WLwssTcib50+Y/7irnZHC3R40iNKcui11zwZ
RHWQsSQ4yo6/zIe8jHmgwznDOdms0/tFNVf/CHyp+qShjwZmTxik9F/m2MHaVCMY3Sd2ZjmG8Dce
grvP7YRHkGGC7d5FSZL/8PCJ7Jw9rgjJ4dnQrvHYAYrW41gTNCWtxjIoiCU2pY4atU3fIfH1QVX/
bvoCgFsQH78jOxuzvoF6pp1gAK2gEGyBunj1MObTiEGLBPts6nc1vpLXUd+Uhb/1hhZzP4vqi6D1
an7XrnCmph7Qf2wJq03ZoTmNcMWADM96SuZa2j6jgvUwI8tZa4zgMgwPDMwqCAtKKV1qxtY+/oC5
ailXY7B0yHUVgNxFvY30Ba0+IH13XcC7inZ6ukuQDOA/vRNb8O6K8MRSlnhrJr/8zuDf8NtjS3oK
neheL7vQ0lakB91IiyREv18zGG5To5mqS07NimuK6x8IAVIYerLIyU6L4u4Czj+jpGmn/1rBGi2j
xDCrww929Nu30XT49J1nzsicBzATaGCq9DLSh07c22caznIlAAIvkmShTksbubM/NvCIFMBnB598
uvB6hqxBuMvquyOjbYwY8An0jiDafbQz0gOyGUXhrPmm6w+1jSUEavo0RwKn2DVNXYtvnPbkoRk6
kjm6pZ1oGpq1sKoP87dQUpdJjyc/A+7NRHpT1t91rvAcEvKyegbLQup3BTmAhhFFKlnIh900+HBX
qLhj1m2/BgBfGMjdDHCpGxEyi3z5P7h+1TbL2SlofyQDVzbI6FVuj+r3FTJQt2mvgsDPXkH3XUWr
ngbb9fKE72lgAflhlvlZHnysAAEulbTrCQs3uKiJYxp5HJPoK08+xywGLIFnCzT9zXOy925X5rWU
7KuM0nH/RgqJoSfZLe7alZI8DKNpoEtVuN8bXgq7EAXcjH7upzNO6jY5fbvYS6HvmaKCXPkkCH7e
3nYRHR/qt7lUEmpb3VzmX4KIsHRbepYK69Jcfl92r9YpuwApAKSMQi7CJuaM9CXQBY/8If+7xIbw
hxMeOKKbdRo+ss1VqXGZhZJEzJXFeJZVjtTJIrgz8NWGmrRdb0BUtCRIJxJCZxI2z8Rv7baZHblq
AVv2vXKbAh50PHE1aaQRwQsXHmVGCD2J0X/XsHlsDCesZO8C5cNXazljNzr9zUyFKdGCL0fJqq70
iKMqaAGscCdFT6SHo62EU+ztuSrbFWawxis1DCV5rAakonTPlBnRyykZD5Lr+njZgKFWtD54wpg4
gKdwN3bnOAmLnVN1m/bxuMSP9zlS5NNo6lVghODsaRRhAOtWPbhQJW+QMqXX7d+zYhBdSG9sznTu
MGUlWeHD78Sis1SVGculd2Rr4KbdIdw/09lv3Przw+qJ0nxw7dNOlgBshsHWcCt//ZbL5aYT6b+g
qdb5HBQBha3z3fXK1NUCJwyCD+QonVlAdmRT6boIpQJBg4RetWTSUuDQY61bahk8QDK7VZtCLYIn
pQnPF6PP1QnfgL0dqWXUOIT6ONC9j0MPtAIxPkrEdD7Fd5j3jW4X/S/jWGgnzLZWf511Co0R6Jsb
f6T0WggfQqV7JV89tGnBKnDoCGNpOSiCmlEw/cSH2Wri/eaUZGMHc1O6CWbMLOVSNoIK1xeaoDWH
jVVHPm8MuOExH231uiAOxZtY3EABBgTbZGD7/qmtH7seZlNX4WfzOsw2dl+dxywi6T5Pe+C71uKW
diGFQwkgbLjuHtGPcGNo+IcRKe+JT6IWDlDT3zyYqNqiOhOoksn/S0+sviTR61nvrdLLHrY9laN2
GnmyyrTjkSCq3KP2U4ZRCDQphGpRMHyEgx+4JOQawh1Sto7gba8HZL4TLYudIIymcgSQinfElnKL
FWFaLy3kRNBFiPs7cTC5gees4i8or8Zh7c3HcdCXHU2QCGkYMy/OpGnCoV7Iqpq3EVgrTHeJP4QG
wFxEteuGgY/hghiGASaJJfkA7N67JjA6+lMNiTL7qhBkCFoM8OCRKH/YJM0gNHcmsFdZrYCecoGr
TnBrMW+WouQ/w2w1yLIVBRCt/AxDS5Moe4qSjKayI5DsXFKj0u9kdxLkVaCuzPtPGCzbJhq2Kby+
lGcfvYhRgHrFLKimsb7aL7T+WJ8hR5Iwfc6xbsPnkj49gffQnAQFDwVtiP7ahNHN2GeGCFWLfAc0
n5+J4wowC2vSSWyV/q4kv6ji2ueltcYp9tdO7n+17NVTJCQkoWJQYCEWF6g1qiq29EIrBmao2SU6
FX5zu0Wf+RFHvhkwiUnMBUyib8Qtm9lwxogc7QAVjMbvQgUAH8/bj8k6js/z60DNzG+S7v6GpLay
6A87+UkENFfRutFw0/dRJ6MWOXTrnsOpcObCt7B7EwRtdB5VRz3sX1/ILg6DotHUuEeNFGlX+bbs
zcn8t1mmll9IzWO3NubzMKgxzyfC7Ii3pqntVH2yYIUiBT3EJ4eqTEg2LOjncL7mFFllFBcT9TwQ
3qYi6etg7EUavN6rGm637J2sALmfmQnq3uZ7HfA6wAETfmVb4dToBtj8pihxrbb08MPVthTGSkHV
zsaJusdbmgcyjlB5/+b6AxWvB4vfDNmQZR+qFOAo8fa7rfAdAHG1FwIDkQ/seDW/QOtacIVlqOav
V5PKmRYfHsoLXRbyKx4dPemPbtsDxQR+n7HQRjMKN8Vq0diHp7wKNF6nZk3QEoyLSzNfwMeKRvde
KY51tCvJADMKFshy4xULbeRdv5zGhvNSrsFPvAQXaGvhO1r7+BGFN9G3Mnws/qMSTD67EZ7Qlrab
9Lvax/vDSFHjvyVQ4LsTuCnXUDLee3TLJZgWwSqsZrPaaOrl2mv1pLasMN3Wl/YLp7bMoJHrvBLH
bxqxTmA+PQoPa+lQ8++Cy8k+vakuQ7IL6ZxYgCttEjXjUSPg5iO00apJrLGFHGsrPzAFcMd/MVOQ
/CnIFVzXaP4EhtdVIEfhYuabUO3IlmPt4SzGASLT8cTeFtxVx6PPRSEgy8pS64gf1PA917hS8NHA
7+sVx6FP5+fXgkaWY0mM9CofH6sU7PJqfzBvIw4DGchvGTKfv4QFrYYPSBmP6KtJk3wQCDQ9SbT9
elpz2VtIrfeIVEOmqaJDb55LNOR+b4tzWBsstc6XFqWBmFXCs9zcnpATyFApIsuVXwVOVTOZKebO
Kujwhg/dYY2ljnYGLSe6Pbv8HxuMKrfszp90R6ByK8vP1oy6EUKkM7ISQlnEJ2t395uybN/D03xT
TE6NFXJKI8qEByS1ia11d2yaahwg+sC+29AeBj2YW371XvNkB1EtxjxbQIjV8GeUQUNzdbeawKnU
dgaXiZzmmd8HbaIE+4+YB9Fdv0/SQNtYZcgtOE7tEvoxzY6JD0L4vadLGAI5C+D2ZnG0YIuA4a1W
oUnczQHWkqTsLyXEJlEl0YCMEhAeVmWRw076Mnzpsv1m9HDcncQsLSQs+WI2Cqd8RgE2u3e3pgL6
S2HSjQyyNCz/j62W9NsH7KV8NSjRKOWTgouGWLUZ0X8RHYTYTtv6gHhrfWDl6NMHyIOeDGcK4m5c
T9+rtpAeukDqVeNcIeFxrL/bcbjtZHIpYMa4g96Oq5ZqW9RPZ+AxLHmxuIic3yutQhndAZ8bko82
xXwOu9l6F+DU96FbCfjj8bbDNyeRRdfcdCIYNKawAed91USrkUoltHP4WzefvofQLHjKmGk9cgje
K3l6t//0kPPYn8mYGXMsr2UIfwIum/rkgNN9+phJLt6nRxLjjVii9ynBC0ysZaDyJvmoW7xiNIyF
HKvA4WY5BRyiG8FQmFKXlhMEaDrkq48BquswNvHerN++vxU1q6Dk4mUoqDEhF1Cb8Q5bBwPZvi+r
IB7BnXc5QT/sBlp4oZmxd/uK6Ls7v1cwVfKvsILy3FPM1VvnBmfE9XEHXdbgcXyn428RzIEQA9q1
XNP6PBfcoc/9xPiU1Qe7/XCfxD3FdT6kUxBIA201RS7HR3iJNJ5jz0bA+/6mQWuRNGlUrmW9iOQz
RcTr1+MjWxunVNExaBoaATbjhdEk8rdzNKVCQ7Tj4imEZa9+/h7gbXvKNmpAADgkL4yqmWQImQsg
qjdCyQJ1ObJ+JZHWGASkpsY1KAFm4MoR65OmvMHaVcIP1jblwk25ROpy7/WP9wKPGSlS/qMOaTvb
ELQki8L3fowlF+ylznRPoM3SdJOLEiOl41ke2bskJNWT8PeCVlH4FIb7vzV1j561QkgurkVrha4t
5vRXU4472bEMkxqn+c6wpLYj1KTT4EJyZtBWImLlOICovj6gYlEpHLpKzLnd2cLfeyaM9WVAldoU
jgHLLvMpnV4Z0MBs6FwE/wlZb8ajox/QTQh1XZc9EOWK+Aphy1KCs87BI4Ms/8I5lB0K6UsRo/H5
X3KJ4LMFRDNsDrqq6eCxpOxNHdRQqINszOFwwL5oT4AIVvMP7RXkhx4aMytdO1Y3TDtzEz3cChlI
MwJP2oqelttykWyTL5OQsMtrooS+WBrQK8Bz+c426GQPDELfDZ4GyG45A3/WJ2oSvil13+rWXag8
8Wnj37+8It3qsY91Nbozi88dduFcJHsp3LBoQR+SjVe63iSOYY2DLj1J64zcs5ovV/AGPXVp1A5o
2Ud9Ri7AYJVmnDhPSrq0cn45FwOtuKWbUawJ9uNovwpuAArhDZlbKXxOWUZ4YYag6u/iXb69hDmn
PBdOowOqEtgYzS9Ian5YMJwAjUs3khF45Cv1YIJmEAzL59LnXGPrK3X9chT1puWhCLzXhSBwt4Mr
lDz1Vpza0lsMS8d2r7IG85t8bTrLe12UmZxSBNmStdL8oSnVTOqOXUKcHoyCuGOpW2C2iCyrf15y
wMZWqzJdktGms1pGQas4SB76/L1Iye0ARyKczgZxVuvORxr0TM8YsQ+jgUMP1kCYd8mdBBoJYbyk
MNXi/TCBawmqiUID0xHnWq3SVwvG1m1u3mJ82f/JhzTxYy1c8Ml6aZJrtjkzv3/Dto3fSv9eKouv
dABJtqOz+n30N68JhWGmkotyBjJBbmWaP4gRbJaT9oknqf91ThThSuzJ+ECKmXX1iKucMZaOFuxP
T0eUKk4zaR98A87aDr030Cmdm9U9Vso3C0VCTPtrZKo6d3d+FaCRtj3qOrXqc2STO5j8uKSc0brv
brhBrekgAUY0J8F1VPcnoNLClLXYjwuHgSPG+oNemXP5mPaAgGHHRienucCLwhrAB5trg/Cp/E9x
K8YbaZHN2b/zbCVZgp08yiR90S81kCV6ypvTn2Qfc0kf3Pny8y7zoSrL24OrmRx0NnsutO22+he/
4dZ/LoZHPkH6cP9WTsD8oSswoz4qCArERNo50Tealibni4874k5ikPn3FF+BkyjxCfcZth2J4NI5
/6fu2T679zsc0TQghbU5XuZnFx7y/eXijvEgA/sjEfsrz7oAHlum6At1Km1Cno9H3nVhNMVCEl6A
yylJBoJVKU9Qm7wbVmAKHy1I2e4PeaOxLThcTq6KYFUt7DL6d+4swTowVjWU30TILj1wFvGi5sPD
EOgrJWm3Sl6irqmmrvtkpLG8Sh6iLS4DNjdpD+5Qejg4e+tivk/cfEo58dT0Hww1poBjvJMDRciS
I5Vmn/09psceryPTbUirqRo/nMHpkjXdi4xLlht3umL73Zrt9H3UgFVYQF0tHtAfidLQ7jvNtcAU
IiBN+7oA2biDQsDsvrlifSYuxqTYfJWCJQiAYYAPtaVcUCZ6KoIIXKEOYxu7+xTab0qjrKtIrlh4
nSOxPFDUmaFnxPC7089sM5ddjYwVYHovIqp04rD30XSwTfQOe/pjYtqnnw239QwCCrn2CaVYaD3b
y8SBlSIULkhzKMBkFgeaSr785b7z4LQjhTNyCAJTLnpPWQwRNJJe6lunjiBA3PiMnICAlibBfFyv
/jMBbj+RIuLtc1QOR1zzxlT+aMr63MmhVUpZAb6Efex0rS/T3BtkHC80M5zPX6xZu14cgh41PUvu
FjPYtyPivRbsUdyaBf30K4O0gk+uMl7/nzKUi6j69Sd6JDHKQv2B+i/1Rldh2y5z96ogO8M+MBMr
1+0c/HLH/P5t9cwV6UyCPT0GHtk14Nm1tKXjll10OXdDCktm8FSdenMyK6XkoNoUkcpBWNFUgxb5
MxtgXMxNccDincKxxSqHfd4nC8i2XlRpvgAM+ClhL5qLID69oE9W9oSqkdszZ3O38i3SHkUfU6vd
4D5ML0v5ox1YtdLEdzwFOEo/1HTapwp5Xwq4LGdp2m5EPgQM/U/aWpiUjrjwRTonZSti2TI/sHmL
zaFATG4fr29QylyMR7O9LSPgwLQ4rh6VqpkxzpvCVboNfhvcCqlYJcCzBje4FNVOqg7/+m8nkIvq
R6BbM2FIsrcQuxkqgsQhK0P7sbsaiEuCVVhdKKHwEIAZHYvpubDuK4E9/ONuG6bBUqms5/2NDfrb
zbo1PGK5dfABdcdv4Gtz5RvWc+Ji58jSIyURg22tSVXbcsqHbQahXcDT3nCPH8XcPpO7XroGaYtR
bJfQU3XpOV837s03QFR7giIFCq2AkF9wudxvJdhs9Fs/PWoaitGf4w1nGwR2w7FV8PhDAzBYh/Hj
Qwgkm+I255SFfbOw3JkOrpDJytnzRVj19BMOPPnWJbey6qqLy+aQaXg8D9EB09ZBYuAuGt0YDRS1
jfn8OQqnUq0VXkJo9wAYbSfgaDVGsd+izqKAB0ZerFL98PgJQgoUM3GACIUGr0SUqWNeTBlvDonj
sW09InLSkDsBuaprGuC/pMRx+neNISvxOx/ei8q7Gt0z6q79JBXwTjzc4CheC4HQpnj6EFna9alk
KO+wWiy0pAFcsZB/nSFLqnaWi7P5LrYCSn/7vwt/vlncG/yWeQFtlX14zJg5XJOggZQV9+buxY5T
WaH8+X5ZClbmosne3KkS+CyPpgB9fKmqg0Y1/hS/bR63k/RUHaSA2qjCTyzYf/2ygeNxdHmaWQ7r
ZyaTWab8n4n+91jD8sThb4P/iibYxjhhJnUAweMIIFT52YreM6SciCLBPrloQ2MidYThApMNHiLv
EzucasYNPog27+xriR5fGygfhoA8ncUdl9H36gmGWfwnpMJyWf7aZFyG80pf9Rz6wzciAgqUJAJ4
8o94ruayfBplxCkwXWKpi9PsEl/s7ahdUlha/ursavmiu6Ana+pQlm3CM4AM8EIbAnMgsqQA7tjX
F29g1X/yirsXgqNLsbsNMOhr0luX46vzYOLW30z3AGq21mf6QuapEgYD6RrjFH4fLmDhMCI+Fmtp
JCt+C9nKuhSCcwXxy9ViXNGarUndAr0KHBFdh7leUr6ei6KijxQ4Y1/oTPUz3A9TGBbmcxato9mC
Vp6+JLMYhopYn5UMIl/CEVaPLCy3Rcmpc99Xm8WLUoa+R+RWVgcKG5FvpIurI+1fYdy/Ph3QfXP5
O+nep5a9thZYaVjI1SqDp6hPD7TXonlLsBEtBkHuXedd+kegGA856WPz+nzYMWqgNUuO4SitSfJs
+cRVZOhsQtZ82W41pMU9jzpLFoNfz8UckVRPrkacEtUucu7EbNBxhZTdj0RA6p9xZJP03SK8fHzC
ISbX1uZJYa5oMeKrnUgOXrTHveBV3YdJKeDDB4pQlDwBBoahft+gENksNlj2KqD6dnFqvHWWEIkJ
M4Z96CaJqLZQmlR9CJgQDGDicWVIPsYyJFNgKBiMwMikT0P7lZB4HaLYqRQKcxza2/oYnAh/v/iF
XHKGI9BEadI3shbVolLK+1zxTAt64uV8qAJ6axLrG1yAzPtITYVflbRFztItfyWC0UNo+klQIfqa
FbGwXrornqnogqzk9EUGdh/hQ4/UGj1SMF2Uv24hvbJRI+V4mASgYqspez8mnT8ixrRR2+TMcm33
ECBuvBUD1w8O7UJc0Z30N+K6VzK1cYWPisYBP1muXpoXNBv2P0eJELgUFpFNJLN5OcW6jZanhTJx
hV+yUbCN57BaVdz3vE01NdUDVWLWPUgZXuGzLnJrsRUtbu9g9nZeKzQhmtM+pYmPI12mWv41UGxp
w0GyT5txwJ0mKA9dG3Z56iGD5bdMSdVW5uPlsjG31mn/bIouch6EPHNByFq/ND5L9AdntjlIOSCv
wu2NNyRHhZkaw8cV6eUQQYOJ81TNC2nFNqydpek3ZIDWRxasHILwZBoO4pYlJJGnPyGr++KC1sE7
3+FgbCgZgdSfkjc6QEV00PEXCtufBgE2wpLqHYqsP7pFCk5dj6R9Q5TOWnsz5QOdV/8qK3beM5ed
bfH6ID0XZQrBe9DaEUGs5SvsL0Ha3K6rSLQn6pdavYJlG599lBxAKsjm2lpqHLgMn4hu9udcclI0
pgIlPRAx1fjMjPxhahVSWRmROnbRXYRJRfeLxPrS7TJVQsCRxe/fToACwYQ1ekBLcJLG7EuzDWzu
okDBjHAW8pRd1vIGt0YreSH/U6NUToDb0t7zEU2dXNID5EWhCv/P8VjytB/IzLj0sr2UFfh0vYff
brWqvXIQRoxTh/3PaB/CRfEPDho5z4NySOL3ZaKEXeNQsKw6PlcHCq2mhIRjCczT36yCiXyYC/7b
DKVCD7Y/oNd+IKnCQZwlJVOczcpDCiE+3qe75VZLcJ90dP9HrKyo88X0cdopt8En3NMsi9KBjOCU
4xPQvGQqASyzVHsKJsS2OO/Dq4R1LgIkxmKFQjjqdSFRoQDJkpRr79OYPVLO/Sa1CXcxS1YAtpPl
T5N+gc5cvrfZ+pEnKgDUeto1PZHNlz6iXMZcZmhDBzO8RP7TCPRS6DJXQDHp19rgVAKAqj+lbYxY
8zZRFu/gvp0FMMdg1YysY2cZRJpYLj4O0jWHU3mgdmVNJGUEhbjZ1sbv0jtHKd4CUKmY5FY7qs13
ulTWgq4kwhuAejmF28lxYbb7l0LbDoCszgTqtHmPG0Ci40aFMuQ41CBxJjklHZoMhMuC7Gf2sk0S
jTTdtoI0DsMPSAavs1j2M2JI1P8YwQ0iNtrerJ618gwZzZTFdaQktitgMwUGFKFjUDRZZfU6omiD
bG7TEI1ruCJ0A4K2W5G/LClPSSPS5NMYnZQZepfceGGqDYdGmXoEFmUAH/i0mVQYnpMrzHnPKtaS
7YEqKx77T6UXN22+Y1H0VdLqxwErgJSKTdRWhIWKAlZulS3/OGKG0/wWF8tkR0p9/mLf0XxY7oIi
/B/drjzdtN3Fvs43G/VQaqoN71oqROY9RiuguUDkZbzliInUHrj275ZNUfsM4Jcji1yzKisRiYtJ
i2GnLo9PzEdCEQbLLKgsTuHZbtOe5pJKxsQqgt6qoMJQA1RflVFTTLji8XTHRoAbS4VBMZSIUiAH
NOV9xF8PwM4rXvyH7FzMZnvSMencQDhvKXqwQg4jkrykc0YWlUepGUTGbNN+O1YPPnhRpLEfAQXQ
NKWd+4NxJpSH0BBfMXko8Q9M8VFyM7z1HXvrmZFA1oJczEWHlOyHBTHd4iqsqS6WL0/xo9JPR7RY
QPMME+S2zTftq7iA3PV3EpDqvtjuq4QVQjAnPMc1nkQoiGKqn1Zivm/g9yR5ppwQT8SLRFZlNSlb
6TLYgjgh5tzk1t01/WJIG8Df7vsW5+ez9d9Gk7VZ63twNW1MaWKU4kUNFKZquzkU7bwm4DLAUgue
yzTbszcttrpUhcUM3elbrVqwE1vDedDEXP2RNiOV6myVV9N89EugAF8f1CjvinwYxs3hdeWe42Ss
3e6QLSGAK331Vvw7fz073wvuZvYHg0yHia34t2juIqQMN9ILpx1+cIv5UQZGQRDDtA2nqTmxNzZX
Zgnx1sg1rRKwXcH6VxN0odvZlrWGxoAuIEzUSlmH4OSeysmdw0d4TUjJ+1RfVEPMMbPp7SboP/0J
xRa7O1+VJG8T0MKIa+xM77KXBUKWKA35GczutfywzjO4P2X0xltfjc7dmlcVvPopfZsKaMsoIFKN
8nVCVXEsRZ8ynj+ylkey9wOgRm73lUd2MVs87JiAEx6gKghfVOiH2fcswaLjUcq/3OAPnawY9xcN
iAa7/rrAA5BKNKiBybNC6CV6nLl3yL85Ff4TmpGFa9FrVGC2sEUKX1OFK9//+u5pD+ObMxox1gv4
D/KBLzIYKPECjeEeNp/4lTtMhj//oWfePtUY4PIk3MOb0YUI/7vCUlNLBt/EA/zAOEYJak/NvH0/
HJq7dVUaNANfu+SWZ0Dk+7pDlx3PxVhjYaNXmWVtI91eegP4zSTy59yxlc+siQe7XgR9S+du+6DN
GtqBoPPjw2rfupEKYQ0k17F2Txd+M6vzosriHKbfo6svQyK3QiqxoFY2P+zP1zz4TjjhEl9Z4YGR
JKLiumhMxsEmrYoSrV5VfFQjgYW3DQk+sMwYvOwPM5/5A6v9ZLssxnBeiAngRtVsf+oi87vgfFVY
bsl84IDc9dvJ7fPXlaxu0rKWPqmEk+w0e0fX/CbpLXWXcATZnMhFW/BXyssUtZbS0Y3Xm1mzbnQm
Wvv5l09HNGvMKrNEuYFljryNO2GHgmIqgIKtms9N8m/BwKHoDThhfp51u2yd8L3Ylsu5D9nOXe00
oDel6SZuLNZ6ixZdRAfxbgVpjHYwEA+aUTi2scKnMzW7x5nJ+lzmcDCfQlUqBdJpsjgdL8ZEt/GE
Y5W1KTCbYxTbP6Z+HgvDp7rKt8uU7OKaIFxLQ8OnDoYTVtZITLvHYo/1so6JurOLZq3hLgGSY8Ye
C++Sy0fzXVax8P0My16SITCGEYTTHLLT3sPGywsM3c5d6BBu0w530B+laqGRHbxb991e85K6yuy5
Xgs1HGo1vL+oT7t3mSDA8iAKKzx1Rkm+DnhdJP72XQgD8QvijkTmuXj8+7lvA2q0fOPa/l+VSGXw
hQYoBQ93XXZv5Nmko6B7W0kC736I57t5fK2Hv8vfo473G648abP5SR1bmQvuwCibZafciAoSqTaL
kPqjCTnwP+hmudFLRiGNhcO/slqU5Jl+Y5AsgoqhtG2HKoINWWgI1Od5bjqmjgd21fMM66IA9wb/
ujW+aRFZ5/akcX9zGqgVQWhZcal+qOsMcn3SfZdhWVP18Pscc9qA0HpChg3mLaQhDjoGMlIKOyLK
F7Fm/+E6CHLXIUlIfVhncKg1dlq+OsAkXeV1vd9twlTH4PfyuG+7ylwL9R1cDdujhhK4yh266uRf
Vo5HxZD4lUiQlX3zatbVpQil2WNJLba3usLQV76tpD3+lIfMcE3lEn89VE2FzEQ+KQKucGWYnGJS
61rc4utHim2FCAeGC/y65Y+sIFyVZ8K3rzGPhetKNv9st5fnPhK5LxzjY9Ktw6e8xAksDcaKPAUO
qxK5M29YzI1ikclQ26sMedmkL4MXtnyFmyNq3eol64dYjPXMpkD/nLy7rQEB3T6MmNwXwg5jqSr2
eAWZo5db5vAvXSOUYv3UrEnH0QZS+wmaLolQnF9solWYHFhoTKftv21m7Ul7lJbr9KaJ1n+vVh1S
SWsRc1caKQgA3XIXzIV488L0I1QJUjWOdbOK/Spg6lVpJ+DJ4fKJ8i12EinPPiUTsxwzqTdbd9WA
Pz2vLAdhITenx2pZyt0u9ummmGrCT6jKQVz+z47bQG0r5p5u1HdIzFQPj7NDNqXhvc3/y4x16ycb
lJroe2MMkIaHm9GCqKEATQ/KHmqKzxNJZv9anK58KMe4qrdmSXZIPQsjURpUgzzJfREA1FESC+GN
k2MAPLPA13PwyXY8/zLd9J3sIZk/RR5tNYPVuhi7+X/F48wfcDRQQzvDtmE1NJXbqXzJTONNGyL2
kk4xZXYTYaIN8yj6GBaz4xSEYEJzTHUD790uPmrl/BhITsmCbvCyYPiSY9BEEf5o0oX8mQoPd6QY
hnFJEqCMVU1aNZIke7aCKPk1MTvO+/PMFqUZny8DQX9SjmuRA2Yy9EusRkwOMgvZhcWKLz6lhagk
UnwXzbIhxVsLa26XALsLzuWnjKdbvH5xBukYUbDM4uJ/cWaKjRVq//pgXY+viKXeQk8ozVFvpgsJ
V7RGV0a18cF3ODHCO4MCZ96pKoZgKCbs3L7VWcS4K0l7bpeSpCADIH3h0LuHEjZv36vEt4+Kpwew
nQmFH7AR/+a1GUNNxoY6YUBzn43bGPG5pWmrn/3ZK7qXT+BFVvDf5RgmM2V+WfBRG73K6xmF1Vgl
jZBykZxgNkb+mxH9PlOemB5tfGuRa43idy3EyxszIsS3kNrYtespkR7ToURngVrR1ePzUIEfLNC/
Va8pYNbpjsgR7gxOLQOFpxtv+AGsoicP4tVkya8wXOTOyLatn26+DKGLNTijanegFAP0CHvOr2s9
/8WsgVWPvjS8HANZOLJiXnZEBMjv9bYoCiw8p5AUHvBVFv2yjlbJKeV0NPnOudwo5ZzW7AyIAjZ5
C07xUHJg4pA8f4i8/V/etAHLHvXmcfnXXzI/UD6gnkIQemL3y8IDzyBxmebzKi6dXhJxmbT1Sxon
XIpiUaUgDjN/ItWgo9l14JpCugOnxisR9YSfsmUz+wToUztbwbtjc1KtFexfE68Sf+LV5Hj3kgo4
QNC7iw91BcgO6EwWDrww9sWa8GuaebpfYESVq48VXApkHRZNe7AM4NjDPRXax32bzqF/uYa/1iYl
MLB7PqD8pqGs3jdeF/I93mS5xGSow4Wg1L1+V2h0CL2ynH9QGrQZY9rj3RQN59CPecyqCNCVqxlK
8QQj+GEWzW66v7AZ6XIW3vuw+iy2J0oMfgH5/TbYVq2q50fZEySQ+X0VhAH6hunEZENpM4QW29qm
63790aMR/sGpSXGEJAWingN+NSkob9082pqmGZxSfe1aKVdGI49udqf2ZvixH7Q8HhGXxWIENgTG
hhJhXmTxGgT5AsRoBQYP5i79UqGqsyydo9juptpXtFSa85R3MFqehb0lKuvZdZ9AyeBgIJbh2zZy
7BuKqJXF4aLngtOQr3E5m1sRhEp5oDn12RY/TbHhlvGgkQ1iurZ2trG+HD8q17B690HYFfQ+55s1
LawKaFzerD5PjgXxNze+Ku7oyeik3siehnUwJxcsNcW0Cs+a/BbmjX1d8CnwTReD3QrGlCvqfZRs
lqUEwwaMrz2sT90DAv8QCtLIVUDnsKtHWYQswi9s67RmtH7d/j2go2v53EAgC8A7b8GBTUoWRLur
gUBxuis57mG2crxrJrzUEBzmEgjNAlZ580yr1mlSavtEtTfnDQvHYyXCZHpIIIxODrXTKJ7rga+Z
XWkZNQ7W0wzqGcXcPsDp01ocR40a1ciHJBhwRENaz9xbLwqZi3RWHHPckE3IBHTDcwHi+B10IQ19
Fv+lMfNmttk28I4Lt8f0kLg2n0wpJPfWimqyzO34D40RAJe/TgQNzBOVQnnYYecNIkmty6UoAjYb
g2LnR+x/lv/5+1uep8vlPuwpkMWOdfs1p1Gjb0grFhTgjELKLFcwEKhm7Eh6WwSiEjpPaRk0PWTD
Uy6YYcEd+0UBYDlSUdrCMZwevUsBskrQG9LwrIkkftSAgisHU29/QcUb/XH/gU3H8XjNLkb5I61G
+xs7VZsWmYZJXOKtUJqxVYctcd4JVO+7Ppy9k4ZdQX9vdOm2ghM3Yr0736dFy0CapXqUo3xwSKXH
E/hOFMIrXZ88MkHuWdkPrVjM9twECi5Tr41ntAKLGmkT7+HnYRXjy8+1nxx5CCYl3dWxlm27ympC
7iGs97Qt/cf51f29OQv+zFbK0z74zqw2R0OtjEyCD2qe/pXQisvnM5eFEvCBIzuFzTYE2P9XD9kz
69atYvl7BlQ4MTUWhvM7Tm7La4x1YqmX00s30yDqS4KkUBlOKVOadVFPsyNA3qn5IGv/5GkMKiSY
rxOf+hlm0Kfnj1olsOkcuzxIO0HmVphJavZaXTROMvcmxbhZGXaETbMsOb+X4MT7TxM7q+tvbxNq
4bCp/XyEZ2g0syq3xn6DbThBlngbN1ClKo/b2kF18XkvyUsL7aVaywOegp+7vffIrfkD3+L2790n
J20w6qVvZZTXX93EHbF/zwHDFdOMsYSDftDfMay62ycNHHzGDqjcSwjBeL2n+Td+TODrZu/eVTwX
8BKiHZRTG6cYZjMWVd3fa7UqlrnXbdMsNaeEMOzM9zOidXiPYjxI0g/UTnQdjAkDi43jN/ZBVQ+9
vkwuWlyfQw3XxwKWnioUsPxgZ49FJIQLfFt1+egXg3sig1FO5IS7q6mDlS4mx2cdcqKJfwKbcT+k
jOjtq2Ee03Ho2uzqyjgWnYIS8ioxkYOZTGFX1d9O6+cEYYtMuj1kORxi63oqDB9tj7nXODQDe1nq
eAcoTTEIAhL0OXYKCJfqiwStMUZ/2Q83kCM1WY/mXudn1lsiFb+m7GrukXk5k3bV4/ZCOIUjkSIx
CkL2apXkRBhNV+TBQfNjAPNezbbXc0bxI0OSWXc6xtD+ZH1gu7S4yCUhrxxnGTkiGKk4mp5JmDJx
/w7Rdcrtk+/+xBYlDSvbimd5yD9011xoOsKSS+15llnsOBMtYuGJlqdiuUcT4vS7OCL0MED9GnuJ
qivjvavnTz8flSjYesZ5zMbUg5wmz8bHIWE+4N7kYwOu0Z/Wt3b/0mDKCZdEGT8ipcaCsQI1gwMp
oggQDycUobrz8UZX/mhCyJoNkyrWytAAYOmVISKhhilUAOhfTzjPLDbcf24wStXIUYYaQN6AN7nC
uZ9rzj7igzE8zh1pc2FY2f3XUwBCjspnuVPx3NOiaRsyKCJRaIyYR+IXz1tBSaQljVmtHqBKtN7W
hv0ZJn8TFxYgd8KSoYYk5R7JnPNkdl8o7fSv9CXTnAPcuClTpB0GV/5w7gRwjCgZPx1CDH2CCVa7
Y0JG9qGZkh9e+bscIgTn8VCcqXJYGqeQcjYkMwx+pDNDGLOTlidJ7Hx2aSQR5rGOk3g61kqval+o
8ANWi1vzyGKNXn5szWyMUob51gp4FUSdqoZgmaouUOQugvJq0JJa5RXnce8fA//BtD6TuedvZ3dV
PTRLsiEUNQLb2GUm9inXsRwRwx2dpcXtvcc5RJ9b5NU2TB1yrtOEDziSSKJ0CDFSKM70mXSfx06b
WPDg1oGTuJy3+eYmSys98EyZbiyEuJb14FR5GPhFUtS73IDevNQiiwA4dRn2EYS0lC3KAJjJNvuu
H6+0zWD933CH3h+Hlg03BfpEtFAQZQAtn+kabU/pE9VZs0Xuacx+GERKeQaBp+Iq6wjUPVdG5ixM
S5sb/+Oppa5jJ0wULSuFA5nlsAKeIEu7rDxIopJRloTkJet90kJbpwrmf90cmM3jMp3mw5AjI6B5
nRJolMf8RnOmhsLpY2DUj7L/bxj6yJQ7UeCpMqgQhCqCBuVJWr3+AaqC5+yRTuAY+KEAiLfYDCJ8
xluLK3174vsAer6m8CPTGIICwcRcveBgsOKxPbNoKlYw3cIRDQXMZrn7TplR3sBKoHfzx4s2WLEV
hNhWmCdOjWrYFSoOBvPAXtbb9PUo2KydQ2DO1jF1iw6cWFroQJmLTiePw2nT+cnD3jchKlu31yb9
KhdWLN8oUH0dDU2Ro7wJPr/brLc0H6i/vBGRdcf7/wU1UXa3qTlG+n736Na25scEkt4UV4pLoHsD
29Bj4zxu+Q1ezGMn47o1+jzhPYaqT9q/9g7nRrWBVFefui5NL44763kT3GBawM1DY45HvdwJ9+hJ
1O7p/ZQjfOAMG3gI+LBYhqGqVnYiTtxx0MsmH8vxVdad09QuP6wCvogOStPtvSb17RBzCDmQCfR3
LtI0yjfbVT92pI+SFmzTgTdpxk/SjPP81X1l/V4Wn7e6WQVkZxe+SEkOiQYjou40xA2H1dO+8wCk
AWm6LyYtm2YNLaSeOMYJcgIgHY6HZM56n0LSjVvgIjYfLu/QON8pvfV5aE5RYmGNSbr5L5MEU7EX
TOkYaP6cVSIekRCgtUqfTzkHzGfybHJjlGB6bJSwgNqqGAbADiMA840xgPBaaCHL7W2ciSf/wnlw
ioU2qVMKTmQx3JjKwB3Be17nkShpoLpRf+oJvfFPt/1y38heGRmDmkJ7DvR49P4Az1IW6HTT45Y5
Z5ckHrigjaUJV2D5MW4P3eaxpqk3HX40F9Q/t2dd/YM8bn0R6g2XmhsLgX2mVyCJ4Hc885O1vNXO
40sw4JotDV/kK+qYLFOASJTFcC1/JsnVHakTCphEWBqtopBG/Mm0gYsx64GyHuMiNeKEFIzocaYm
0QXYrJ4HDDlog6dqFhWZ/QL+11WR19f0re/qhXKWVps+gLospS0/8He02HXRdviIRxtYMGUX2JcR
SFlN34ePTs5Au6FLcW4La5RvGec6+uC+EwI9F2Kq17a/idI28f5MQnEgOKZfdtFCvPai4uYZ0VU+
cZpEaOzjmsj9lwYSgJd8PPHMTCsZ+p0W8HqfSv3s1bNRoUDit+QdbJbNsIgLoj5fugdL3KcNF3E5
UH31qPQzPgm4P7OdcNgh4utyWwTkwuVeFDLPth/Ujghn6y+yVNtsbAfbAgzGH9arRIAXGAvaDp81
Z73j/xZI6sqZRsdkls1kuD1IOht6SsOYc6V4vRPsIiXxGfUvw9V6xUx2FrSCKdk/s40gHilmuPxb
Nc8rG+KSP+Uk2wqlnNnLEZJ3DtqbG+jNhg9h+udSJ7Jp9BtF/wqn72K8LLRvYI03eEz2twLSPWkm
Ct06OpKP6AZYdGNBqceCfGbaqH8WhxRv/j2nr/+Q6o4GbrmpkOPB/koTIyXP/ijsNhGBUXKW/nZE
KqK6E8eEpOioqK6WlUkuTFAtnBEXo3XqktVSO7iIbAxEIyfCi1J94lT55L3ndjkIZBt6SycLEmCD
edulWV6eW6mTwcqfHq/anru4TpEjc86v2u76V1WdeOlDjYqoWBZs0/9f4AD5Vf/whzfyZVfMm+dP
9NiwSUkfGz96fQWdFIlIE0/1U6p1YwCTTsb6e6I64jpbWg4qbVofQMculKuy5vKL/KYxDzHlXpzv
7KSQvnXGItH5+KjUPFAr9kIkt0qTQghQI87JZXcmNaMJgLNcQ0qH+hk8izYtiA2FoCwOfhLj+mBL
brL3EQ4Yr1XL8QiX0zVcw2yZ9lJznjD6Q3aIAHBKErwomJzNh7twn8qy/1MAqEk0NvrzpJEyYQlC
E0TAawbMCTK1rVvQbmYE3HSq5Fy6SZQI9fj7a07mTUD2sQKYGYYbqqFezoXqceWkPudEczmOMXkN
JO/HfajKEGe76dbdwuAyHvt+MXLmIOctmNAnFZyuDW70QhTttytpgg7pUc7nv3vKwpHhp29C9ODE
4IUctgkZezdv5KyYA/rTurQ25JwP7FYX3FnxzD914Bqjet1gzytd/sNYNJvRtO6BRT3jrPQSc6p7
JiqxTBCaI6M8IWvM697795SHP4axWGOFn0AQDQXloMYFr5l8T1nPuz6yPyYqdQXzKZLdGPlEMiRH
4lw5FSDvbejuLrHBNkcW9IAtidIIuWR4yxPSAQHA/e8fIrC5/9/+9jzwOnhJeK7BcNCEDbcMg36U
DJtbzg1+Hqg57gr781bniFKkS9/VKbdFHA3vTcyQR029NE25dDGl4GOAdBml8CO/ezmuuBs+CBp7
ZawptZY46tqArlHPexpuNw8mVI7IdTEcQNMjKs2DEa7WU9UTfxvGo0gVanPYwShq9aQ8Bhh6FdtZ
by77VCYEsCDvxUtNxSQ6YVbJIVxa8SeaTp1d/uNHaI7DBMbMeLz9Ih6ykcVnh4SA63ydkGg1vaqE
jn4jWaoAiIN/PWmonN07qc5HVvr4MuCN1c4APu/Jn+wqL9ehqvaFox4n9ixu1zWng+K0w/VDM44/
d2OCcWLjvWZTEvxf5V/gSod3zGOuUJ1peHNTJ/VMwB5UwAm0zwwC4J+3e3g4Gp+tRCLMc2aPIXTH
IwhuQeqWJapNjpfNGViGDgo3brR3P1dqTlhJeBg06wx25DSPReGTJNPEU2cnBdrVVFcobvv1EjWA
U88HELeyXq370nZvtChAB2YVqmNmnl3MYXunHk3hhNz9D7a1cQDYi0qP30bLzBHE/zxrgdAY002u
TPSSsgUAW43GUyhY8opSnGcRElS+qPvtRg/foRJtOyM4F7FTP9cfFXdJLOJ3Y55sOITVKGrPI52j
CarSACZolMxvcA2pWdRM3mquNnD5f3jm7+afQyz+NnKakeTw1hcymb7x41KHiPOGa9FU4cbGTojj
F2K9qPdFmPi2xQGZbkJBf+hGmhbZqwsVcFoIQNoNA4nY0DBcqzPRQu6LT3/XN3Qjtewdnmz5F59W
CLYQyh8gfK17a5t43ie18NqZUzVFcgTaw14jL4fiXQH1Qgwhl3CZB/54zcgqYYBVCX9fQCBIZKAP
5353/nRntto78bSdyPUCull3EiHOxcIwEaybnwk5E7m0PED3TJ6wGpvvbSCSUBPRp9KKOvelCuRH
K0009GjJCDe3m40ytmcfU9Gx3crkPYjIh79rjip2L090JnFzk1n/Her5vl5bOAtlHmWmKx8+fq5Z
UAK4THUvLAfvhMJyaVGqbqZ1Oz84D8O+jD52OS/MK8rk5AhFX8/O/gRD+BFV6NvzWK6OLd5ckCaL
IhzOPOwp3UAgJB1Yn2Hb4xKAs3x32lCCAM3QJPoJj4WCKzlGnTCUPNtDHuz9CD29p+yCFX8lppFt
5ajsbNhToTB2lyXcgkY6QKj8pdHljwNbpAnAem9gSO9GbYOfzxI3BdiI/W5qQHsHTn34QrI6Eiz0
b3TL8JuAc1NZqEXutHfJ9KKiHv6uQpPK3cnNYL837TKXbBQ5Fe6Ts1toRzhIkm7awI1/ysheOb60
Fk9646NCsXiVw98Eds1VCpMR4VmInyGLEPz7liDIHsj2WDmJ5+zCuI6EgqEmOpnqGar0w298Vbp4
L/x0p5PWjxv4eNiD1VvY4HQ51h7Uy2VYrlTH6nGvTZs/Z4IUPb57vZcvmBw9Iq48i0zWqfFnivLK
lxiQocg7X7cW0q00bpg6/7KjAFzLMxhMMcKqfOfPFDwiYkO2tFkBz+quEf2FDxxikQYvW6p+JoZC
cNaCruSd1WRJ+YZnXwFLVPMnmou6GjTGsVRtLEuBO9FLn+vMpqbuMyS0jPba0Ez2IxyWz/BtnMeS
NM4Z4P0rzTsXyUqxQBNwwa11m55zRYkr8eApTLIHQn1T3TVpbYY6fvRDOAkV5zQWz2hx48v92xUG
Lc6kyVt1HMBBcLT+B32sHsqde3/JGdxbWH7tEDrpFmGhN4rBbxg+1aF0J9Wxp+lJizYgQLbfwBUt
/0YJ/1NTQxhWo354QRZ/T8aotZKBz2RY2IphawUBXP1ssctMrE3JuotN8dNYzvUHI+kupBOfURMP
vng9GyCRC5OJIju7r5UCVUXnEMLOcBo8ZAC2K3teeCa1cbwNHCAO9z9s/fSHhh2Ag80v6OBDCj1H
ps6MO80MBQq9703iSZpsx6cDw6pQ0Q6jBgfGYdQ/aCbU+rbQYFi1AhzBklb6zcQOvdm4Vz60vgHA
VxPUkHFQ8QPvP/VSv7XxF25cCfgFe2SXigeK2WEZPWpOXjHcNNXdjOkcy7+/zCc6w1Tc+HnVkqra
zdbeZdilhKub6+U83zHW5dcvvoP/pz2l3IsK/MWpBeIL/qiNIZesJij99tSmuSmMXCwPYQCBGVc0
hweeFf+tT7ZtSMkIZKHBvlr7UW9Eb8EJY05FQS4b5qEfRd2ai5spvlaspgrX0cpe8zq36TKVzJLg
jsWB95+S7dOy1eKfcdPhVtAKuxiySAlKq7kfvu+P6BoQUqfjvncHNl5kSelTbTOTSMUsI3T1qVB8
ljcdLbpQJiIMRDjxVuGIPOWhGZijGWFKg6J6cOOilTK8LaJAGbpSf3jISuhsGJR+Xg5Xy+WPz9Ck
PpO2KAaPe2BxKADepsD5TzLDIRIqE9jKpl6ZAy6wwFPvl4qIkPro2d5ibPUPS5rn3YG4aGoule+O
17XNzRmQmtH/+2K+DEVCgzqDdeocn1gUnvZIjx/FQrixw4P75zbF4aKu5tqBMNg3E7+3iCzSfnWk
Dnm3yc231uJJcZr6soAPLnyQ8xcNNIz/4rtM3FIp6jQViuO6ZAxk5a76RSuHOdxGVicxxLTlgSMh
OWMsVgpyQM7HWST9QQf9mmjqfeWUY23WI+AdshpGhG2INWdOVqPdQy8T0rxpXGVYNkReBodPd7G6
POmauT4dMXRMuBIOHhzLslLiWJ3NZYhnC0KewVsIn9RAp13SErRN8/FlCwkryzi4f+A2wdv0TSv1
P8V23zTfUUH//6seI8Y2qHSejOPcBFWGbWhjgKjOhsv8K6UFQ0gM6hQR2gKcgU8hCfr1LAIVEw7F
0WzcWEVa3sYTxM0P9b0rEw4ZA8A605YPqG10JRiLIVnD8sh+4/sOwWmSnVH5gJw+3C6HfIDmWz4t
9lxcR4v00NZj1IZJ2eU+dZIkSfG7L7ZrvtEO7UENSWUJ//zmE0OpPMlQysIJwEJ63A5HSiyWZnNs
z7KWofoqMByCd3e+jmuvpuUBnqTfN9hluKWA0Qd2jabqEZk+lsXCIn8YbrZJKgYlkgiFLrk9xFye
fhF+ZJQp1+o7MlwvgQFQi6PGA7Srjqpu6Ab/gj5EKkUTXjRhjNRA6BY3P17dCoHdFjH+oUhWYPe7
kstKknLGwFmKC2CifCYh6IkyiigXuZwO3YLzncXbE0eFCbAM7ktrh78J2C0/e7Na3yD/8nPTi/BY
Hd21BxC+n/lhg7ceBLqYtzR9k2s23FuDcpIK/1pipWCWxz2ND1SQ7WcbsGeGWPr8HT2qxbzBkZ4S
sJaj8XXusgQ3bHGrf2yGGXJqzJRQgKyktwE1G5MmsYVEWxyJ2EU8XUNtbF1hzI8X0kxQAZDQfD3m
9EstM8r6/SGwPFJJZZtNeuqDrZ5kkekaFc/sOOa6DZQ8Opsdg6/Y4eQrjroaY3nxHQBvlDkwxNql
3++SCBrqHJoxn+iI28zm1yaWNGKXzpvkHAxzoeACvlrQdhUsqmadAiFGBrrge3ARVRV3n5Q4jehN
YS8lsPoMct0qP+VIdkiDlI4lzUxEdQCBzKpmQ4AWQJgJ4wI7UgBK6IF71u7FKSsjBjqup1d7h/mJ
TqbQBjbEdZ6uwYzvqm+mGJsQcIkJqKwIG+uGfabPXhlVtB7FdOAjgBKMDFm+wshuAkvWTXTbOOy8
F9c3aj4UKk2b1Vx0OoaC70vv8iU6DJl/tBVzotORdFVQjqfi5MZO7BUiSU2ahbl7fWFaDmnS/AFe
9ImR/0fjT8IDzfgLTTwJfByTximHoaqi4H0ijUOwv4Itu0SKjHSd8AYfpgRUuxAvDDIgcitj6kxU
9BJuV3CVFq1Jq7+O6r8TVjFcEKEbIDn8z5v/U2JtKhn48LuAY/+GjSfUZxUVr7PHl3TiYV3p4WAn
CG+K/SP9qmEhbQWBf1yKnl14N7qpKXOQzwcIt7mamWAph31D4RSeDq04/lAiBNCQRn77/rmuJwTC
AfB2/jt3hH+lDjSet3C7uQFrhd5rY/4G9fIhWoYmMhmoNPYxCB3GZsr6fBL6WRYaskiswJ1sqdbW
d+3u+jeZlyDABCTQ41WU48n/FBBDgiFkBwPk8TDBk1rTRn5z3go+zpf91WMm99p2cJ4ts5s2WqT8
oz3bMlmFTtpAkonhJY8RMAdpfDop3/vxkPLqgPItNJEvl/IvpNzZOpKyA+VTG9MZNdvQS5kESzKD
7J8G3c/uLqOMCsRShLZQcYzApVraKMZzXEh3pG2J9DA/zb0r38sTaVa+J+mcRxH52c2naLLUmbBE
XZOfVVta1e7QsdntA349ixoYXQEHvXo3cIWWwhsqQmqeqXnRSHBwQNhOAEBN1kehpA4F7EoKzT7U
ELfgYr6fyYgf/0BxcCUmvQhvPFmOQ4v6+v+3HQqu6YlC96MpzmabjRjPHC7QKaZrThGnefPAIzyX
DzrLP/PKpZzRnP69GjMUx6XksF2TWhmHepgH7KekPKZA6u/7TYDFa+ofzzQQW8z1qunnuPNCOtAc
vWSb5AAmqlKiI3UEIV7hqR/pWIgZsIEhsGHNyKQV6WK8RRq1Bmhbmy+6/N2VpbgqkEeDA/P01gC4
0/3U/bFRg6lb7W0mvTyQPEitHApb9PAXVtom161YkY3frqnryNZZfm0XoBEGfWssLdHMPJZtiZem
Od1+nEUvZ/XcvX7jaTcTZCdpcXAQhOjusGjW9nDvXrsewfcMhbM7rl1C0fMjLIgEcdujDUu/KvvA
ZWaazg/QkdJPArukH4/OjgjQ1Fl5eiZY9FVAodrdw0rU9BDnpvI/NZUlEe7RI1mM2kGUVfCctz0S
i5+jOZmuTveJq8vcuI0Lacx5zgB3BhQFQWBE7izIZPTGUWkjOWnu9GsnpnQkYz+b/hkEUIcTcSLr
pPoAF7rf5S+DWZDCE/sLyKWEqEfHE3pk/jp0O+gPy4T7S2fUMoBc7DOb3Tvcu9On0yvfU6XUFlz3
sin4+ie21K3bWqfDrJAtVz4zyhFDKo363dEC0HSlgVq1JdefDfBFhFRRFT9z7FChfqxavKaifykZ
os0yy9RZY8E/qUfwJ/lDqS5JAJn01GEn1do4/ZcMocJB6CJa/EL0WSAlew4VPTlXH1hiOoQkwA5c
iySARq3eFiesBs7MZ+O+qruy6jXU9JVuY0Q7YFKAdZ3Caf9x+uoszJEx/KjjO1YrEUS0mzW1WBMv
7vXh0JiegH14EKB3QYYzeF8E3Bo4noP+6iPdo4wZ0T07xWmnOcCK+PTHGRFn8thDzZGDwFQnUI0l
ZrlFY708HDiQ/27TQB36aoE/4rTGe13EP5qNML2vJkvPgOzCdB1Q3p5PyBfZ/4LVaVKBk7kg5/yp
vWZCGBh0riYoQWdGa6srEkwu7cDeZ2OokXQ5HmNy+nXI+HmgHL2Eyy7OMumFXY6OH/+EclmG1+cw
38nbCALRLOaeCRxs3l91+yxvomfJT3Ad914lfPo8zmSpqVdCbOZKb1esTE7nNK0DcnD2/xBPVvck
5ibx7XNnF/WkojgIBbOBqX6fpThzp91LPTY61ZtojBq1EFoNx/TDodZ6rOrbwH4mTmpBy4PNkozQ
0lZdtjobfgpgqfYf/o5+c5UIpn9sRMSSA763D/4dhKwb3FGisw16UWsIPel3wHHtsg00E06iXj0X
oPq4zM3brM+i4qx+l6/Dw3fvQ5kNhaFD7QcY8mxB+5x/LwCGX5ypLcW7Z4+YbURWg9vB7n5NhbFk
5ZB231KG+8syyo4GnhYWn+rFlkyyOiXTUgiGgaUQF30ynqYD25ZL7wjaXPedkKgpw4H/sTz4IRwT
3aQcp17X4wZxHLwfZ+WR9ADPYMXSZSK5FVzy4oR+lzK914KKvIETsdlv8RQ31IxMUcFOn/sCrYvi
JF0QO96fUxH/lT4gG1eJxu2uNdQLoyMY2MQpz3Ynwmza6r2IipxD8Jl1Eazi4i1Ghv1eOd/rYVY6
yl5HWQECOI38gMeQdR3EyLyM66/TRQ6P0bTgzOepe10CkSRK+HY3RWxmiWdFASfl7tDS3pyevJhG
nBOxUiY4CxVr8RR7xBuW32AJk8YEaogRS1EzipVrl4TPrHipVYdSUGEEVCJLN7kyWgHVy6msBarZ
9sSyroXTis6dJE6wuWmc0z6R4Vv2IMm/2zljhDcZR4O6ReXavNCGJEpl7dRnWt8rgh2iU+zcKw6d
xZGFLIgFTIlf7LzxDeQ7vTJydYgfxWSQ1qw++P0YVyAycSX21/W1EBZrq8MhoevgmY/P+jx2Mw8l
G7KTAFEDDaW2CjA5/ImNTZFyISLIYEnYd9R4aCiAHkiwpcxtiqvKcwskDCxoP7SCiUOZU95xgEwN
90MfYvsJLa+2D+zuzDoltOottnf92YsmbljwZqXAZ8r8AQGBBZ/eUtWlLlTthQpUUkrdovRBYm/y
TBKG+ox33m+mRYP53YQAm29I70Nz252VhZ01/1M8dtTqt+n08IVV5N9TcgGydawADNoftBFkMAdt
y/KS2/dglCnkzJT3Fp3uLi5sRhF+EyB/0L7+Ti9kvlVLMxNMcGjo2EVeqsMbiuL66QtRFZFRImNu
fuokHODKm3B3BwMbcz80+mSqGxdHizb/A86G4c22jrWFliVPtTkH2CUH8K37Z6jm/6de8j2R2rU9
MulxMFIV8u3AG5Jdk81b8OwiO4YOdAPE3FHf1Ch0XXnF5KABoU0i22rAZq9zzIsyJQFqohUzkg+Z
XNY+oEFTGRg0wKyUuXBvWRvitn9yWHZ65iAtL7O5ynKy0vupaLN/cm6HF2JPOfpzxL7Y/rplpAYy
FtFjSeHhnPfkSl12GnMmOWPAV7B8r0l0jl1coEOmULkHvazIa0i1GPf6DCIHoPm6/kjZaeD4KGXS
CoxdFtGaMCn0e/5Bhz6fEFT212Q/T6bMx1jdrs378BDDgnofNQOLXLj1wBpsbNS5icfIfyo9mrlJ
zzDMyBC1M4G1pfFbm6/bu7eVDWNSP2F7mzlyjvVhTWh3IrN45jtktFw5f+qxGH1bzrb3WDqz17Ki
J5wGYRWHrAVr9vl0lpwtKqbUiReeaulnRkoC9PYa0hT6/oVbZ3hf4IsUt8nudXVH0oClbKd27CYl
mbN1wtrKX27kVzH3vi7SuDdi73CzoagURPxqGbipYwC+Wn0Ntp+7XhyHwMOgsEUSEVxlaJXvDSfN
lEfp1jyAWZHUBeCviw2CARzqpyT8oyORbBPZkv0lWCBawCmp2LHi7+AtUNIiYH8grAua3uyClLwh
uV0LPTNhXKM8Va5Vru40L6AHXXW3a74GieiIpCdqBULohpKx6r7AN2IqJYYd+aBcracaAhRWxovS
Ic71TXn1iHR69bIOK5jR7cjMUD/48VD7vnFjV1CUA/2aNwOKGonK/jjZyEW17JLLY83OqbOzZwdQ
KfaQUbl+r6VxPc8W9Bt8Nk3aCRrzmvlacx+lp8fvK2NShXDuvvvBt7F+lsEtRnyAxrM8O8bmt1Ra
HOMW3ZTcEQdvGfEFu8TJekJape559lWN6kunAnzYuIDQOFPPyADZy/YRSo9JPUZy8o45rmG7tNlh
8+5Wxig3sm/el0WV1OxwAikhpLDMGeBml+7iHR0b21k1fn0natJO2d58wDoY0GeTBbn8QzGSAiBT
5e/xAcSEP7eUB5Ck9U226ikUDcd2sBSTVfr8z2nVBLYlHBaNm7vDB1E33crGE9/sZnI7jPNfsJCT
fQDSo2wrsBZFyYdYJ+ysN3zpAU07UWkFQYAmf2LEN36iAb8GzUZxQoxoDZhR9O9YpTfnbMN7ZW6b
iqaKI6/IxiffgDO5NUG+BEvA7+Pxj9IvCrqMUp+mlXBPgEI1jWGglCg4Pm95E0ZO7lfMkzhdvnsw
rGIlsza6PA97tfe7slOVuoYyiYUW+kB5Zu9GerQ2/0n8TAm9bTvcN+bxAjgdjJaBolbBfzitVQ1F
XE6I+JVHDYfdYhqiV4FJoPp39DCks8BmgziTptS7DGCoOfl7H+uvXgPGM6BfVu/+U90+omB0FdPL
x+x1VWKN8qiEFwtV1GlvpYYRccKfR/NHh5v40gUb66Ta+D8xJ1LoxPkab/xYA0gJkXdHJvmIxdoB
3XqVGnpLaSa0WhRBjkVVuhXvTkIobuVDpmAUYF8hlqi+XaGPW+ajAKFWPs0M7usYlotLd/EdiGQC
S5dlJf0mH2jotVmmP6SPoAGA2hji8HzQ/OxQN/kFMoDB5HKJNt0yDFGIqXPk8sVyg6C3ndmUH2sB
69zH+sTI8+B8y12oXXmSPm/84wqXOkN5jZNo8Pmri2Nr70HxVqK4AOAw35ovIMFLRLARmpY7EIF7
IE6bw8bN06S6+EPLeYMVCpsdR8yVHPRcyh7QWWpDuMLXGap9T44TRUGMmPESfvwzv/OpWusctV53
WUB7DTLrhW1cc9JY5b5PU4sap/EugE5JulQqzVQiT4IAy1UyicOS/5krQZCslQQQOMDo8CUq6p7L
IU7TJZCLMTOiSJglYFlHOs3qqN9tp6wiKtjBbvXONmt5b+QLmx8OxoOn1WvA1EM55BPEoeaQ4F/a
7lcEBA+QiteMMxsbYVNqqJHb20ITeC3IERMLjqcxuA5BjXl8vyh8sQkH24r55fhHVeO8dwPXF4Pw
0S3fbCD8GI03mHD1oXn8/0v3P31pWwsp1EOZYINSYV5TVUmLUusekbdKlUANBhb90uwg3IfSB6ZV
msls6SPYQB5uQ5bTPBWh0Jeq3C70on6REpsMkgvGKIRN40vzo/UH3jDsong3sqGSdedw1sFeNMLl
mxIOhJ5+yFB8lvme2nSqlq/wW2pQHZRyB2T5OuY7dYIsNgXF3YBrawk9hv8tvtPeHXrQjAVDE5+2
OqXlB2t7QjHfv1OAJ4NcwwmVYggE1qlTjhy6gT+2ECcb7tnK8EXF9QGOjkuMnANVMK7u9r040m5x
sxIUr3w1gDVUrm7WOU3RCUJ162E2eS9DT86OgDyOOYH+9ufn62+hBwbCazBVDWQcNPPIVWBhlGKE
SDp4fEDMOct3vdw/somMyJ80JPkveXSBW5ysRDVr5c0mo7nSjXmRA97E9kZ6WKRPkyTd6FYByo4+
hjjRiYAMR0ANuzKWqiOYoC3KhuY0VMozDQM6vFiUnxaptoDac9CYexw7ozwtPJnNSnme1O62Pp9+
cvV7I9z6U2iN1mGze0tKIRvz8upRCW8riwHd32jZ1YDVW8uqTxGPB9pavIJHe2rhikdogVdJGdXz
9tgHs+sk3QzhnIG4zWZEmqmjI+RLpMobSVAg+koPkCbJWR1dZzCbQZ2eV2vEXfqDOFXGMHHifhPX
gyxhgW3bK2HeM3xFlJq7pUsw87kJ5TR5myCkA095NdtK/Fnv2XrGh0PtWa1iWfChIQhQm1VqX65o
c9cVD4q548WV5YcSkJV/ftQN08C0MuhPXNq+HYTY+Gm5BLdv8MdVMLvcL6qQF0JgjowBfis6BwlZ
kwmS0wUzeuNznTwf9sRg/tIbPM0JSYRUo/6FjmA5sxurNDe4JX2ENAH8dMJ7Kv9wB+XwcqmMEy7N
dD/Ac35qApN/2gLSlhjW75h1ruh1XGFzYEskvymfYenZjxp6XYZSNWW8ySDmNaLym31aPBGnskkx
RnAGSc8PvT8ywqW3M7vWJ9vAgZSjMcTovGAGM+PYYh3zQfuEStGwf59wQiehOOu8DMjK2IH9xlAB
zb/f+X9YjpFrOZQ0IjWJSnyTbBZs3IG9pVdlWsJSGJwTYZ6NdNRzwR/w81Ftwr+piJkpKAhcsYsp
+/5Y4WeCyRMBfJ4mMkATaIe+9yw2A1XWws9imFp4SOiINZHIoJcdPOl4AeWqbcHxkOn/O/+RXO9W
9vgfVHPKbcR5f/XWTRsl8oZ4xnWJPU5hUXb2lL2e7+MK0rUd3r59qpYNT0mEYYnN7oq4nScqQvKO
QLnDHSh/H3U0JT8dX5+4fpwWkuAS8xm7uheJx7w5lI/eNvpUQld/xyPAmVUCV8YQzk0lir7Gyoh+
/zX8/oPDKC75XcjeZerQmDmtEUpoo/1vDIK0jF57QvoGRAoyppORHWVoXWObqnRq9eTvIf/aIJcD
4WOH7dkQrOw+Gphw7WMd0S3gQufKaKGy6F/LRubMfxfD/Wlfz7M2jemHGSuK726EN4hNhbvi4AnG
/vdFTwhqEbFoQnvLVKZE/nzNwrP+E6GhTGAYEq/Wau03sabmF/VlbfQTcOCsJgn99DEOvsrLcEhm
flyItQxKhfQP8mmwXheYepCTPLEc0jiF6Zk+4TNU+J5PYwoTnPpUeMX0P0A0PtaofgGS/YIpv2jR
mdKlYMqU1mIh9IV1BAVA95YkGQ1DoIbKmgBAEnQDFkaDXTOIUzGN1f6iMw2ZNkgyHoH45hypD+dK
C9EtAIP9A3qFmvsGlSJxmzNorgaxZnW0lNQzCN/4oCmQ2tZNlnDr5yOI1xugj9f7HDlppsf8yJIz
hzW2xciF9YvcqYSKKN2l3p8D8TZUKRdb6lXHpOqu8U0qSmQvLEMgxcIv+L6gKeLHZzZyoSvDNa3r
wJbgZX5+jNk8zIcRs4m8+28rrerUi8Aq7qe+2IQEfExURzy07HlfnJJP9YbBl4RWyUEaKaSysJ+r
f309cuybr6eUUq9Rws/kDSGqH6QlO85zN36AjGKYe7gp1dggNIs7Yq5hHD8Ay+VqHs7YMdELM12G
+kwANdkvXKhDLXKujmhpbZ1m0js3XtZnzgXDVCv3v9EriHWMFly44CcmNZo0qnPGboz8zfBNzIyP
WmJ/f9Zjmhtiw7kxauahG8+5T6cxJsMn4FiQQoIIsSaTFnq5ALUUxwVXpFXqObLpW1T4G0fa8WaA
KH/kYOd/HAikBgnwnhRwf4s4Kbn4ToWXSl93Iy4CU4mDAoyrZiQbxm8f0efwaGUtge3AtIzEjcDB
GUnalSjTdbZZd9ovlCoRhPizTyyABJ1ydwZxDd4ZXpqzIXkDWmFhdMlKXO68166KWCuRfUvR1NX0
nYluzbbr+ahoRz9Lnem3eyOkuJMqxpqPSiPH6UvXeGnfNPVkfnsZtpHvXUe3THR1D89vb68FFLjZ
7dcE5V95F8L0VnV6+BuWaE3wGPQ4NEwWx9OPKONseDSYSKPLUEyh5wp8Oj5M6lEIBbjnKa6DVB2q
FAK7xvvTNSpG2hxLuswc9pse+uajVpu/C3nfrb93cddhA6Wr0A+AMGzYcDDzQ9Hj+rnwC8vMoJ/A
qIpWiD1esfOBV/tSFdTY+EGB6XYoQkhA/nNnHwgkgtJ9Etqsl9uy3U3eGEFpaUmm0fT+JCpdmpuc
1JhLK1lRQ77TF4DVYqz/hH2RdOdFSkqiwFif+WN7KZT6eupCqF00MVp32w3SAmObxDE3Mydp2X35
bBfRhEbd3iyPwN36XfBXWzKFWuaD0+c/jMr3q33jaaxHi8kioVi8uUHiDKD6QvAPav7T8Lp9Xze/
njEY0qZWOwbVf+5f0kod7SwHFZ7KLUKEAvU5MN3oMOS4BzojKavZm9jpUElRMy590bNWiEf2kqRg
sddzv+R+ivxrmcTPungrqPoYQ6L2hutzjYJ+QfUPPd19XHw2nSTWTMUfj9oayP6siICtooM6rTfv
z8OorGJvg5Oh8c+731VCd5b59AM43P3MKCURAeZENzHZKMqu5rtkislbWbdk76X69Pji+3mr9H2Z
Y773Jvb/ibmBUGYCBBa87icbcNLhZ2KbBncjgWdzjkIbpSZpmwaimqC0ZpIJ36aBypvbas7eoLbQ
nt1zwoWc/tJK4K9FCF22FhEKmnz3FEacnZGd0LFGfxDDR0+qKfNTUW6uy0o2fkxY6kVcfRC2uPQ2
Cj6ky8Gtvn0WPLu/3t0p1EHlBnNpUFlcOFoXRz6umuYlqYTN8C2TwYnUA3BubFqRwB6CPM931eFL
c25scyI+S9URLhgNgQdsSV6HHbyxsLB6eNJCG1Cj80i5dTNabot23Va+MIHTeKb/vGuk2hqAKYnD
KsdWqT22iWV1dVzd8xxVNHzBRX9ft6Q6DT7GBzVzJdcJ/CqBQ3lcTjQmuRhKX5Tjb1PIp2rjczun
Kz2YD+PJdUU8sXiNRqaXZveyiWpurRGHY5PKyW5QGbfTsWgw+FSKDvuPBGi10t9SPljZiZ5Wqzc9
htB7WQU9ygUhFwoA8ACyIOFL1ZpREUE1iXikw2ihoBUQ5cHVYfPHSpkxyiBFrwfy82lQklE3z8Ec
6Aarhvd7XrXo5Z9253+ccqEHoRFgCGmPUa/sBhNsreW816W7ToaZq6c8T6fnF0IO5HxEVcl93jlM
g8TcL6q2Wql85I86gVsPw/PLVOgSNtAs+qC6YYEXZc6dizEHL3Dx0JMFSp0xMalpn8uRP/VEYjme
bTS+AzY02paJvtY1wKdMsylBNSTuQOCw/hNBzXL4lc5u+9WFDWBP/ZyjI3wSKZN6tUxdVfh9pE/D
ZlVs4/AG7z3QgFmkNMPCqEHfqT/rx0T5+EaFyHIlIV6s5qF2z3MJdms98p0Y6aFErtelycplGgmj
qBvhiV+PzTNE6zf6ojGubyeJVBV4L+aU0L0ljv9djRtKHt6RP3gha3C0TTQAgovBa9uJ7cqhN6YP
LOJxV8tfy/8HjdBeR3Ka/Dh7ZUG6UYuUyJk4fVTY1tL/twsH3NORhZXrL6mIAbCG787Ua7eux8Ti
j4PZDzGW4KyvQd2wJu16udX1PDjt7W1iy7YIBJBOlhadRwtCA5VtUvfDfEKNsCuw0w8kBBQe700L
wwt+o5sASYsb8L+G3OzZkP8HfFuDgPEQENhlkzntY/u76Mv6pHmuBKXfmhFJP8nXCw2WxgeGlDwr
liBNSJ72YEAwc694qyX9pmgEAC6qijzByWb1lB3he9jllXVu3FXtVQ3miYluTkgsz/FnaUcLKRLR
KdGRJy5zZZEaAbrcxpyIw3y0LLacuhhKClYHR4VK4i7r8EumeE6wDgNwnDFPMwKKISiuKmHh6FrB
3SuqE/W7LXlXGpRSRWvhQ14w4iBbIzrHOND6kJK2rtemWLye3KpbVz+w5K+w937yT75tAgXlYlhC
ome+HJ+/Q28dnU++60OWJPbd3Iq2Jnhm8wTyzOOfpP1qFuPzPL2RBohIyNPFLcMRdbXscf59alGC
5H/yoG8NjnBHIHtJL3fsfmI135q/u4dqiLQYRqI7FhEXVX0qtiGVVYeBILmwIlxMM1OGq8WsBIWW
hZ5kX8e3emlKg5hr2Qmja3r4pSJtG3c4B4lddLijchXcPjw4lcWrHqv0XxZ95vz56j3lYGZBClBN
cSqjKdSwj8CM3z3ubw0/w05WVt0DpN4EwmFoe+1n+Vwj+6p+8AASq4lydE7BXhFja385L+lBgn5w
QCSxiY466yLD0W0qVpp8VoYx+kr/SLixhI+3bKSmsJkLBbjGYxHCtIGz2Vd3lynm4xOuu6gJTnl7
D0+n6bgJ428mN2gEIHxgBrcWwvVDJw9pfisVrntFxAodcmxvKLtcvvNRhOunqQtbEUtfz4nWPLjy
DqRRi5QiMM8Iny0DIk2zpJU75GMH1D6xyJREDLkeIDUTI20vEeMvMrMZhK45GTLNGijlFryuDexh
ncakaUmNHiwyg6wzop3by0J7WNUNS7eDcCI5Myjyw6ZbfEpcqGUHMd04qWe7/BsQ/0Pu4jjQ8iqs
wXINKSDgPhOb2ubbEyoP7owwPaIQlgZzHgtTktQuULH31gcJ+OFgLTXUhqaS4bq6OhSG/N0Iiy73
oSBclq+QM72UExKw+JsfQjHnYg0HlMVem1680FJl1pM38QNCnJnilL1XLiFZgXmRr0ySFb+RYPdz
J1LsG2ge8ukw4jYnLKLLqa+ZW9j9VbpeBz4Xmcwit8MjuInBcUP3oYbkTbd635AqTsejkZUm+ftU
2LCdlJEG0dLkN3RRB5TXXrdkvGz7gXLd4AsTkQLrCVsZ3R2lLMszskjMyKyZ2PDXy7W1vEDB8lOW
x064EqKLsHO3PukSAWz3ovVV6kfHkQ02cHvB/mgOXrcQP2UvLZCu0hWR9rInr1yGFSvTceHfkqzz
TSzccagXWhzKinqCTy/SHhZsMevPxwzCRD4BMyKmrmYtOqd+IhOREfkcAueGyku8FeRWNRAPDWPt
jaGIAWjWlmauKNCpvoCncLKvNRg2mITQrQ09eJqgChw4RqQIftH/sN7SXpZJbAxto8qgU71/y7Ln
aq4wZdVV4TmlxOFP5tbx3otai7XSJlJZ8FulinMpYQhUHqw+mNE+vIF9iJ1kMFp1otYDHnT7SQm8
4up2Hf4Qq0aE6prRzl+yFSJfNSjKuWEorrvZWnxr9DpClAQ8QB2kPfRLeLG89UbXtleZwLvVfLBi
iehqSu7PzHpcGg40QFyDwz9LjDLAbW4q1s/3zFf966LkyBE0HdXWYzVJdc+Nu5NHR7IWr2/+q0o3
w2Id8g6fd4K9fKHOJ6dZEagcs+F/iQA5M7aTjeGTZCR/uOonorb5CVekC53zFr6ymQK/8age2bRa
a/Y/5KcyhlJ7d0tDX+dBPkGxDJ36QD6YpUi0xQzYrDOSzalPQHxxCJ7qW9mM6WhAn3tzTMWDrvmz
2cld6pm49SPYdWGrMFvEOdGLMelHqh5rTNJ0p8U9AVtDQ0T2MkZDo258a9QLXwgPxT6xmW2xYROH
jh+K8ejklKnRgYcZ6ufyF2LbAx7jqsoBTD3EEKq6AC2HVeb2cBUNXDKuDEib+Szl4UbZkoKr+m9i
Uo/jAwhztnRI9ktL0ioFBSS9CH0nQfPdJBvtw9J0F9BTtBcIrZ98PQShi0KGEa8cS94cqMfh14IH
OCEWgO+YB+4W2WS5Ysd8gAXNPt5XHXY8dbFt8SDCjlhYjCmHSYJOJVwLr3tA4QlrL0y95txuwTz3
kdYvYzX5SYjk1fV6sfE6GhDB99xW5FP6xiby9iQ8dXxE7fOFD8CUCbVeFK5uD/PGvhFn5wW/LWdD
HTJmbUk1njN+scB1YaPdyEBLnicL7ccktjqsvmWi/LhoUvGwvv1DH5Fmxa6vq9QCqZbzHic+Cuds
Sw9MNOyR4YM5+SlIfSUsyrucENG6vTTcrT22KszNybE24O2hOVwI1QzzGNnoglmQhnhINrKBkbOE
qDmXYHijw1KiuZLkiclOPGSEpOfcxqNlopmaw9MD5wpuXOoNXN2P6cekECILzoCnlE2PNhi0UW5w
lBxCyO+6QNLCVk+/zExaPcZkTrVSZekRoInp8AJYAVivuOyIBnhztRLPf/s8eAHHuVNgQTwHcTe7
KTGJoitEu62lDUecBHyIdt/A9VhzvYL+95pgpQFLF9kylbV6tt/e7DLMCraQiQGDbHBBb/vr0r/J
w8rjm78arkRDWPYDlaUNIMFjwGhQVM3XdOnKa9av0NuwsAbAWbC8j5KX90ctHcOHnDeS4GbBv6Fr
YZnXa9bMnwmqrxEvQHWgfFrLl6cVcPQHrFtWECygQ6nwQOSOniMnF6aGQm3GG9eF8KBfjNs2UtMd
n3gB1aMmguI8CJnLYWiZvr7a1RnQoFu06MY1RD09efOckgAgxrjCSkHvTL/EWerorbK/AutxS9ww
VYrgKa79VUwtodTnpI71YLaKQXFeLXiVr6jpeUQXv6kNjAKYBOKRoqBKy/BanjWJhjHlifdOV8/H
E+ov2HmPmGVsJVCQosrV09DaEmnCd0PT2VSRqkuzaipowQ5nICaydSpELlZgtMzkeMN/i0+5k8ow
imQXL79z4a6tgEU6VyN03ZxlbZ0ZUy15H49tnmFoM5Flq2rDOhz+pQQVHGbpTLsKiSWaACFuZOFq
XYUyEJ5IQ6qxOAr93/cC97rRp4tGeKta8ZW6IYyCnoplNLyvt7hO4vFcGLGY/I5QpIbZBHw6VX/t
bZADy1OBVog3ZA9zeMjFVz149sq4QxLlsqWiKlPqp6x3+u2BEmhI24wutFjs7RGvd6TTFzi1PiNI
WWeJQjNPz6bD1+a4LirmV3ZglK7mXpSFY8kE+ETW3r5fu0BnbWoXnief59KHgnZhvciU8IW0hHr3
qKPsNnvL/arIjZuasZwIA4FTtXHLCIHinRrmxoLvBbwwImi1f/tmc7qMU8OMuWMOFa/VXH9nuvn4
REh+Ed0THdsWA95VV5I+63ulymWiUOaMpdOVqD1KO7sUzYIb9cFaKnZuC0lxc5+TozvrtvcpSuL9
vr/Q9tI51aIpKB99XUL9cFa+thBULSb3FV7xDGD4KVCSLJAKXZ4Y0f97WQ+yFOhJ00TKbjC0uzrT
dPK83+gxUuQMQfGyO0b3flUufcj5B7NTcUMxC43uiFq3pc3rIv/5AR1NamW5lkoNaDzKBWfEQsK+
DOrElOSdnn9to1D4syA/eAmMiM0lRIhotssD67rwxwFaV0l9c48KijwrRaggFQzOkNd2lcFQiQ67
eL5yB+j7dYKM6DtuLxRJ0zPQ6nY/9560CAYN5TGjalxOSXH9ekpIikwtY9P28J4Qlr7ILKxxanO/
Hu6+qQguvvpO4PJ3jsy9zAA63jZkPxdLXg4gQoFnzQgiP7rdTcjluIznr6xaxdiLoBOaxsOwvQlT
gnuE27/L86OC1IYESSEPISYFlY0n9v9nItSIaUvQRbeajj+pztAA9iD3YPbEtZvBFlOFRqqAc5g1
/6kWNJNE3F9Ri0lyRLsNUaUpenLzUBrp+XgvW4TMs2rkcV89eZqtEYQ9Qn82x/2GtbYMTx9Tlhb0
dEZtMxIFVPc+zDr34iwE/vEdSYF8y9gwv/j1NQWSTjhflBk/jzjmXtG0de2ojwhmTzcdUZeZdTiZ
KFad6+oQyzTGxgA3P90wMCmV4NUfKpMwQsR+msMWNRHuJ4nNWUb/OZIEKSQ+j6HvpFTEVzj6VvKS
atIYmgU/txLFpgNiZNM5Ea1V3Qty4tucBzHYTG517cuXlDE9uZfPKKhaHfGMy+oTgRvQPnN+Ex/8
hVRKmZcx0XponEfNC3mZQuGNA2rNkYs6stgr+cb0h9jM/A8AIXDqiIH7tSfrlBE87vruZEaMM/P5
ySo2N70pIxZ/b/jHFK+NClMGCWZJs+Pl0PQHq0rHbXdQLmKHQaER/DUrtdbMCy3Do1YgZXUEsxqG
6Zzm0UoA7ATuYVOcgTe7fkavs/lNUb0eHfi6X7BHZROqRiFiF3NOm8f58WYVf7bAchb+4nSKb5sS
U8+5hPkbqA3pt4gG4h0TyulpnpMJF4ozRZHy5QplTJ2bNJnm0xI6nPp6/b4LiAAS//PJmIE18I83
3XyUxKp6M4mm2hcmQqrZW/Yp8AQF1YReOpBGJ1ZWbWx5Y3D4RKIu7CTX7bPC/uFC53XcwR1xp6YU
bv0tAwoyZCCtUWtrEOj9m3LKO0qRrqELtQbrAtn94V9sEZ8t/IpxGOdUYdz9ESpRFKShslrhq9Tl
eaii41SfJvo6xrg/J1itJEcHPfccYKtVnYpIsuMM9Miwpya+LqzPFd9zgWdZzUKM6UG+EEhT+21I
faLhsbMNtIObCuQKRkydjGpH2nKIb9D+bHL6hSvyPUEf9ICLHB4jd89gusXBYWpsp+YabwzoYpZT
PY9gr48EEvMy/fBhNkM7qXKKQ0ALNBZGozOsL6aZJKvxO/H+31j8l1AuylxA5jAmRsaNhNK1XWtY
xe/7WCoL6mJQwP6v7PJClogSXbplcUy4IV4k4D8+5f7CcBTc/rEIwakRxilBi8nROARplCttRSeH
gi2OJQS2LZLjaMrBeSen1NIFCj/WXxEX8/xG/IIn7MCFvMeFNW1ZVnJWsaXMInr7wVJ6rfz3vlde
rf1JjcSJF/miJ3THtooZEl3Spmnje6wdgeBjUJ1lMlZnMb0p0Mp10Si6BSRKSDIApcJJ5MzVGJ6d
HcT09i/NNliQatC2yuOoWXxdqzlBbQdsuJFMTQkKtCd1REpXQoR0BglIJGssYxVNly7Mxs2/J7tc
+JuH49+NQfUKSI4fSK7anqrmxXcI6b8yNQf9KaZdXCfqv0XNco+8wzcFiFAgMuiOW5oxVux4ex8e
f6NCfJI2bVun+7U/QaI6I0grJIL8gU62hmcbBXEe4Zmf9Y1ptdjoiVcaWIRYBAIAooL0cS4UuXEU
tpfmIh/6jAEZoLhmCThnISU4qSOjyX3v2Y1Mx0x2B6nGZJTgh7v/CiHK/47L8vfUBYbZXmoeHDwu
Auh57ew6XyZncAnznaJKJReKBkmStr5nNGS7zEdFFWvN0attXw1Sc9DADj+Cy1o5mtC1i8UN16WC
jSw01xkV6u4ISZ/cDqG60RU1Jpp/EQulPYH/99Z0Kv7IDovGGAO+pdm9tFFDpy/13td6yzh+d3F9
lcCObT49RJiwu8UeGuv8ZiJh3aNmqk5komiXT/t6JjPp6VZWbrMSqyPFnpKYlNofSa0QfapikB66
Kzj5a9AYRuqxmfqQua9POExBtoTp+ShLmmpz8CZ2+zk6CR8ikdQ0uXcklOXOZdKpJVSqYRKPNMX/
3nB5qtpdplq7MsNNdjYsoaHg5sQDtEy0KSxbYjXNpXscFdcX6Te9fjpPsbiM9IJwWrYNKK+E7oeE
5aLW62hiBiRr9+lMV5PpSed9V2ZswiwZIlB5DrubHXaCd+JwpRsukYv3WYyHpCNZsj4nm1/n2a3z
o9L1Td8vMXVBXFPDYVZ0hlQMxw5xIsYrB6EXEFDIrFyCpi3Qk9A8p/1NlhBipYBB8AceMo6HmAhb
SdUrxspt7ryJRzccC6CeKLGnPOlZfzJljZresHAutaj0sxaT8gnB0O5AMJxh6ubGz5BPjlze//GS
pm8FliCCBvogSw6R+2jAzaZGFsFfAVdgUu0VmIEYBcEMz1y3LL4AWWrEol7M72ddaOEtfYWPNAnO
0AHvRwU8tYEXJW8rkTDCAwZISST92M35VFJvB0L3BlTfqVp4g/JTlKwg5jh0fcLKsfOjJre0KvS7
dilk/jm6aUt+PekI0oYSYFU9nCYvjRdEPq+djnvU/P+o2ADH70LJVo7VqIUpLORsFk9ViuwdCLBr
nOgM/A+/l72vDqptXPlDeQiTIALyUefQz/GFXfwHokEm5Txp+ZSetiYXUqLqoElox2Nqwh34CNyj
2hAwq6QIeHWdUJnmrET2KGbYkotqgz5ro19QSmX8DLzOiE5IwU36DM+tZV8pdyaNYJDjGaEnNUPG
lF3+cM9B9teKJ7q8s/kJQcbEOuuGZNGGKwlXCy1i2AaKyOLKhjwn97ZT/TvPbUJWNwVbVTqL9Yjr
lwRsc/Ev4LzRiSjvgG2eOm8fM6HVXumC7dS2j40IkOT3BFilVa3FES9DQmoY+85lR+ba00966JJG
urvPiKB+0UWNM+vVddDIG5Bcw4E8bOMK+JsZJRna0d7xh7gz5fo+7MB2ifzyj17XMbZG1D7Gt6Ky
XS+EYGA2xiMymZC8RnXd6wtOBeDRFE/tNCERboBrNy4sevdU85lBCfXBEbpAyglaHd86BzXjYioj
hGgQ3i0wxRD9JkyXTWrCGACcbSKmRiYBnU9mCuxZuNGlaSy6j0bkK21pxMBT8s+H2/K6xEudI8Li
+NllF8EqYVMybBLHP5lWPB5MAY+o0fLd7J8LlAhvOro4FqPnRVsOhOBJ627r3+Rt/rUBkqkIX4rn
jdxdvWJ6BVvfXPEVPY4HqHOMcj+jXDv3fNnzf/gWHJEHNyR/UW3zbrbA6wjJVivPHTUYvVs6ASuG
lsMr1fYh8yz4L2frLU/HQykr2meEzjwpnqSCB8btxvR/t/dqXVdEUCIjE1x5oHOtD8ROBq0gmg7j
+ljA/hXlJqxWc3XORlFj5lejTSLUBXXK7KeQsEFuPrgKuCsXl6WtyobWnsAdLST5NmD6R6eAmW/C
NSDG4btPKj8CRLL2Wy2cjY9ZXCglZy7/x3Hrw01ZSkVKvkNOl2j7xsa047JCrtK+kKomP8IJP+le
q0BhxB0rY1Jyd6dZlSY2+O6ai/lp7h/J1KE4aVipeYe/dbalTIGkINGsiZTyMdJ9Xrn0cNlS1nAP
qdxFRkP+qGMgvjy5O8s4jzFaiRU2ukY0U0+hKk7UdaMAI8Q2EnqKT2HMjIBZwo2ilve/q6jKrWiA
AWWwVTsKSpQJjLrsOTjxsY+E7FxmGRfYTMyB3uTOKHVAoDJqasQQuJ6+URdNihwoVZ1/lMEtZGSQ
xgjyqR11z7bZ+WnNHIsvXi1FkvTlJGVcZMkLAz/vcwA5KAAghRB8JyeT2e3NqdR7Dd3SDKrMyf7c
JqMYZ7DhPA1orJ9HHp3gGJRbwDfEg3v2WBRyCG31YKZb7n2RyRp4s4NxOq8A/ZIS1sZ6hJlUhdQM
18eMKxBY7q7c6k8asc/RuLmctEe/aHN/z0zRX41Nb5UlYfrV2w0exR0DKzl90Eb4kRM33Jnndd+f
DWNYjtMaUhBHsnRXuGPaMwsWsNl86lhky8rKTWc18iDmrbkjOZW0UQV+e41rhJk0HeX85zyAhL8e
Jo5k/yPl2uS1oyGJtmpqcPa49aZbxBnxLMU+MdvLWn8QPGF2+yjs8d4OgrRfZdhcgC2KxS5wI+rP
J5mx6CMofyeeShHyYYOj+zqBDaNo+I7qmLmk2ghuu3plKFywrbi6lozIXxQxcRIpWHZLYvCKm+CJ
zdhNK+/HZyrzbXdXwiD1csk3eI0s8634sfweLBXY2UbUHo/wsUiGnQ6fuE5xgjQfA/jXTpdy4J6F
MLf0tVMVpIq380ZdGo4ZawmNWu+MPjVKNODO0ss5BDMgc1YHakqMzimg8WMia2oC9T+lBgV8gd6o
C9u/vGvmNrc5RF1HlBZLlIJS/uHyU/eMbibg5FJ5Wfq0T3jXE6vQIjGgGwmQ1aabvH9VEZUWXBGO
EIW9R2a+kPcDik8z550RuQqSOLPUZVZD6qIjxxfQBeOJT8iyU1Pd2Z4o16LBwa1V0Vehia1oAnTq
V7irYnGFJ0BcRdHuhUO/EWbwnQMPlQyoTPhA0UC4wYMLeu0m8Z9d+p/8AcI7S0UXMdrBVnmLSzfW
/Gdc0ACu16NQME5vzkJUHSGk1yTNxodi8o7B72axYcjHScduVMe0gutQDY8pzRLuGkk6ffgB7s1o
rmU+StonJa9WYogYv1ehzzClCIPAAAcD/fVb/hsz/9jx7eALl4iDJbTxdjaGv5dCw7FKmtHFSMi9
cov0CSlEUUwIuCUEzUXMy1woUVzMzouqkKNpmhXokUifHpZ+BP17QkyUp95kBntoOXA5kBRUTans
/uVK+rEt6lkAy1hyRwGXLRsLnBGvKHT2h1Ff60pECP0Y531FShowRgXKWwpbneCt4fizbXC156b/
Kk5Y9RoLAhM+kg4WqRNAvq8c4MaqyxtYvjWbVsGi7T8sPq44vAms5Jzto04e+HptCF7MztA7V+HQ
60y6dKV278wWt4vxxXcMnse3oNfdV1lnjMvt8SodvX9YqHhC+En7n1rK8iqVMA7Fz2NgAtbfY1lQ
udcce+SAAc1oHskqoW/A2c+n3disTe3IB6hh+Gp40YXj8hoq8w7yTc7sAkcrt/PS2WvtAgcU2CWq
40nPsGEjMw1HU0OP2eC5OxRGAbMkCNra8kpzoSO0FT5bdwxYzTp0gYiWxpSa/C6Rrq+aeG50ynAO
A666uCBSKAAfmM9032F5BQglo23knBpvI4118E+D1eSSPaVthKMkAzTbyuSIfiyOw7S3Gt+wKnr/
PMeTOEGHRxy+o+qkC9gtn8rkAAdi7ixl5SdjqAcvlJqvX4OcpSutjuj6XQPQOQ34vRHyETL3oqNZ
zC5tWrhd7MmclUtpTUqNuVl90pKkEvR6dBM6PTjdjTxf/b0TeRolV7rE151FanI2G+kfUl7h2pvU
EV87XK675lnQv2x9HYdHR0bPOmYQVy7nAoD0CVnHbkmHgnc4I0WVBM3PBRtlL6kLbcVurdXV7zVU
loEe+iS/LCdZWNH8vOVbS/xE8i8tO6dNgAmUxdFwk/ZE55RzVRo6HBBJywQxP6Jwpm03jQP6kitS
DFBAhImLtoQLPXJGT5bPZEEefHObTMySP1q6opaR0Ri5pf3eJBVDahMiMovye/87V48ZfMSMZEet
SPMRyBH7vYh4ejV73C0OcJvc0L/2l0YEpGOsKGCqFdKaReDlhHl29ALAqZxHtXCmfJb/4WwcYCu4
5z9pSVaLtMRrQLoYYQbYz0j7QiU+g3yLx7CnVJZ3V5FzDdQ6EZz58aMKJnzbif+Q7GNmT9j6w4/P
cZfp4m/2kGo7rq/1ZfAPDwBqIBIbYNsi0gv6G6jh3UIiBDOWM2hEVxMo7H/o5PGZfY+rEm0dzXR/
CAcuQblarJnsS8AH/O+bGVFp9r60JsoM0nqD7xSTCU8CcyT3n1hsmYUpRjcEDRFOhXA2AquXL7B+
T8IQs/8TMpGe46DKCaRxbGuKTBy6tkT+b6C+Kz1AGOwhNO2W5E3IYeNtFahrXOIflPitXhlLgv6E
D6MPq3Yx4Gd8cw217r10RMhIgw+TnWwqENMjdCSIeYMT8Kjfo/UmI0X4B/TzjNkPr8L1UhcD9NpY
YpmkNddm16gQCo7N2Ov8BIf2uwf09oAZ9JxM9r7CXJXdf0h9D6+KznVdHC+MnJNlt+GxjHlPL8ZP
9iR0iRgI2/l4XTlED/d1/iOHz83BJnAWpYP9oU5KG2clESCqjfrubw7eZtzhIEH2GbkPaiiVuoKg
cAFAekGJaKbJmJm/yuG/Io8eoBIaZseOuUaivp7PXglwCj+yWDNPXJhdEk2Wv3X3yCk4KrmZO+Ks
KFZYS94gA82ElBArfP9/iJ3I/MQwThV4x6o+xmC/VB8YbDem1yDYdoQ8m0/YcCElQ49x3wgAAT0W
ushSMJuD4rtO5nJoDyLyF6h6iuKTaGnsw73jpI1aSRicMAHQ2geeB7UMOATd/LV1TDsxpfz8YlWB
2VXk4PqHa14t8Qn+LlKPxwwJ2MwwI3ep0UIWcbGMuzOhxWa2QkrOg6l12z37Pz3nflleYzgb3dQA
fdAIFoqKMG9TmgGbmEQUiHbCY3lwD88AtVMVGN2eO9lBEo48j0tiAyMOBad7ip+LKlXkXT6soEtx
VhpALtj8QwyZhUagEPTOjWu62iolIhTHoEkAtUPX7WWwj5x1dyjz6Sn33nbBLHguaqnhO2hImMKq
O2LageURMHokavt2U0+xNzm/2Cg3JziT6Q7lM+R7PMWk4pMaTnxKImWhwGGB+ObSeQO73FOkaTmp
lMdNYiNVZnJL7aE/5NYGwDadGElHvQcb2JYclTCdeayfoHVR6ffgA+f6pakblaRQSxey6LaE+ots
RIFzsc766oP4BcgR14YblQgbz1VbJcSh5wE+dsD0QloObzNn2R+6z+ZtpFyBy/qM2+DPLDIrFJ3c
+HKke1Sp8gZkdmanLYbnHKcYhSuAFHpyB+fUR4mqFDYqUvo9dd0PigkcQZ8ik3UbjVWeaWwZejdF
k1EkEXKWhaDEfcZ2uRCMrZj5C0MY0Wv9zUOXmRLccY+ZFfWDtq9Y5ThnXGH4IgujFrkok5jvkYce
qzY9EboolshuSO+vAbwEybZEGVr9vg+X7ePWvSw+uInhRdr6B7qUT7uZnUaRsSTbyjBatFAirudF
1AT5Zt6WMU+0FRBLkk2Dw3kU1XhuSj13ckMuZVoakO0MF+nqRwSY1MqC36mKLU61yuDfr76blCk1
URz7f7UJYyiNNIc/5de2Rl/ShY7R53m7PjmN+asoN8sRoTxMfJ+ytyWsfe79zfTiKYPideZd2cNq
vUH07RB+qiL/KyzLXwkNbQfMObEakfKtgMkr70wH5Dhp5C9vS3g93DgWWCOyTDv+8okXoTx0MQ6d
IDL4y87kIQU0mKhLrqi4a81MsE32X6gXbAGvIiUDWq9LTREnr8vatk8WAyeeqdcQobr2VDvQw3kD
TQbhzHed/S+ZFVzfsL9nKid6hK1XUP40/Nl5UzzknjKONfOfIzaOlMPsuApGmZ90Sd7w0htPMSmB
d0+KpIh/Jb6aLzf0JGVNcnPqfIDv306CBKJqv5hWU+S73OpCwySxOlKO26F7+hQEntcvOa4vKFOf
H69KUf06tcgMx3E+OFrVY4LxWz+dhJk2RXFdeMSeB12KW+L6DSm9pjcmAJs9ELoRvT6GcU94WauR
WRKc7r+DGQ2nkk/cJ4dFae2L+dCz8/Wu3gilpMraVfJ9R8CY4vMoPHBnxj8u6BJG2iz6GGKjaGM9
xmWhzgtIrJeZJ4BaEtld9LPLWFFbiy8iuqW/9rJz8isgwtRdrnFnMfV0LztjQv1h0R95EZLXj0Wq
znbeZRxTKq16GgwzZ17ffvbEyyjeDuBV3Sz0s9PU/0m8zHSmP9fF83xA8s9251GyHy62G+Cw+dzU
BbU1zufLODWG+TgzrWz9zYphWjhrWpWXQ5lEIDXpHNyKQpgQXtVmApx8UZE7bAk9wTL02NgH+X0+
fG1HKqr0/Mic/9uLg3xhrkfeLl6cH3QP/WgkO9yxAX+4QsHFCmO4xDayVWqqxyp4Cmy8TU2v1tOe
w0KS33zf04eKBm1Ya9er2ltgTpUnyZugW2XsO4w8LObEouo3OVHq349vz8IQiX5O8eZt7h94kgBi
uarRHBjRePR6tIKOKOZzCynhixqlOBgjvTN6KrMDvi9Jydf08Fto1khkmJB0T/ewMfPi2clPp0lm
ig8wPVmqcaftrDl/mhc0MRjOvi2OiMhEO/CmA9pnNL2ZZLPuFZ2iVhrucroajsa1Mg/bw2m/Q/Bv
VlAxPHYQ7cSI07nmg4YxkuYhIkv7Gd7FFAJpPi3yVMOWzBXKZd2ySNJiyMggHVLRmilkxsPZ3HLC
K1qWAg0x/U3tJDhb3OeY9WyL4CN0oVDmLqYgeFFWXAH0gq4N21THHz5yPj1Ey875CRi8NGRGNB4V
fI3f9K2HQrgsCs9rUPAiIirie9xoVn/RwaaWVRFcO22oHoRHZzEvUzIHO9RYIYPfsSvc+ZkOt1fY
mVOaNl9Mr74nwOqZqu7LhZoO48gD90By4Xt9ZkqysqJ6duwhzVqktncHoX5Cq3LPqgvjYA/k9w3w
k7S6sSyDvSmy2psZN/FNUNE3suJhRpxA+0qhVlqGN49uGFDbf7TCrk1eSkWfqaV4j9Oi+O5JGv69
JHV3aP7+NNUPVX2ZV2UBH+6vE7A4eSS1WwoXjy5bV3H8sjQpkDx8W7o70DZQX/DGImEFw8qbWpyZ
Y3xL7fTHoA6hnHCE4gqTg+jyN6Va9XXXNSDFwLLosc71RUVsV1n/zbHljHgf4OwSJb/NlCl29Yyh
j06WP2RacG7G1/9Y5u8L/xHcOv69ZinpEGCTgbx0DpZbpe+AB90poTJJuz1QVLjhduUxUu2eOzSI
WAMw+S398Bf21G7WJIcEmt6MbdHJqNlmxmXR/G3svOtZJzv+J62LV/e3yJ21NBdhr85Nbgkk2T0y
0LVbu1IZk4djwOmETdLPKKYUMTF7qDXaoAUXACB72QgoZcb6ovLZBq5hfsbqBO+fgoPE1HMzlj0K
jue4D0FgFinBLk+qg8oPs7tpAvpH35bxGpKYuuhXbzK2Np6QRFFQ4cKgijLqvFIXUchVtwdKdgno
UOxrn576zKgIHj1YZa5dJLfV8dvTDUzNvqhN3jcwB9tWoewkJDfEGVL0zZnVI/SRt0xFJw/Zs6Od
QESlrFEdsHy3HvFb9DZjH7f13VZX+pI3q6PJHPlzSufzRUcuA1ZXlq5/OUPXS+JIzchrbq1XUw+1
Pamxx+ggGb2Qh27ZsXmvnZTCIEt9sTpdViNyivG0/tA7js4ooZbyuoDf46Hz3prw/QBYfwsv81K1
Dt9yd/fLVmiyagplmHNE+j89ulsXKiJE6OBT9kgzCBwElRO0+pCxkCDl+xcI2raIh3DSvlb6lfdY
Dc2xZ77cx5Ak4L5iueiHSkxreA052uV4fUtAZaCBPnoD4RgFaqGObLhxJH5BihJBOa29On5pl0em
DobvgDDVe8clCahTkfbB2DEzD6hVo/IbHrE/04LlYriYDxBHud5TFCCMl0l9bVi7WLoxyl0TwtNA
eg4cencfNnYP3x8pYcVVTHCa+ko9HJctU7S0XDpyZHuBdi8pMjr8Ous5p4BuJtK+IbvjUrV458aa
mBU/oGig/d2NFnzboN5zoYTsEBOgWWbGIc5t2Omj/vgY8bEvNDls4h48HEzaKjtU7vAS6L8TnL9s
4GBBxjS19yrJrwqoQy1FtQ8KJu7zInoBDvl1GHG9MuqifCjdJzVw5LfGKOAo1fBDg+TCkGjeWUw+
zuBJ0VZmUNLG2L/TyCK+5oxqdxiHxf4sCu+p5znnkbD8XABvtTcQoPRcSI3uB2i1GuhKTR4o1Cvt
kfaFPIxArwUd7u2LB2BgOwbGidva7LpWIW6/yp7q8kLMq5YtfHEvxAttYMk9JHEJ+5MNoVRvoFAb
E2IgWyDq/H6FjcGFOYjOTf4BDuh4KrsQ9GY2LnRL+2D6/En1yyxNYVSmKmnYifk1AYcwC1yuyQYd
lLxBQqqbhBl6vwqQLjFYHb2QWpyaQU+eBoohqgZbY8Q66rdZXSEYRArfXM5HYuQyrurbCS/7BV8U
qxMK/Dbgc02Z204mR2MhCPlmJ1nb+J1+/nnSheVsdN6rbkWvskoZwxpqBUxfNhNyenif5Q94Mk5h
EruZWf/ZDuoll2JR8Za9eGPx9F6bwsYubqW9ZtmRVL64WIH4uk7zid6en3dQk6HIZT0vZ/mzCkXm
qy/GD7JHJkqalznfEzUREugLhDa31+Wbtoru1e+58WOwrjZlyZkwpSpjbhACQOkGU3Htams00Di1
JH8lXcjslMbegSUE8uHiMu963Ph4r0n12I7ve3BN/HD0k2uRUM9/Whl7vbswYeaB8DKZppm16c1c
k8vGzwzWpM6WesZDtsG1f0G7wqdb38YdLONx3QAjkTTvbqWC6f2rBLMNgfSKEylKMPwGzLLrbLzh
fba9U9flppdFNwrzpPNFlhMk84TcpH3HM4YgLQzTmx1PHOFsM/aAUQUs+x35kdJIMzOTwzjN38cQ
HSoICUT2pU2q5h6x6Fr13SwxS6bGXlVWdJBuiZVgju3nEY+uqwou3S8jKwl1MfNa1DihIrsEsFOR
rMFk95Xk/wi03JNCGafi6KOn4LZ3VOuxdIFjgT29JXObEkFmgvEsNLZW5GtpbnYJteaugDydgPhR
FaTECXRKFboIb8yvTnkk7yZ6EEEu6DuBiHo/TTEDpTdOdC6bIqnQcDpe+DOds6CMJCZ0EmAnyTyR
SevQBMtybTRFDHNsOfbPmBRxXN0GGD6ePE96rTam35XqFK0fGBpiU3lfIUWtTkaQTtKx1kZSMOg1
WnuwUHk78ilsNWhl9J186h+hFIQ5xJXC0eDOJubwraX2aA+UgnGRn8EwI1ffFRQfqEknv5jDImTn
2oPGtHHk5xZ2E0/lWNqdHKI82vZ/1iklcQ9q5UWl3H64xn3UrQY9xSWeoMb24Qb3jwdKAqGX8xbT
VcJbKJsQeac98VfPgiE7u3hKSDbdJO0lIjr9tiKmBcFjFhiyXgeNYhF1BNDT7iZKAzkaBFRPu+L1
FE4Gk8CMtXaFUina9PlowBOuFXVKHxu+0HrrixU+4PpxEMtaXdcqTTAAR69zIXzgx+Z4P96GXmdk
yyR7/3WWNg+s1NT2K6sn3x+uAIBXh4ovhxAde/NUInpyEegCNKVFg8JxXpn0OZObOfeSStP/eohq
0fgn/cNXSGuZB0hDwylOSVaHbxSSMJp0ereJec/pCN9dNwYX6SVjO+I2mJSdu/Alqgc0bRRDgL3M
UmemR6NVoeeaxJqFvFCKBK/O9Ov+AWlN0qCIsqgRjqPR0eaePqDhLHKvU9g9uXINEmr+YaDavIUs
kR50P3tW+YXz2slPhr0bNIRipwBNA4v8yL9PTFH15mcw2F6NQXCF84vlRMoFd1VSx9LVu2WUe8Jv
L8fWBADuyB0yuVzX0xt7eE0DJvdRdftaj9ui1nU220vSVr++sR871F5NHWaCsjioH55mb6ByNuyb
J3r7q+7ZFRiTHCTC4EWmYDaZZUpIRwsPHkG8sfvtk+Yb8NCRAxAjO/j5CBW8JByjRq78/OaU30gZ
Ej2DO6tXpsEQyvoTLAxkcGeUKZ2a+qZd5A7rh+licygEuwLj4j6avBtKhcKfvVSBUDyYsnAl7ma4
vnO7nwLx3WDXlP18Op6seKyfOZ3ybsNtsneJuOKRJPQ3RQLlQAvy4EVjRB4eQrSI6bywINfvKjGp
SiE9MJQw80M6rkL25Nyg8L8vK30gF+hEyv0Q8x9GkyEwtzkwc860yUJjc/wWY2C5iFcalIGm8myO
IXSCCFIjPEwK0uXnB1wOHFp81M0f5QMERQcVQhMwGfOFl6OkHdzxd967N6SoUQie+h8zxoiGPPum
8I+k59qOjQzg3qMFp0QnynftM6YsT9aVBIvzs/kbtGDny0LcdOQTlUftJD7okn40UV+kQZ0e9pm8
Rdv4EghBw2RkVFXu6wqa7+a5dug/Z47XU8mDJzNk2BRZnv5d5dgchoPjVL8xgHHxOcajDtjMkwcT
qglb9yfzYqkDOoHx/xbYqmTwoBtGwMnSZgBt/X2vWju+lvoY5zrRj3Q4mnX1ZXiEBmkq94KolKFC
Kgj/2ssIqYI6nvUKtGURq5MMkuL5NFvH0RQkf+q+CLXCEoN8oPZ1Sk5AvS/cC/NMu0Z061bZdnLV
Iw/d5AAerIaJGS6g8QCfmWr+F18JnmBWzyseOX/MKfINzBJ1rcPJVwKvwfvE4RE7ZVOpoHGFsrS2
fHsjlDfsJ7HrVYXPzU0I739b20/2PaWxSpfwuWIUWkYeUEoSkcRLUynbelc9JFQQIYuBXVxTz98k
F+dGdGm6EBZJVaSwFExraD2kXEHx86kPsLyeAkexHaUYBW2NA51xQdyAbb9LY1jejXL6HUUSoGJp
GubliL6v3WIlwLMT5gN+4FSYCkqYRIB0bDU1KKbZtJPoWvbmkYKJ++pHS9YJzsEFgaVUsV6rw1kJ
bTyG6m2GOG1UqoIf1R1iCYw3JQw6tV/3x4oJTSIcvQmzAOEuETg6WQynf3yULsdKIaa+Qkn9CdHj
ioaduYu2xJbDb5kkvcRac5ZZymytC1tE6aTYEV8jbTUBqnwDIN6rW+u/feKGwGSad4GVWlQI6ZwO
yU5/cbzKdad9RtikVsv6lJDgE+8Uqxdr2vOckaS0lgBjG+WbecwJwVX+SWDjW0koZUURwkOzY+2h
aX8S5r0q3vLjulNeG7ixs76krAsu123wsvB645d3LzGCyd0GpzLqSv6YvMMZrdA25V1L6Ds5e3aN
jNKYgx6tCnjouTiwKt2gAtyse76SL+ySqKL3pRZj7rv3RcOfe6WLFq0eG2KgsWAWTFdTVsPcK2X3
pA98efkGUf5SgrJYlJMLfQCGmUe4H61zvRr0cOe7epsI2k3/hRxjJqufxpzH2cVnfcMaAk9224zn
r/lcLEo4DR8gFSnZCFVX+Jy28wDaT7POU1fPbgxLECynNm4NQPHGv5lK71tyJvekxxW5T3PLmhY3
4nXImdAhAxKH0YY3Y62c20cqjpxDXhybfDP1uNdXkhwSPSw5xvxnLb/jqGovtzlkmNAQY6Z77GcV
ckRjb5sAYyUPbtY0oKaikqfG7RtVnk7rqDB7kyZ4tnGqE1RP0U5nc/G4cdKK/EpgnDFRbba2sJDm
b8i7gbow9QvrnhGltY4udtmHz/85X4K4U+fpKMcAhYyN2X3Qy+dWcdNpA9O0vr8+PDJ230cWiAbN
TbR2TgfCQkThDlA5ylsGePmWd/q8MnvdenS9B0V7PWXuG63vw0HPbF9VJxyx58Siz5JRBFD27TZg
3kTnMItUf62RZ+TR2/zcei2lxEJg0u4gY3OaZm0GFAvGCSAJjix5gqQYwB44C85UsWzaHzjZs8Mb
R/sNyPsbdNINfJ2UTPm9jEEzW8kQBth8kGqnsbdZ2oE+OPazZWVn/otzrQp/jweI0rBiU2W8QCr4
R57WUKNQWQuQUwMAIzKJcAz3nV6uM9AVSvoRZ6Pwjfm9Jrzf7jSWSLONoJqRzVKwGY809Jl/s6Ab
klcXKJ7/BWawurGkZ4gq7/tLbWTfwgIMpBZa0R7h5UCP8cXBI+etgbgZgoFexG8OUC7TNuBlXwEa
UQLNLp61eNUXgzJKvMjNtZ31BPIsXgWmjAWf89enK2YEG3NGiH2h3EhdP/V0iHhI33fGUhmBsy+B
rVzfTzqqpXQnoxPwM9TyALdxm8kcrVVCvO3mXHrkRoAjCN42VUnLCz1rBmO7A/cFX3CZVmfWt0Ti
aFS9jl+LAyBdbO/1piAVNcEtUjol+2Ly0+O+if8oE1BJypp7UvDn7+cU93oD04HpYYjN8st7LrFJ
A2sxyccK+SdIymCiplOC9LIrRa80VgbG3wjiqXxgfDFWftygYEvO9NiA2pqYqJ817BO/Do8IGI78
sbimV/v+hB6OEtXlMbWV3OFd+Z/kw47LdDy57ehJ2gTl+RDLKfXbs6pTYslMZMTrSM56clKjtg2a
HwxqW0A5sNmNOuRLxTdJ45TZZOiKrVjgUQ4ZJh/IRRtpDBH30+yl2BihiEJASMQElkf2WBFVyeNB
1qZfzUMMgLHqXPjDG9gOdNpBHp/lQOxyJReODWd7xDjx1tKyjxcA6W1ww3rtolI30YwUanBYTZQl
/9AlRjEx6Truy6DliGqPoTCCHpfJMF6KG/uthFEAfaRULlfmepMqEDbl8SvfJ5gbz/20d9m31gMS
3hknFVjaXNlUjxBbxDMfgzZOLib7zcq2Lgk4evVCyo8wAUf/eCt+cHGPdTCA6vwqWkkJ136iNZnz
s1v0Ul+6WV27SAS07+0CTEjELLRjPhKHz3oD6GvII1yYM2Iu9K3MHRw7PexR/IvZrLAXLzdIuqz6
H++qpWYDOAsavPsWtnI8QR3e0myc3rwWxfsmmtq7YGiQyLfrghI+xGMfZY/AKt0fb+Ok6/5gqCmt
mOUT15aY4Y8mPBOSVMHTzv1wBrVy84Db+kBNZbrZSyKmzxJKF8hzztb7vXbxyI+OP3apFom6dlgx
yd8ML/W2YOuAUV+VJL1xYKJsx7MU52fa564tjmXkp3dRxV9zhphf08+ENk3pd8jJZNlngnGhoDbp
Rd2Gvk4kJoCdDizpKixPqDZidxtj3G1FeOHmvzMmzOWiEaHRbIrb4MBAReGshqDGsiTJXgAyAA8+
PgdNrTFdz1vLkxmcgYVdoyYsewkQUQWiTiwsn+K+a/gjedYLVRx0bfTfvggLibfH6VtEntEWbIfd
83HgoFGPYMeF/aBMvBnNnPTvynQNmFKdcKdlFM+L/LeR25g4Cc5OvHYqFbCc4fSp4xUKDBamldjR
ONZDu993dQWkR7F4Uy7Ri++8Tdbs0jKbfTmg+utSSlTlETbG52F2QdznXpORUQ2Wkht66yJgXze9
e5La+UdVgDZSIYnzngA7+4mN23F/KkoHi3hNKWnivBssagZh05cnFpuZ60qLeITrTaV9S3hTtaF+
Ge4ZIF5If9zXBY7CuuSSMpcdc7a6GCF581sjQ2airUIffRFB/6DeaAMpN8m4FVT7xhxPHoXTndg0
9MRR9bm5ayYdMbD/RchMHEHuyBEdFy4yXZ0kq2QgGAzpEFaFVefVsbCHHFwEEYs3FlSoN7QBkWMO
rOQis32vS8cDGEi3piTdmH8eaC6R3C1PbcCaQPMl4SvNtNxjZWkWoVtz+sGGGBG5Px8jlp7pT6VA
IvoJXaCj6z9hHDyiyXTocgIgqd7yGSGIyQm7/uB+J0j3CCXUCCTOzIuo1c3BgfomySHB/VUU7EPV
I1T11AW7uk0iLDt+RQ4TzcupmdzeNUFFJSU0DsmZ1+piCoFjgkbdxWyy13NnUFmJ/WRhEV5TnfqM
YYxQoctrvH2NpeYvID30RjpX2ybzFE/t2hlw6zdrhu4eUd9TlgjSLKldheaHdJ3PzlkpS0dwKM7N
VTouYzrIqGwhXj7+Q8qL7SChCIgBRFsPntfaL9Ik7YfOvABtBnk9aI+eENhX90k7xFgUTSmPkXPn
1IBYQF5r2KzoZDRUi38JXUVLOsAxLeYj+uOXvAcQ0NjDQ1Pbp8fvEfGnqLF9Rm4ium+1ogBjqIyx
oDxQFVHQLlKEDhhvIXueXmSXy4ATSe0wMFPj0ks1+/7v4ZSPsQr3rU10WOtS73I14ZDlVQB98cNU
3KMhRjnPis+rVzZ6ZV7bgljL7/t1iRgZLbv9Ajaa4hNc8+Pvajhk2pPAslf12i3xDmunlzCSPlrR
Uvu0Jo6bB9gdVFlpmCYX8yCYJJkobpbv6fO4HGIPYbqVdbof/asJV3YkvWJHZEIvUg5JS/4qx8MK
/slqezBwgYX2dHwv+Qd1jBtP8XdJr8wad8Evv4tKBAhpjEwwQSss3s7HhlwBYjgA4f438dOPe7e0
mDEDseRfZAF38jQ4F+L7VOhS311LpRwZLgXgY5UAAWOCZ1W326pOMPBM7N7OmxBo0gqoAxpHWMkU
7Eg4bP6iLj/QxWqK1v0yKeIABHpy2ygVm/Naa+Xd89GwqTCkfJ/+VmdT+auiUInUw1Ehc1dsOEO3
BHdNjlm1JQTT5HC+cpr99tNHI6+wMl7rGbADhsABTGh1lihWbQgkoCK35ZvtlC3bnslcrvkH0p5U
uQL3j19p8M7Qkjy9xgOM98/iT4e3+lgdHoqgxNv6VWJXcoXHWoHvK96Q+OeFqGaN5CYpLUDAAuC4
wCfEtJyjBjvb46xzmMQRuQbJM7q7gutuTRdU9/uJkRAspqe5dy6+aH4W0jNVudoHZKhCCeaVyzSL
pssKranWPvMttePphqWzy0LzHe5gib4tWjEqR72ISi8JZOjPzjFVvZxE1TyqAb8PIORfCvd8mpzH
u3y1XuKCBgGnrGsJevUg3ZDuVnEBpgeSvFFRBxge6X/yvlPs5gzN4e3NK7/oOsJrYmLu9T910LLI
G6drgzHlzKBmz63aSx0Olvq6Toer5iLitW41jWiQ5r0cJx5s8+i2YVi0oqy13jzvqWAzK8Y31l+k
lP/8biUzTlhcVwKam9HZhwBSgVjG3Ylr6k3gxhvtpDgFu9ZGbETS7vzDkjhBKUs1zTWubtDt8Q2g
E3heWEoD10SZF1tZ8IHFctrNFAuFrh6ndqd97bxmTiojkeEk/LZ37UiQJjPszXpejTOGOfzM4rtJ
STRbSgyobt5B6/iav7JXpu5MZDjpTqYVdIpm2dWykrQ6hTBY4fyPKG0UMvkATCJ0O+y1EEVIguHT
8BRcFHOtCQvtHu3/UyCcKl31DAiVJvWMg/znTvQWAV3iiGueZyVMCyp51MVp6+EaxBm2o7kg9ben
qUbnfEOpAfkalUHrE+LNI4YgynnQBaJntbMBk/eE2BVUZpZPCPrBPjFdxbwBvjs6uAEoIDeVXV6g
JV/lDcU0dHV45Qs4QNMAGGfBCjbVDppwVDD7I3DeR74W4IJCg7sQIzV/HRcHUVk5mPWiHj12q3DL
hUeIBS0GI2WIe7G49FSTXlX5PRJn92i+1yJOxU/R5BEoCYgwyeEL+cgqM4sAXu/mNnFLtvZbo5sU
6hU1J5fXQXWv1QrjaMOCdlUdr5uHHuxx5iV35X9hczwt3sGFbSJzKiDQmsvh/NruSp/2EaXpkuRR
6pYTD0qxnG2Sx4MsSZaeleFcPZRKG8ABM0NAinG5KZG8XLfaUdISrGZbrDRTN4+9LAnBYDC3tLc9
xF5s1IZv1uLBUFIqd7NEURjTAs5AghTAq9xsNHsq6DcnXMwwT0XeELao1G32pSPvXiq8GaWD9Mfm
D6gPIzwhGlYq8dtopSh8J7nAAk5w+f16/gJZp3qurqLOfIe7/tMTCpB/uIthkIfw3A9cKix9vlVR
P9EdHXFDxQoCkUTx//asntTwb/LY458vOJ9G0V1n23ba78E8/SbCkPMTeqo0Nv0GXhzc4xvYjE44
HeiwYHy/OPntPXAZzRHJ1YTqWtnvmCt2bBz4ib9RFHG4GobM11/eAuLrPfRJQNrLJHBDiHhUvugz
QBstemP9xSaM1xJdiLLvSAReSEdkMsO1ejjiMYCKN3vJKdhxVIyrklZ8HF1xSgCx1rOkztyI3ja8
5rlSw7LhjkXOvuNOk6a4TmUtuRHjvQzRRdHm15XRDw/MY5U0N+Jmu59vanIIr38FEw0cuhCRxqzN
U4o+iZE1At1cyilZj+BLBT1FGBLW85RAs2hmoH8k03L+8g4A7VFvTtRubOoXb+tPnI+tCnBYlXcz
04jRYufRMNNmqQSb3kABIPfRvtV8NkI76FJ+P2Nmugku6eUnXZEP5DqnsM4KBEXtLgO2kCgBk6q3
Ks6ZQ0i4zWBsHLIMV5q2aJwFMN2+Yflqta6dzy03g+w3cBaIfHM5JeF3ZXTlUl+c64rjOh9f/F6f
rNXi87vd7IQV1rkNIPe4+dTBeOPazDpZN2s2uiSCn+N/9W9SkR4e8kcfFNjz+j/wi8ON/j7arscj
O3/HJSaafRTsNVc56oW0DJm0JMkF8HPYqfYYgLgqYEW5BSw0ifofwxO0wg0UM5BgjSFyBQMHPtYG
orfQH4ck2PCSAnyDeRwLpR5H0NLaiFYecmpSsNIcl1yaVrxaVwH36Kowew/T7LZkhvRATY15hiM6
yFK/pVdwLUzSygrygYBFjq0fuRha4JpGUefwTw3uHuIa3hMcZc39S/GpULE2PD7hcoCFxCFwWtiz
zQym0gNJiaAGAX31GZs2KfB73hCHCLvXNToKVklzSbOCqmFalDcvUno3Zx3qQcSRBuvJayj8nyHc
AK9d3UViL2xC0ABtoxSlOX5FHXMhuv46Hr/E1S17GJofruQLUS3QPlE9yGOaszfSHF3THJDxGSco
lCadnTWbR40ucW/e493EPBIaH3RBdJ67v9SiF03exQ6Jl+OGo3QY0ZVePXKUFJpJef3sCPb7Oqi9
0tObRmfvCext3s/ROBK2gMszfHjs/1CQXuqYmVKB1WvlYtkg/UAI/lH/BtmjQeSmj5yTco8gz7Fu
IHkPviktfhOm/zmkwGA1D5hlyVRNIPNg4kQfYniiTsjqpdQoxopf4TP7zd+drto8D/m2x1dVz+0Z
zy6/rO0BrMgxfxLUwXAMoXfpWDN9ncrYuc2l6qEWM100ZtiuS0YehGcNK6TKYkl5oSrLms2Oyy/E
6bqXjIb2lGMH4mEZiMGeb/TNe1N6bB7MF8hVaGe51PpsG5ikBV/xKvBwahzAC9/1E3AnT4unLoph
0340TRt07hpoJ1sbiN1lFlC9OcRIYxps1thPmlGhDm9eO0QBnvQq/+XSg2y0NNAQVntQmHM928p+
UJx5qEK5s5L2QOEwZEOI03PZ2UBalvP6IPbtjZtO6ZjfXgW3Pa6XYhLhCKnOSu7qQlDMUh81f6Cq
Hdy7LYtB0bFQFIBCeUIq89mKySMIukdYpoxJ8lTQPH+gBLFbNfX/4NOpkSoY1g+yP01r6qrqlBtN
yJuBwrRgalpGjxdo3cXrgWJYSxnrDWGF7Zu9Sgw5NJwDf0e5MUAS09BYfOXZgdsNdAibWM2QNPpV
1rTKWpsk2IsjOhpi5Xi9Qy/VlrUUTq3QczqTCymvwdORSFhQxxhD5TUQg7RIYOwcbfhOE2WQRvMb
MISlplHihU+kMDaj3KEofN9tzivueqiLM70z2tE+OL31AE2PYDiFA7Fz2pTljbKVWfaSajRxe7d5
RPl5jhSiNdKGHRZctIT1/Hf8MPLufZ5sjTkXStHG0m10RdFsU6LawYfJKZEPCuyi9KxCtyUB6BMb
Lx5k+GDh4lzvlRqLQMY971/obDDlG7NiYV6RfjUHMdo/1QHSpqWVfE8NIExAsNc9vVXaWKREGbDK
yzdO7cSpWXyrt80zNMJqVv32IGjVWgO7tVYA5FIa4K5Z7BSAflFOV8bWgG6EAKd4OzfGJSacdLxY
pC07rhyTPcog8CX++AKMGJRJJ8qrSA26EUcOGE7kV4bPU/1jT95T2zx5LGHmBUIwH4zM8ioFSkpZ
vUlCOb8ULWWDYP/59EOTY8uxQVWcp5l+7Tw6z09+6QrVRc6SnmmYtWap8ExN/y4f6k9+u8eKo7IF
5RviwML8YA743nlIzkJ8LmijaOCa1+NFcZOt8jepNzVkH3UdQpMVyzhHHG+vN/h10RC1mlrTTIZT
DPjeyMIsM6uWJcnsdqc9EagCumLKEyrSc0nUs3cA+OtYOlwJ7749gD5gfMEoW44FfcS2yb5VPbAt
TJQd3Vvr1SRufOoRF2ncyOVX1P1B5qCWiVsQXm6mx39X6UX4qYK6ry95Q+VCAiJ5gjIYx2szlqsj
8DVLUCYbxcAvoJJpw/oVlsHy38y+FCRkt+2J0AI1xMcL0+9yvq44dFI/yz/tpsvDynd7qyy6WYRY
2NeLggtDgqP0YjUHdbZg/QtF5GCAdVExdQf0/1ComBugB6vi0XjsdjFtBO2vqhPuyY/R3ZjtNw93
9yG0HEFqeGrt3hVLH2s1RnobR5MlH4TGXOXDMnGgatTFQ/pp6EHyYcpuWKEV7D3WUm5DziiP8U5y
g1beSCikKiC+fUdySIODoxQylm2Ie1DPqbwIzoyt+6UOzKv4z1My5fc4O8Xz1qXcIY9SrndcIp+M
FdL7r3a+1EZ4XFBx8hnePAai8NHYgmISFY5iPJ9tTd1pR/JAse0fLn3ccN2Z0Vvo/xEKFgD4n4j3
8dxh7nJtiRZmINqb0rxA0u613YRDDB8s7axN+aAxJLlCXv8SRONTVLsFvtWU/QTIQLd8cxpBQzfg
Apg5fBe8DhqlQ9DWjm22ONb4Cu4Be86FR7vnbGh+AKn6pDy6Jv3fq/AKvPjQ8YzIP6Jnz/B5IM/U
+YGdlJljQJ841psXSvP2dJfTovx659X1p7EutkZEsOqvZGVwELvT2g7HctKo+kvC90Rt9/lxF1Y4
cKjMMbHifojG+1j6NfpVTOJbCQcuNCrsaXhlPVaQc42tKuI9Um+W+TuAzmQpTFhKMBTucQWQWjJP
/95kvDpY1bYxxqQYCJ3k699EEQphbFfQK9QiUu5KtANYgujbWMz1DXaqmSVY9HjkS12KqDT3iz1E
sC5Y+zCzASApG7+fufmNUBsTMSmWMupjZSi6sro4CTU0Gy4SF0Xg3xNdTAboC0rStgYtPAlyCWA7
m4kQVoHtTYHks+89i5pJobHOft6/icsTw5YQZOMz5u8/FxOVYMB1KdASF83E9DIa9DFBRcHzOOwm
0uHzHU40NOL9fD5Z1oACIPusQFgFZbc9dMzej5d6Edh0g4IAdObJY9aIji/OYOHCE8t/o+9fYX2S
r+fTHh0jSh4wR1T3P63EBD5x1zxhw7iWwJYA6vlmJ2DqWbUFTJ3ii+ITBi/jC1kwD/h6bRyve5sB
ceNLM2ENstoyuaYhMzvgvY0/NiH3cpQ/JqS/vG93t+r1ng9NiS8DXUVoY4GovCdlsxmZ82MUIbni
7qgFyJ034kpkFvQtHKvD1zwMFC9l1s4iOBbM+4q3Ynaf0V3m/rPPK9v1kVa+yT2lZX6jBpchi5/9
wv3+/Z0ud4khUp2Akxh5ZdcHl6k4XNyBnNK6wxuDppR+1iAClWB4Pji1AeEVNLynpmutYmGKLLYX
Q5gmU3MFPL7XB1ZZ5py6v3WA17MOD2ZsFpkItC58xGGQPQgSOoZRh363JsmGR3I0+U/7iFtBf4RL
7hMlCqKxATqOIfHvaYiy17XeV+sXmm3c/vVCZ0qFK5WR/SsUIb5lFHykeN3PsUQs3ETlXDYDDYtl
qpEPuE8MEn9ZghtTGKfazr5Q1BeGm1yt1PjUidMBzNDg5wnJ5n4uxvSWaAenOdTITkY71dTgFtnj
L9woh3BlFS0r7kz9Y3cpTZISI6VN82pd57hH4XqQlwM1YkirW/0uC/ycsJfOltYVyCNc7RlO1U4O
bLTZ3kikEdhzdWN5YeeVlOgrTw3lV2ny1FVnt07rdmq6uQDv/A+tdxw30MpSvgvxbXAGvTTEPfwL
0OqOa1sqhEtkXXEnWuBDun039nh84hM43QrauYq8CWC/QMxFf7NxjirfpenI6p6MsmqVjyI29dPI
NVDGHYa8kw/82jJv+fqCamJQSsUOUKmIf7p2YMU/+gvLss+0R7qmi/YbMoHY4HEfWhKYHkQ6eDGN
mbDCqkbNF1eSHSDezszFEQ3XnLP/8CAmwIo4lmiDBIt2Q9UHwHJALckR1B3nfB6EQ3VP2UsST9iS
YHAIJSKD4qHDIi3o2d73KKmCVWoIbRFRY16NjKnfR5TVCUPjpVxgDDzZ0fjv2l8RJ843iwj+sczA
6JG5uI5AxgqaIUWcqQazbVdBq2q/O2lMy7apTTsIbslBcDdpI0VbKA3a2aljoE+XvJ4MtWeYHmn/
DyIKRfo5SLCtcmrcR3grNRz5hztT+mAD3naxmIDdNKgna0czpY05ehWFCN4+NXwBHVYELJ3qYUPU
RQOPKegfQmT+2CjUoqZLjjWFnBgGSX4UMF+vfyjAKorXiFOiVYQT8QGr8O50+0Ryuby1zgpMWXiW
ZyQmoVqG9NyZfVVqggUPNtsGP1EDELqkVr7m+Rg7C/BGISZ0bk0v/suzC+UPxtTfNRHIFLAtu6ls
A09dA5rBDPc3rocnJ2GLQitC4xBDNKLBkjkl4vQKyX7cZ64aMFl6p+eiV9H9PAptR/4BkvYx7tam
OHdCZx2poblbvffhTPRM2uZWfyb4y4nstjfms55lWI7uDrGaCbz+Uc7SRV4s3AMn1OlvqLwCT8pc
0d+22JL0s6PgllO1DgrPV/h8hqnkkTJiEoZuoqiKysjqmfsrlBywA4NAk8nURqYq5Rw264WVVrSL
h2U0FDngzDyai5i4b/wfNo8b5cy1m/F8N9vt/1ZWhyDZkwDKfbUuSp4SJqaZYlmGfwVU7Cq6/IrQ
P7bd0Ap/3flsn/WQ5dRF72B1JdcIB02zYQwX47Jit0mZzQDepqv0witUExH1vx4r5r4ECbcDe6y8
Tqmyyv9qsVEj2HWWsiHioI8FRyddBV5TT1sE6pz/9p5/7IS2UC7P5uqtEFBJmbYlrAx2iygpxMue
TSyAI9WYbbsTk9dIJlq7rlnjmUpUjKkyXtvaKk3HsxUeqEf4wRenZnmjt3x0ZjboGwwQ/N+RVILK
un2U7x1xQeaawxSXlAhx/HqOoDHBKllUPuN9plVKeOka00c8JJSqO2qcPHkhN342OlxCkS5vcTc2
pcafTnoBiyPU/u8pj+NsZEc0K03JNawK4g7miTfUu9Blha5yA4DTXbqjWBpMT5murgbdMhR8VMFb
aoKyYBbBt9TyqbhFL0v/J/aFIAotB7jd3D87DWkjq24ItrwenBUGCRjl4U9kw4mT0xD+LZEBuxzM
4vaxiT6rBE6oU1lwtDhDaxrYJBlkDW98+JxyYP0ZmsKDBLmca/yJJxMtM0dr3Qd/AErtQD83LCyV
3CzE4j2qiFBlHG/tzdmKbuN1SHQ3SgM4Ey7LOEQ8WuZqybitgAkBLMrJ+QSu6UFbMW0f6Csexm9V
SWNHm6HT0J1+mDKwTvuYELYpFlp0kLmh9VS0sNJLBtqubQ3jmLQQFjaPSefBjj74TURxk7q7fgQ9
CEigJC/eQMKV4/7ixHtrqYMWaLXnqj285gb++xDG+rteXunr1WeffCEaOWTlyePtANiXetbD7GIE
f2OrOM3Celf2uC5DHoZxGMyRHx39H/3sRfIzkKiTkOHQl45Nf6V3YKs/+R58O3QNq7J0Q9W3woGw
oRMNrprYBtz0w4D7YQDJPnY/Cit9ae56KoYqd72YpJ2f1yuosptDcgBi0xx0j/ELy4VyGon/lyZi
DZTHlGxa2QjDShJhsmqpz05N0xu2OwRwQpEqAARPSV6VN8w2vPfjUZAFz/gGArIvneOLxnqgR1a4
VANWwg1ki4RqxHAvvPcAOdnXP2HZ+c14v20+fcUTnO7Hl2GYDIaWB0j/OayZABezdmUEbOY0R51g
ZHY1XyffLa3LVIYLyU1CmBY1tUzogkxNLbnH0sYZljm/7LMCBcbrFmEAmEgWpbaqDV3gzIhkQYhr
bImmycTv72T28eMZMUsBnai1X2T0Cyv85y5iwWCqHklVpBTqbANftIBq8c+y7DZYAeiupKHrgBB4
PWMaICCdSLl2GstWPl7v8cC7hYTG2ME4133p7RnmguZbWrc8RMkOPNVajV+I0zYM5TXyckw2iyNU
15/VDkDc0DxaBWPDZzSEZ4j1RgSovEnMynpmEpEVjZZyPYJJsVR+n1OglppUMKMai97bL6o8j/+L
ecAGwYqvWtj2iywkTpH9Q+cI6Bqi2f7muyrgNBtsqJfhqVm83o8upnydmvNIEksQd1ow1MXc51Vu
mvvroZMmv5fNgHhrzWeHUrlZEpl345USDOvEfmppudJN/5sXHxnUjNZ4OEqGFKh5qXSDM/dKgmUh
oqbGPwdOY+cXXoDoCzqqM/KnVU/2lOtkmIjExAUHeOrLLFpP12XNePSnphqRvGY6QQ7fTfm3TeDG
FGj2UVRctyG52LBA9gISyCrUc1r15j7DoXFnd5W2sZzXAbx236IL9Dp+V3pZHy8DHOfGHlCVJmC4
W+0BZy2UAxTh/AC5IPfzrhlLcr77pmAfzSmrecma3+Bq/A1icKHggpiX8RispCY/Mo9s5rtdqyZd
pzBPf1r2dO4hYwLNxMdgP4mBE4Fe8SUWHqm9a9hXVskWy3G1JNSJgfUNeKLr/BDXiKovbDyAIyMj
9C302aCghdV1Wbzno9UgtGMDggv7OuiVcaWgism8YKu16/eaHWNsPvqkKhQDuaf/NfQKvOeCQ3wB
zuKOfrI8U0eErJaWrbizPestEiZo9XOowYXAA7Quucr3DXTRCRB0JL33uk8tFGUlOOIzh5oVAHKy
y/R23sKF8xMEmJxcnmDLy0mXeU0idctAd8e+8M3xLsVQzg9bLK8L+3kPS8kwmynN16ciwO268Qpu
ZkdCikcN33+xyfa4qMAd0mqdiHDRaEUk13X2gFP6FV/zCwPCD9lSxKT4H4utRWCy3HX7FhkdSt2O
Fr29K7BsWNbohdOEkkxb/1ObP5RUaguSiUo4iNn4IA2JFuPdLLbWRVGvcjIz4qviVJUSUOUxeCNK
8QirLT0/fdWnT/lXCMkjlGf1kHuOLFI88XN/s2iH77Z+n2piQDasG1PcehO0qv2b+k87RJbwWRQp
UJEriOGLhtaa1f7WHGw39MyraJ9Eh/qw5gjFD4+Z+8QgMmWDYEtVLVdj2r8sxgpxGkyb1lOBvExY
6ZmOLYaR4l/Ei/tSqkBIjkvWwHJkZF3b2HvYZm/koqGbBIcYmsjSUxZA5JdT+stAcfeuCHsZ4iyU
mnO4d7ornO4MbON5nEvOGoLJ9PkA8mdFX2a4L0JPdzUWy0qj1PPqmRv1xcV10/2CGc8dYGB2PQ8a
XR6x0RtjMNLzr3hXyvdQXid76cxGJERGfVFmlWbgav9fyQ1aCUSE+hmX2NpIAthsDO1/1GiR9IcQ
TbmFa08SG4Q1n5dyF9Ty0xcDRZx6JyANjzYaBXIY31maPchkE8JQBcMILQmLn6nZnhd/egKVHs9C
Sfqfkg6ZNb7GLZF+USa90sjyR5kc4HGY/QO/OeXOREt5IhOfhX/dsiV8eTJn3dzQafXVjmnT+bsg
rmc0as+yaiaclEFq+ervN1V7l8AkH0WF8ZVGqJuZsxN2c+XIoCAK/Lw7xlq13eDfFT/2Yvk6X4KP
28hUumO1NW2j+740V/nnRMXcGDv9Yg+2mQSen2cQainswEeoZzz7AkWKc9g0d8wxWpGN95EqBkNv
z/Y13e4K8CrDr4SNmbDUnJ/L9iCnqVquk4Eia2uQ5EZv1jFzgNg7qLYBRXprmNiw7Uovnw82rkWH
1AjP/Yyjt9xu5j1nEIcyvqX4fdL46VLyMGcodWgq/kZFrZVlm1/C/a/+hKk+h8dpzT1VEzwKVMzT
uv9AxeFtn/klGxBEe/T+26A2Ju2CTVxUeORA29xyyWmeVSqhbch7BIdZCHxF59g7WVnnHXxMelDB
bJuFnLxYnHjV+UZPUIS2Cpim0N6ySCVnA7iXStJmoXpQOLX7QiTTVVmday59BQAFDImyr8s6sbTp
eTvwH5qk1SHrsIwhtV2H8iOobOPcBCZ0NnUKBlaQKXwT1tw748s1cPtat6R7+B4AC9Q4ieU9fDhQ
rudPSfpUcQI9zXoq7POYNmY6iElyYi+8MML+forVwas1wl1Vcgl0dQ3L7eR3RgokELepjOuCRpbJ
GWm4VIMgM63xR4tITDI9Ioqk6kUZye9maFugr1sOiSgjl4J6za1Pvlip0X4MJ5Q3pMFaPxPCgLNy
S+kDunVf8ZcBHM3iNn/8eox3R4x7Xv4KyHbjB/7TOYd/pP/Y2gevMBnBCCDvwVJ1VCGxJEcM/4G6
XDUHxDFveXdgobVgmhSn/M7Wk0+py47KrPwseaL4bBl6DMTYGyX50zWPZiHUN+pdLBCDyPYTK0jv
Rc3gH8VQ7xLh7WnZJ5nvM+9J3TO4Hrt804GtGMuE2zhNqTDJa3Ng5v8YmpVzMZnUv1cjpFobOJSx
FmCqB5nBtFz6wrMTOWAckHKcQvhOeTG80+ibrK5d8x+PpOf5S47LDMsactrZpHZqaGYWd12AopNZ
NoYkrFaiKfZaPc1u2wMQPhpwptDgDoV/kJRaFu6B01yWvbLTvbhpta71B0hdwWweAXjJOVir1rpF
jSLcO/JT7UxBeD4vLwvkOxqrDsZcWtsqw5CA2EF5vDRwiYzpwawaUZVA0+D4tzZCNKnKGer1yMNv
qq0hK3hGqWCP+zA/7zWx7w98uiSr9Ze30hMnZws8jojjQDe8LGkhwsAUu4GiGExrcdiBeGK+uRpv
QT1jJWkWzG4H5y474PPa8zMLbrbbpHud7EEqIPMwfhDwHdnFt4UiD4PuIm5klxsZVpfCEp1RgGLz
IGqxl2xlZSXp34t3uD58LV9WVX+YZo825H4WVxoP0BKDL+gVpCgIw2gSV0OjXOyRcsesen5+erV7
cT/V5dlwaCaXxFb90m3VxLlP8Oyx8Ivfu98dVfED2pFuYY6ghL2KS/lJqyZ91z7yAavcDWxvu6KB
D1FLAffeZk2eWGotCgPp/0ID5yrQDgzwVRxyS+DZ098pPh0vgvwUcK79ZUQk130GNf1yIcV9iZet
uEj3PhcwBreLfd+WSougfHtgE07ygdsGxAwaUpb4IMGDRaaQcX4MX351lHdsG/JTU231o93sfQFg
MFyjJvXwJt3OGJC4U2lsZgh8nwSbMXooENOCh/X71b+EabT/OluqyhsyJB8OVcrGzf+6lmdOZCgF
xvNmcCYt+M+IV2F7JSsDA2tLu10mpPu+F4IFwXopVUUDyuuuM5DVuOG+qEAcgfP7p3adphUc2YCF
SbNpNrKN6/4EL5vF4vXCFe/z/zAg4PUWekGnc15IgwJBL8rN0kCtUGoe9CyXpUBiZoA5yeu4hbgt
Agrs9VmrBjYiFhgTZowY58wim21kSGsDa4fmVCcyAbJu6tynE8p5splasun4uf7sC0wjDcapamb+
j7QKR6QUMvIazmATFrF5EBNTTseYuOoeaAI36NA+LOO5wLLsxOiQOZr0zBzz+nWOQ4POH+TBXKaL
D2/sfxnwKgTBEEHTqKWwowsw2/Wltg2H6PH2rW7ATXCO21vdYZ15BOLq2txDDSL4JsKV0bUvhguy
Wo9vTVw0cKSzMZid1zjY/v6qHIey30zhy/vSPQzg9W50ng+QcS9q6xf3rDFlFn+2F79RLYOI75Qb
4DOLlc//2hBiZ552Rau3O/sHmRF58sNVYq7HQRgdd45Vx+seTYOe0WS9i/CmhLYtEw3vJjbGumAy
uZ3VFoDtA3l3xQJPhasaZvPR0vz1hWbuHCpSR9lYxELBpVu5sLQAJjKzNljl9agLdcsWA7q81TtF
S64rPyIUT2IRR2HrUfmT/2v6OtPcg2LyIpsUyW1ZpXuPsiTsuBk9FhqjgLepVc0KG9LOpjaQd++C
W8qjkvAWzXTiGa1hpbKzrvOKdWe45HxhQE0Ie23YMdJoXmzVJhi0FTKhp+8KEwp2YG8369pFcio9
vJ7kSxFJOcKl6EMTivn4YvNvsdAhYzvWmc411jPmp8koqdch2cIhG61KjgGqWOeJ/XFpCE91tfD8
B6nenRmJqaYce0e7Y0ITbuMcPXx+yo0oGBMLcAbUDoAPBBUBOBj3JMJPqFSPvWxFZE4A5VLeRJ34
96KMLpLTbjcyn/3L7sTwQwsseMffLM1BErxvlPW7Zo+mvCFsQRfx8ufWBcaTHG79Vd2HEGHS72bi
sKi2k01g+PGk9zyWSM2ZIRrIkPV6PVGtssy5tQFfvKDtjHvZOD4CaSMY+62IG0oK+zvVkwKrHh8b
xBUyU849dM/urYjSxM62BamvrhOReuzCQvtYCW1V59rcpqoKMU1TQT8Hes/z+bfxHeGC/lGtKOi7
cZYBA1rCTXYZzajj+Ox8+h3Ba3WuHmMOEB3Fpv4MqHDWMnWnlSUpnZs3l/aNGIJMVrAhaK/mmHBG
smqqjguAFV9VXOnVWdJ0YvxAagl9d0D2/KDK68DEKZgbI5QU4s7pDl5KOR5gMLlNaraxA9ZGIjVI
g2dOOg+/C3MQtGFk7bgoG1ZWKbiKA2iwmqD0zvucgmRfa+CLZuGOAHPlhnAe+tSDiMFCHpISAL9d
RXwzk/ncg8/pYao7OHqDxT/N/VL5i+SQWG5rc/i1+jZqvt09m/6FLHK3jrk7MFIdXvXVr0n+tDU0
QVPdhvgZ1610IOE/mz4K5PtmW+9P+lwiL7QACw0647cI67ijVqHqnVRnmr+4H9UM9PUltO2KfKhb
aaazFf/bE+XlzBERQcR9uXJ7t0hKd7NITXOUCDNQznmVpaNW9K4WooD/41i451Nwrq1ZOcUx95l2
wmvmlXEQeGtiNqlBklsAczLw6CZG++SkJPokk5dQEuriUj11QkG/N8Cg4/lPHTvS7+hekNfDlJFW
Ppo+AVeITr7ByWPyRe2Uiu4AKwWXMcnnnbe3yXIPVmtaDGWSk7bKeS7vQIe+JzEZRLUQ+/xHp4Ag
bEjO8SAJUXR5nDxD9xsmSug2BoBmC5dbLOnSWZdkFdQEgm5GGVtZP/KFzlTmQwK9h/oZbckGsDM3
zX7MsbEtbc+6ODaiIusky/4QXJwx0y57PSV9dPTFJlSVcib77bM36jnaNNpNWE1clB26EysQ5U+F
7AYmZrg56rgWcC7kH/Afx3PsrOOjPmFPlscARQGR5IX5pUDYA8h2hn2V8ylV2AnJCQ5r4Ej40BZ9
kzweBbCd36tjpMhka/wUtaKQwypUccssIZ32zDoxX6wO8K1KB5hITGBPK6swjMXTGp5GPaRA2ICP
2+O7WRSYtBdWgN1aomHds758t+ohwinCzST5Em0/dJGvYNFvFNUIAhaPmy5CMLDW+SaDG3p0zk2g
wQcVLrH0eLfBVaFQ+DBAJWMQvL30eMNFQolDTWTZU1aNh8uao0Ykh6PdnxV7niu6PBMaurlOGLon
qedINTpxxXw+UzpZPbRj5Rsahzv2dT0a71V+8xcakXjSKAkIY8+dWtVdaUmLMFTspTwQfuzGh32u
g/OcfAvObkyxMgRitCfREMjtrsio1wIMPw1VOIrAs0e6qaacBIQXbf8GrcRBoufRNiHC/B2b8mck
QL0jQvw1E8obOpAWmj+WxXyWRAEDisORIKYAuCGaprSBWtC+fDVAnAp9WcYVBuvQnE9D2Zk1OuJ4
GS7vpP2D2REj4/nryDy2kYTLI5jauuqJAq3qmg5lcE89ko2EGy7nJXxVKeRHpaVB0gAwIPcVrsWq
9DxQKICTZitujD7VAq7pYcQIeFUGbw2hWS2zQp3ppDLMmm7DO7ky5QGdQ/ymNippGmDA4xQi5tL5
9IugmtKyTJRUSoRcC9/THq3idq6McyAKrJhD5uocPIS+H7Con8ShDL7xmoi224EUNNJQ7G+zsH/C
EDOK8y5Nsm6R3WYWuTJEzryo2as2uVWrI96BM36GqEwyfaqwTQe7l3X3RrK5sphqHSzjmy5MdPzI
VnUVBCqQU64btSjeQUOu0DEzAtDvp7Z/3+5MWJ+3InMoF8V2ld94fg9ULY/bYp3kwLyHeQTcapXT
BiEQNBzuEH3YrdJs0pAxxqQKpflpZpzw3SMyB/tyVJqaqwFW4UaaAEQ9sA3OY7t4KUU3E4aGC55Z
rY1e54zivG/eoBjRDKptFsGdQEFiJX0WWUgJkOh7MovS6Ju+y2dHx3HEmM6i/xnSd0yQCGbtfDgz
+dLXwQ2jXDvaXrDxpsQ+EqmLrPM1sxp6LQ9Ad8pzHZZjshyt11exsSTgmmut/fAxIbPiw7IC7pNJ
+hz2ep6c3222p35pvpbESs568sMppUzt9HV2qNlu4h0zidGSPs0uAZVdqsJXnNwVPET47zdDGwKu
IDoNYcBvCeUV+eKqD5fS7D/hwvX5kw7oFsjcLSC54BNiqACo7VEg/n2iPKvz4Wy38A5U79rDSiG4
rg74la4G2BFPR2HJIV3aD0CkkO/Nc0nlHJ3wbJc5sX8UazpYURwd5eYgrL3aNRDb0c8aurPEGGwd
Db3YFB/WaoAvTcxCw0fOmMLe6RpV9xMl/3tMOlYeA/lABKszPwZXNGjyCLhXFQGgbaIKrovZ+qVr
UBW94wyf+5dMWA+4MvFDPiVsLHFe69CAmabcHVXJXu3QKnjRJAy8v8jtWKzh86C/yZtD8gN2nDXH
YvJl9oCBE0zPw56UYQqJ3PozY/Q69VQT2JegU8J5BNiq5yB0mZgvRph0e+hehLeSDUUwwFYaFwcb
yoEEIGYaZmpxw19Z4RINVB+7VlZDnywz/qCE8Y/b8HPom3a7xm6myqHZWO2IqMHo4ZrplpSyLWIi
dK1XbWJITXbmgIHFGOhU+2FygbtjeD6BZGR114DsQ5KJcE44CU39m7uIOI/d4L0NLdEl0JkB/XuV
HzTo1QF5dDpf7h3zBoRb9nC90d5GGKc8qmKCiqqQVUPlfz46xtHxdbojQGz0agBlj12oEoRZPrme
rHZPpxtKdQywn6DEF9q+WYjgvvCtvejB76Fo1d734xD9JdQmpM9Jw1vZL5FbWg3fqh2+T3xIInta
zp65W2eSMdVUTM+Hw2SEfC7JvMtsZ8q6VefZUJHKRamadTiF+KB5tHafcy6Wo9y2Q2ni2qZD80U8
ds4EEtJUlaJMnFdRG2qq35/UE7jBopPDRUo3yP0Hf8/g8mfVaoA3QVIzNKskYRJH0W1MZY2K84iT
Jp3u97EfVBxdc9HOyGXMsS3A5mNtlJp8ZJCmlC7NimKK8dD3XRxbTw3PdQL1jNsIwd2NV/8y3qWO
FipQlb8n7t83xKZwWC5PSaCBPFRF6+6qGF8LutILcwg6mt/AO5Y/Z3ybmyAXeH67JKzc0+464oe5
aZivFzFMGHTHxh4vBwZ8cX6YWd1Zs4RlV08K3WlnaoQlfiuQZcohA0DIbrvzmSiub4B85OFBFIk2
MEEn1DipbrBDlF4vyuQ3l+bNubblgmcGM9ZLgEDTrSQ5XsVu44MPd18xOsowD/d/TYzY+HzNx9m5
JZZrt2MbUK99/2PT7gRW7tT1r5TroYbyf8VjFSCzdfCWEsISvi01UA2FW4PP6VHPzD+uZiAcbBTU
YnBXgu5Tw5HpOtN3DSn3dkYO3l9YgNbE3eWQnZAXcxoA4F28Wq7T4KjnITeeQw1xpemufbRLwTwA
SFkgJVE8UhVfUSQGAovFpdDtBuWHX6iXoLypTimJ0E7BWKGjNxzInWYCMPkwvn5+2xgln8G+zQMl
EvVpa7Z9pn+5mb1X7HAFUE8a1uUmguL2/UDy2scNV6bsNhDCjX9M5gzyWK5Kcne3SNXG/mXQjx1Q
RVHRApCC9XBifyXFtSfqijDKC8tfX7Oi7s2myd/OWOgk7SB06QzgOEfcY8mArTSJXOpO3oaEY2Cb
jXsW2WHyfNiyig2MKr6j42NPXd+20B8u4uM4HHB2K6qdDsLYfT/NfCTrtuMhGPbDW9O6zTNpT50A
moWJFIaOFGxjiD7gwuC2CtYMCrZBaP621xSVJFmBZ1evYvPvLZG29+EgfkYaBkbBJ0XqO2npzt7r
0PhEJ9RQusfytTbaYNj6pnlOFh+g1ZPmc+GEHwjgIquzWW4O32BHnQAsnUq0HwT9PjenrnmG/Eh7
Ne5kklJ4tNSSEUy9ICUO31B34IfAOgBVgx6hGVRs8F+qUrAW6pS382/jJMBbpUqtXTHfQpZOjpMN
vePtYi1tSwE6FNsTR0eKdQzUaFeazUQkJ4bF+jhZcKiCNILP4EgxOAs1NFL23oW2Gab3Bhij+WK4
oMMyks1mtf0mE5JKf1RhqHikUbDm1UZFjRm0WDt4TA+6E9z5rOb69IfeiYLixJ0GHfRWVoZ5KEU1
jKCRgEdGzj6kDAu9Rqw44sa3VdFork7cRFYkKpVXcYmAVn4fm4/oNG2Fr3YqNvsOCz5Wnxm7/pn5
JmsGYtpM7e5+rmWQ4/SNZEI90Dxxk+rGX/oW/dJdrzu9YRRyeTWhBmPUsncS1cCe6/LBClEi41bw
EJwyMCbbvcurs1vUPmHPqt9d23UHBN46u9RHF9oXnv1z7ohwoYzBazZalXvV8mZjf5YNvv77GrD8
NJXhrYCuKKb+QPexkOapCUpiXABcqco/REZxhiZD5Zr+z07leShFhuzxrC0PVlyLsC0zixvT8zGW
aLK8ZkomgA4a8lxFHqgHFYDe6fWfRw9dMBblymbjCNP0WX1wI+zbdRuG0Q+Q3BztthyOaQpNRXeT
LsZIF/zQV/R6oiQ5zIc/wJo6FhtHKns5+tPvnZIoL+F4+Kpsx4dEGLrGf2OCflt+K+/S7xWD/ucs
XsrmtvSRY05rVyc+xWylxVG4/pzzn/IWM5AUfeBCvJylxfmLsSJoxqYkXCIsusbSUEaXBlNQWm5Q
2K3aUPdR8n3j5wIdrKtAWcAn3HtmWZic5aK5zUlpCSuBSxuPwKSalVMjG308YJDN1xikeG6D3bOw
9/VXvrndm4o9xmKGsvWdfOVYPPe6i/AggHIqS97OrAxMyu1aLgkEVgoZ64ln7IvxlhsMBTd8BdMF
IJPH1RDw9xhapZhGbtPOgonByTpPhjIcHSsUkp1sh5dnH3HF6jWFn5P0hnjRdmaZHhlsARq9PNvi
nJt/ZmcDWQVA1vNTAdCTfmIe6nJDvhAmFsLxs2OlnUV4eyH1HnzIvVrgp6eubz4Ion1H3kzu6pG3
Rl4E6jL4OWgkCEkFjKvy2PLfQQNIiS/3UM2pOqPn9ndtionPvGXkuZdeuXdkThMsKi/snpIifEbT
y7aJFaxxQFdHeO0tdH1g9Wc1XkoDqolvHFXTBZa2pXkuuTMC2y6A/lFLBD06PyK3HIZUSy2THAHC
fQWS0pdrkM33TmCHaGbW3Kk9i0joQsyvu8C4GiF8e6u0xAtjuCJ7lUX8PjsmwQLdyaC9nSRCjHK/
gXQZMrHsS9T/DIfrBfPn4QMxhx82ePt4F0APabX7eGjwwsmZZ+OgcRmT2fWwSXGYw/ROfIvRDFNX
u3krKnBhb5LN9Ig5kibh3b1hoBI02xB2peiXg3qstws1bHAO2voemw2gOXgpr69qcqy6cr8yygpx
FQX7L80q4weDCiYDPkow6kK0xbwX8dQDH4yLNiCn5K/PsyS8FiNZ/U/rf8Cj9tTaRGNvnAGR3fWy
2kg4egVGuNI06svWKo9duPH3sN2GXnQTQsHh9QMbc/6mmNyY0Ecvs5bBzLsKaDI9xE4pQzEwOOmT
aXeMF+JDvvgYXsH5VPWVqnXWzxbEs/9dfznLABnovxSm/Yq1BMOOyVu+i50Muz97ApArxeR8Supy
vrLEF++yosDFwJ9Z+R3kXe/gogwLjnjUc+j4xmSEA8WbB2/OYvXEUWg6DbTgQf3WZOrajvrPXqar
EhEA/i/O0pR3CMi7ZFQPWOxkB+t2lf/G4My1yELJKHqmwfBemLJBYqyHBnTqfx7aFBBgeutrwtIv
IJcJcHaAvKj3OVbo/Sr9nIJz8625+H/Yb3zCrPbg+2OrKB4DoBfIvD7f6cgMvQ6KE4kqz8cWX6/2
DtQ6oyjtI/G5mUAll5zAYi7Ogt3Vp4twuMWlV8IXzCkIYifaVmnGbbeJc/tDLXjnlz/pSW1Oyk9d
bzaZm4ovhR+LyI5tsZRpXx9gneOEPfff/nbXaTmYaw1j92i4LOF+lz49a8U3y8x1CFOrZjmUaxGp
KFXNqrE0+H3xCip/sIYTgljd1CmZ6MyXDMcwXrcQRtL1YdZaUBaDSEt70LZA7cgQVZ3GKWtxNSPL
UeHeb1vcog0hO4ala8TIz2LgH2FT9HImeLzP9znC+7k0aKlF9Rtj+WSW4JZ/yS48AbgvQg7cY/gE
+auMmEMCLG3nbG1/xs8qIhyywtld7L8PVbjRRDqBXqtuFjyxXLbZsH+vf9N/l/w5yo5kSMjBaiNp
ynRrBx+19hp7nLrUVtH4SadR886KA+tLG6L+PtbmYPSOME2Ui/nQyjChylEv7IESKNtfxtQD2LlO
eyE4HcboDwrbMvYLSjROgTz7BxoA0d1sshJ5lNv+Fl4lJ8u6ns0PCl2IQnR1Zr7qruUcxAJNmDYW
37JJ7XxiLejFvcJcLXStTvQA178NYl2FzzTClYczjTzfMijetmZq411r7gjfd1qmscU+47iGx9Eq
Ms6Z0J7+hr3VCgrplkW79rkfHZ6++jezzCRe70rKRiLnlGu/bLpR2Ru3XLv4dTNYL46i+lhKRtgx
b473HAg5COylVPHAJFWbELh39rPPHjTG3batYKr1BHwNE2TzefJ8JdaUm8VFpqsKTgeFoVeSGJ8i
13I7EcF3bR7MyjndyiASJDZ+YylB+CcpNE6a0Y0VKqDfQHIWk2+nGWB8lY4rPbFhv6qZk4g4iTRQ
qKKCQuRCqpCLr0VSFogc6ichC+j+06qGENvClRXTfqKGEoz/paj+kK6xvlSFEeSDWaWyL2RYkko4
UDkJ8+o2r/ckruAtnDJaWclfX7gz9KvDtkbU0RWV4df6bm1MJQiivb5imEYmTRV/KBbZaWa+qF/r
YOEjHBIAlx6ZEM2vVd/tvts6KB/sDGE4QhF0LS0J17s2vBh/tBQT9Eso+FKBALvvN/ekrQDYb5Mn
Urve9zcoTzfMhPYW7bClSc51NKqSl5eMGtATkIKZRj89UadcDi1ItpMlyeQdaZc5q5OeHcRD92n3
4Z0dkLJYnKlYO4HvNoZC/DvtI1Si4gNQXsyRL8hwhlK8td40y7r6yxZqoTseg2glagx5EVLkJ8QU
8KQxw3THp7jS90eK0jS9VSLSLFAXqS5sPJuXPIz43KwqkMZd0S7jagOY+gfdMG03F3s3gcoVWm1K
hHubZg3S1/FmaQnK5zeyNU38EwTtXU4ACbrSHaVnXi4O2igqZGl1oCHt4umpnfAI31Cs58KhgIH0
/kWTIrtMGJuiaXJsSvc+WKXbr7r5OFBPEbbXDA1XQ1yn127V0qMwtyTdpC8ecu6FQZE7i4P37nOY
p8skS6UXSBG0tDgd9Xq0RYPf70ggzuRY+ZdOFdf7HImATr++gTCawnJkB0h0q9L4LCuVXe7NpU2F
6INBP63k18/ap+M7/Z0F01ox5d/ACFPgntoyuizV0dsTXXxbOEXXBkJA6ZDH91e8BojWGASCbAXx
22TfRxnRrUt+5NgNXFbx7TL5S1vNeJx+AuI726yHAdPRIfbEJTRiCKy6od/AyQ+aZ5Oo8kTRFl+W
ghYd2pW5z4TSR+BhuTeYIZhCCBreZdH7ZTn0LImGaUjtZbvBJH90zAHCi0lAhmVd5R4Dl9sO6TYb
7hsqArB6IsB7mLenA4EO/qaX51/OgbieLYkHiVJjkAstyHXWEtfylX4wdEZfv8qu/yzSseRl42zN
5yeeUl7FitMl/1dIHfA1XKjn7nt/ynqv0GkPm5mhmH7T39GVG0gfhpvDAPX4VQUf1qd60XevkuYm
ixjSzeFRBI8b+papJ784qPWywVe/On11pFNmxbQdVeb6ZFXgw+LNGAqiWcrqkrQqdyDb2DJ2fHgk
IQsogZJo86XtaxSr9Guf0wcaqJ6TF3GWTWH7wT9TIq9uA13mIm0RtSgJ0SHd49IYFrcebnuAdspW
FlfU3CSJmvLZP2bk0l66hK5HQFJ1Wl56ZFhRsU+lY03W9chZJj/r4+3CfKm2B0fj9vcNHysULSDT
Zr4+TPn+TK4fTm1gDAI6km5U0UlCCGOUsZyn30WC0feD7UyaT+zCvhbFRJInaVQLKDBPwEOVTcwJ
oazXXREdylNFckfr/d8KzOgCQYKay4Wp81KITaFNbxsLcv8jUNoIOAT3J8cdtDB5f4oHoYNjV7pu
8nzmFQcawUyAxELJ+MyueQeMGFBJRYmHBZvguk/QAPdOBtHVtRPhC3QucPMPvGdxq2JgqHiTm3FM
5wagmj4mr0Snblpqs72I/j+wc27HrEwD2VjXpRL2+GfSSQXoq+WQSssjIhSOzJyX4RCYbIc7Is56
mzFOZoVaK6yLpOtgOM6yHLM0pHw/GRuYD8bVoiXLHS8RpwLXYV4YEovqHHnERurH27BxrX5ukyR/
NWsTR0Bj3HTRnq4k85Nb5XMWDxsEF0uOG2cOeUVMFO9HFmWbXBG7LBbrPvqFL607QNxyyf2w5TeY
rG7Un0fGijqnytmc5od1+rTIoQxmVnZbp64PIc2XIXYAhKYrKf8FE+uRNo3QOWVyKB6HzQ8YTOfX
fB8bQK31VObQX1rwFteu4nlZ4bnWRZovtr6c/CVy+n4A/3GZf3YKew6WnpTe8+pCUpHIPeDPMxe7
LZKhUEA9Oo+WufzD/Sm0P5ftZd/QgOCEMxshXN8bVY002CLgLheGp5EO9dLWjxSLRkSwjcAwa+k1
JKrkEq444LeVD9cnHEgfN8JECj6KS+s4yjPb3mGcC/WwZJa/O0FpWNFy5Kbzi4w08DKdbcgByrZV
3gP4fi45OH457sPbTRlddfEVXNlTFgBZTASdHjg9s8WWNC0/6SIzM5pjeoAmpMrBdhYHZXNInnCd
w+F+3n5D9fWIMAptTOuHk4j9CPmAL8J/scDM1PGO75QLiLIAWPrZwgsNiaBnN3uVCQR8vvWMc/Vo
izCKVHLFAG/LCL/39xpOKybx4FqT1L2tYNfW1uBOIvu+LYAashv+eFQpTvp0Gc4ggrONAkCz1Fe0
uy4TEQzGR33cwSm4UL4TXFhMnBrJJKaIsnG01wBdXzRMoRpL4Oj2jenGwjALy4aumbALzThk8kkj
To+oJonFgwwFcQnYAhmGebtpMfWnL++tp90e6bl2WAfTsOOMV1aZ5SXM6uxKBzuIx58EYsIBqjvv
61xrhODWp7E0iPMMBA9N9J06C1Iy/vAQWJ6VzWRztIzbm9ycaB7RrNCZpe59B8sOjcfdMwspWTVG
nqdGhmRyiuCybFddT9KuF+CsUPilk7o3c3dCHlYQ8AB0o+1NHVSZjKsXP1nbfS642Mzq66Sran2T
/RmINGHbA5a9fsukPP5T5lElRdFFZ9jc0YDfUMDur4CbpGpsbXtq8Ra8/u3C1go/NnMfdNeknnLW
7lt9eiGA/yk5o+KLRt94CJj1FTeWDvTa8qXvlr03YGa+0GblZDofHQAnCApFjgv8JJzJ5A0hJsRP
sXCMbGdIzPB37VPl6+DYGgQyEjSGMQJG/bwbqmp1LsCsJ9dDfxrre6Z/lUsrNivO+W97oTIyKprl
utfrB9HxH9pHQ/Tm3kEQZE4aIVu6crAqokIV2RHbYF0ounUjkDbrcdSzms6E9CCp0tUcL5+faczc
XuyD9cUKa0rkl0Ax/QslfQy4/qaSWgcKwXkd6vxlxY3cEYSg1VtnDLrU1SV0fAsLOQqMf736vFFY
xrucdc8djkaiXaFGH1wSgk/r0rstfGnitL6L2w2+selXgKEtA8UiP05qP0RdhsSk7qwI9mBOBmeJ
63ntpHApbc+Il1hAId7VCeOpLyioyMWKZc+CRL9Wtv9d/qOtbRnEPBFbG/AG2UaeKwJO2qg03O5U
juQ9D4EVAXtkxg+EE9o3KB+VwijGRVHbYJlIvvUIccA36BHzxl5+y08oHPW1A0j5tXV5OOPdxZXT
Qg6yvPlH2Ph1U/bpYs7C0xwI9H+gpzDn46WaojY+M2Bw556IV1Zi6cPnVQdfiJX69cfW44Q9fHl3
WOgOQkoplpYLmJJzdQtKbHZft3EXfhQJbK94CSTCQ2P0RmgHtPLTxuZf3DXY0MTOuiE6SoPhSjMK
dyoqOX+0+aenJ+4igCxmHWNxjmqwsgyatJea9slEp9o2VGdZOC+Xa58aYDGroRWFtXh9IOkJMAFb
Tm1jqaZYlyL1T9Vrb6W+nTFE3k6SYhOSr3a1Z2prN4BuoeK5hmq3nyX9OaUj54ao3/lNtwtNWUT4
Pw2f77JzIGy4QeOcHlkKQd4C3SdsWijX0JgpAEvN8NXu7+uQ0zsH/m1lsVIpyrQAaofuc9IQ6D0A
Jy29QxlT9KrX/GeISA1C6st+lDj0PUJvut3C+80X6VIYrcwn6qoTyYVzra2li2hvEjw/rbqwG9tC
/s2igw8GZ/tXKyJRjiyrlE74KPBSA6Ed+drq4CZae3xZGtBkUGjFPoS3EQfVG2ii1xEQea811Sgl
vlyXaZtuQeV0cAfDNbxhSrEZDqmPN7PJbKscbs3HHIM9OJVASMSXuxcHyIoeruu7k9wvxNOVve1l
FJEgKBXgVO5lacFthSiAuNZrNZ/OdYO6VLNvtcxcrar41Av/h8apFMDEORO0WPLtyQ4Q8CvFjncj
XkazPUwV2PKOyFmsPvP9GYRcVhbcY7LFrjUAZv03MuZPYAor9PRHJrN/JgIYX243GNemMHN5JwpH
Pn0VMYKdAJMs3f77yJ6UjwKQ2AZCIbKaqxnu3RTTPlODLkQjs4/tjdyZYLqBJYO+JfN12HI16aUP
eflkckqUu6+mk+/fk0JwSrdkOS1OVxpd440mtK5wJzGkSptrPaMwlLko5CuP7P36+JseUsbGIt06
J32BQe1PQfrodC53qFys62oKgHWtElbkB2lzQ3o3ji1R3VY2/wTij/d1r3yAQuoddQWUOGNkb7RW
OKz0Z7M0Tqr/sFmeSsEigkdgnS90HiJhE1SoRz17ufiZWWnpNBKJRyiSmiO7Nz7DpAhlzC5v/ffP
kTTg331FdlpztTx5FitfJ4QdvJRzTPWmxYCBiGJ6KZm87Cam1GjSVNIKH+T375AJW917oOwzgmIt
wrWPZtO7KGMGYPrTNrjwTbbQIwCoBv8NyfK8JeN6OjlKgNnYiYae1K/fkqWncqrJwyYKwlqskwzL
FlZ1X7Zk6BL7ANM8Of+mDTCODEZLAlSemN8CEGiuYgOHWpTu7HYwcHFt/v90njG/Wrpk81wJOpji
GPioTHVVEIIbK0nXfyiYDqYu2yL3gTl9Ki33OeaGDpTtzYu+e5jfmL6vDiL65ioKfGWKvozA8HAX
zZjLK9RwUVNcwKnvcPnIrZLaEX7wlsNwEvTJpZRUYb0pQXoGNacYqxD1RJOz4+Rs/mhWosfGNDx5
U30oXqmrHYGDGQPWhltVsYWhxCBa3z+NoXTCh89bU0rRP5lHAKLb1vFJbTIPrACTbLmHjO8WHtj1
qYMNfLDL+Q0NCbDNyZ4qYk59e3qGZsMe1XxZP1D0Tgo5tYFp7eiVhilNpi6qwPbuBizeMSCo8ALz
3nvojbM+9JUpcKxmdRLuUg2JkDChkF92ESvfc5K1Hx8HMr48tw4mkOAaIvyL3VrMV+RA2lUt8Zd3
kqKJeCSo3MSwKL75JOEI9LYjrTz8sXBCtA7Fl+agqD+1cfGHqIXwqR8oAStZq/DsG4pJNPGtX3Ri
iXPMKiSb+chxQsdYWBzxSiEbHYoGfO0ExlyO/aa8329Vh6P2XxmJNsl20r1jlp0rNrmVbFve4EoQ
MnbuDZ0DAdmPQ0vUegv8an4YXcgM/oezbbwNWbf41+RqowAgvDKYIwgl4PkmnmGHjlJ4PKLbWRQR
CDwRtuhRR4W1yjWF3gfFUABaFQ2rSu0/15/Lgbsaz8soGc60pRn4nt9lj3GWhtIsxsT9ujVMhMQ2
AnhcxqdhPaLhZ+/ReZqKiNpaj6/BF5l11Krn+nZbLcDIjMk8Yp3YAXcUoePC6nCGq8r9K1Zvno8O
L4JHr0ODgY+LqRRZFw9lzbxZBMh+B6gqMUCFkcT0gFtuaqS4PMJFyWexJUIvirpq9wtmTj4NwIhs
Ykw3fojMH/V0FU+6zzvpsfuT9uBrK6bZKmyYhhloY9+eH2CEDnlioNmB90wnv7D/NzvJ3Tda2aQe
s4ORi9K4s4TtlhWS95PiRgJCHWzu5j0oJTdZu/SwSeErhkQ1BggdzPI0cQqSOOhs5H5cEbtIAjTw
ezOOxcO4s6XvAciu68TU7KeZr/UBgcejYsPVyaBWF8hWNj1e6NyNgp+Efben7xFEAYQmQdlFP+M+
FTHROcK44C+rMcN3XBNeqcp7Gb306Mx8es1YUGGcABFi9cc3Gj7OAmcYc1x3npvsBo2ME4xfQVnJ
AelobnKnJlMUkyqBGc3eDnn4Jkb7CihqIS/w8Ed8SbdCYg0c0J+lYxWUmscL4/yNy7J3wWVEOAy2
G/2cr+/b+5/75G1zv7UNcvGGv+JL+qTRQA0Gj60GwvZI7lbzTVg1nNYcLqZ/kuMgMe80+xriQT5o
4mggx4H5vf4irw9TOtCiZ6tezt9dBv2S90KBT7s5rc81mgDR4WBCeHpHIYA+28PXI45B5hvx4WgO
MowsTdtByX29ZkH/+z4jEv5edrPPhig2AISG5rKF2WX8JbUryK7GqJgX1fm+J0l5OwP8zNXj6TNN
FU/11iuBQP5ZEQzSJKVN+Yy3gptz4/cUO3E5uyq9bEXgXIqrNSY5q/PFnRWGTE95u4OH3Fkp1y4G
XbSBFfItemdqG/7SIWMeYxNsjNzlOrX3ALKqnCI3OFu4/0YN/BJf9mBIUowuKMXxrvi3TiYuXui+
bbH1DwjBV7qEfAPK0+Qa8jOGXfTUo1jQfYQNHz/70WCmPg2JIqnZHeShctNf/wtLN/AlkM1DBfrF
inXJMhe+BfTnszPTz+dZdarR9KDlFVmixFoexka4oCIdV1udZMp7a6L3XWedjnG+R0J7xdb9igXM
yrzEK7kaoE95Pdz44pz147YjcpQ3cp01xQIhWVWtqzDCzNLAypKNtuo1OfNWjRIxzrTZvmEazZaG
vkV3E3Tcdn3+BxcYCdXw3jnTbvWGU43Gt9aGMNgcxsIKyb6+KFN7g+dXf4wdsrkBkn9vMSHx6Mf0
dDqEogazguydblyWay5685znSaxXlYpCpEtz3tcbABuNN5RUDb9jv4lf9O33R1PFhuWRfw9lUa/9
HR3PQVo1+kn30d/g6irQn9RUR8Kv6nH5ZMr/kSeXi3WWWsc/F+o9zNsY2KNIKIbUxH2mMMa2SxQ4
VFW9cmz/I119ORu520TzV6+4do6nR4Un+KC5vX9bzptjh1p21w2CSPSJg15jRY4kxkMKjDyhDDOm
/QCycCL3UifiJyp8jVmgqSuG5yyvsuti7hnF6sxGF3JEQBSarIB+FTrwqX4nOvtKdaI5u7eD7w4z
SKTmafidA54ogMK2Pj/wgmIAdCCk+GxxHwbNpqDktUkX2FZ62g7E65BRzsqmBd6u/SaThwlMB5O8
VTwhRhpQHG1AOeh7eHudeW8uaKb+Eq3kIdNqWWCUFPKdfwzniccqqGDT93oF10WikS3dCK5+KCU1
p2sleP+2auDYIj58MN3owzfd/zh+pQKWswNX/axeRgt0lUUY+MfVYWPrnYzfRFm1oPPx4YWgHWkJ
4deeIVvKXRtfFENcbuU/UO0dk0AFR6A2y/4q9rmk8fSVy6/fUAeX1NuBQGDcEm+/d3Y+2lZilBQd
AGf0amFX1Nxf+Re8Crk1wysy03sDt3ii+P9pLbqG+t6KAp/+7I9troej9iEuo/S3h8+NhgqXM9b6
+rbAl3WPkZaHiA/zVgJRFDnwJacRYftu01rcjseSmOwRodUWdpEeiaivfQsEwmrMLTiC+Qblza2Q
jtZnTsH9A58FPNiOpXb6VOa/ArcOAZWQufiFhn6LW1Cs+cjoUaWzv2mo0BISGbd9Dx7ztgJ8KkB0
mxadWMlsOhwmYvzfoC6oJBponGAZoNI0A/wt+eXdUVHDz6BbUDLS0NxiBbx0fwhdeuLrl+cBnUac
64R962M9h8U7ES3vwh3NhvMMvvatNthxhSx3fyLLd74G3VmIu9apv6OFXEVvF8+s+bbfXaWRmHSJ
IYieOv5dY02EHfhM47aPjh4LiCbRn4EeIRdg1UKQmoOzavhRat0Ioe6URmxPoIch4Nzb8tk3PgqQ
bpNvxj9rqBNOoGDpAUG/AV3MgWfOjcOSKSeOcZy776RCT6jDolecrTdX58xXohB8aMs11ImPc3rM
Q51ASgHncubPYxYMO/9WgkgOV7WYJxz8+BRyikwyMm15LrrBrR6U2qxiiF/3IbGTVdi0Y0x2641X
KoCMq5kYi55AW6u5DyWW6cb/s7gZEuvxU9vQ8ODqfXJdyI8k3Pg9/Yi44q7KNS0MseJ3LhvQqu+D
DLRxsGGNuLaThKJnURqO1ejzfpO+NFPJRpbYNc279u5lm5GQQh9VoII50qYEOk3M8hB5+Ng5CcAp
MsHD84iT71QEJP4d6HmdUjCmra00qc42a9UnsGs1tZwQRMA8PB8JZQ3AJFlfqcpWR3DjpaPBrGhK
JA8xB6aQPfp9uDLJStqZkeWZSGlwfcBU39ZZucTcl9kOF58CtvWOJP1cY1C/zThj2+WPYlCfiik9
nTnJHeHpdUQoEB2LFA7RSPKQ4AArIiILf3bwyx+Hk6nIY20+KkIAUS7PROdJJPpl5dT6gdE3fGgn
O0UOFyZ9rsjvUMlO4bGqJzFhoDS3S795/zDQPkSroBiepFaHCA4FrBQyWiSZxaMeun4fD19Ap3WF
duqSBy/fzSTe6OwqAmeQ6z+U8p8rmQD5edh53jEu3ZIHcK72pjFCo27crTZUJz1TQPV4Z/HCffDx
A3UIjkcE8F2l3AidKxkTj8BMJzcjoBy2i6IBz21egvlsrDeRzdxDi3wNlQKcwK/BZHJLKM4j309G
jPlOM7xpslzw1aip48B1orsCEWJv48FHeI342s1fNxjg3yhJ5NTcR1/E31GhO+QSVbIIeREuDsQz
pbwSEyTde6WmepC5CBuTN/d+PP6cdXjoEDJRe5IZdJ1mRYFvhN6zewe03CNx5XdLczM+wo0v5hCm
0tqoUH+HHEP1cVD5queGAb9wjmON7Wwr253gzRvCxIdXsXVv4Hw9QNsDgkxySzI4pYsLZcEkPTBe
QaevrXNywT6ce3AWnunNXxTekmJg9LwRezr0PID3cOcmI5YXQ3MABKJghRntdTENNIjhwbqhhDjy
gZp4KL1Ey9YhZXw5yWPmToyHe8JCEUo+s/TTdBf05JmHTqLIa7dk0ZtNamfH+YnaT07ZUf0+ATBh
ombF5QCxI1jz+0CBJ/Wf7WUbYkzZAylYdvWBUGWpLnXv9lhcwwuszX/RRuIzlkq0pnc/QqZVrWwL
waDPq1kzYfrrPu6b+sAcoe/lS28+MN1H/y1Knjsr6WmwvKrLQXD+grDc9fkh9SZ/96IiwZGG38yH
56w8e7928ZqrwJ4TYNEJ4MS7dTI8gmzkmaDaN4e8tgo2lsRciP3g3dVmjyjPZWwO9OnmYcxuPytm
0ZfE5QFNnCYtcB5QI2cTPwJ4kdtIQtbs7+0FuQPFioaFAtiOdE2FE9o7J/vyitHPg8gxEm//bn/5
29FmABwaf33l67LdM9wzXahjBl+swqOnaUmgu7TsahtpTk+I5yiLKV+veWfwRo1tbkHqWP3BYtOg
7hrsuyZHWGyLvLwpFbv9/IIHMLkH+F8pEvRpdDefOLai9AAoafqUsRD/wc0LnbCfyMfGSS/48rPi
Hd50Sid6RkkePoMVO2Y46l9ANH6xsvwjLgUZplpktnDvkJd924/QXhTpRQzDHJWpB179p82E7e7O
wWyZ8KgSVyB8RVG0oygixrBf6TbiAbc5Hh4U7G0ewBv6PJdtGnyOw7d1J8ZWZCAvDq1g6/tweITP
8gml4neq2WYIt1HL8cp3clcMylvQ1NkakpY7JT0/MJrlpCKcNcNViMyOFFOuZFPva9DD3bkFlzq+
137WeniKnO9I7NeBcd2RBrE2hylVpICIO2Sso2E1ojk3yALl7TfC6ahdTeRl1Y/Em3Md1mkP6wwc
OMLHxnzGyi5bF7GyANRM1yXN5uSK1b+/S8SoQfYUJUnIqrsNuoQjS6mn2wzDsb6ImM7ctYn5RsOV
WI/agHoCyEEI28F0V77/WU1H69lpcPTg5PTSEHOICCw16ZRWT3cOCSsVYLrZr72KIQGlPBXfTcvn
nZt0NsJ+6qyNNSMXzWGXcuazsiAfC9ciB/xlpwowyhuNpeZwoAKV9/Jm5xBv/0yP2H9g8DTwVcHE
v60UEvGrrSHdd21pwp6WSDV5Ad4dCttySM+7wLCXq/TJQ5UOE07uoOaxOHWiyb056pKd48OFNS8S
mrGzBV5nNQcQfs2PBJSnjpLlX1lJEZM59lRgXJO9FcgTiTF9BKaWJm52ytcb8BbGr8ZWnv62LClg
l8GBAjHtMCXp1XmdYXEHBwUnI7LjER3Q7c7QhJd9hnXPqAsJ2vKL5liR4G5IUT85MCNhsCl1ZlVH
InIeLz9mxgTyNbO0JSYKY2wO067rojNv64pGiimS8WeQZm87XHlYIvHwemeoXJKp02/sZAkrqalf
I2bs0qgGK76Q8jWDXYYbGjRn2jyA82yBTxB+wJ3NaiAweHh9j6/hnhyWBp7M4XnGG4qkp5s57RGl
VBbuFpBmdkVoXrfLjf1qMAgPslVQ7ipSVuyoxmVjHs5f8LyBeD9Oy5OlivfXZmxz72cGCZrl1zQR
NNxgR0OUKp75CjeMKFnk0oEbatqxpqpidP2LC6CVNOkuSsZHH41ZGia/p4M0C4S5ZM1lCa1IFqVJ
WsmiojLeBiIapxBDwByuIQyn6YAYjyNMoF6D6MCTc3kmsk3fKBQGwflOVMtl1YlaJIlerEh7HXkz
4nzM80ZQ8j1D6bf6Kt18pv1gqPlhyJT1VrQRml1kYkgCOAGG012shLynXBPhmWrUAm9m4dNGM/d4
lv/bIZv6ZC5L+8jadPkt/WBdC28/LjymDwLPoljPKcNr0LL5dmKfpBygAxeD2lso0aWpLLStstiv
Xt8YM1Lnsswxj8SwM9TNrWW1MMfSvsQhEbA8uSoUvZ01ZO8R6ycjBacB7IfUSQCBkKTHt1dSVEKr
OZWQILR5H3IoN1J0LVPygDM1vwMPnSl4l+xQFuocZLnNhVUKSUKSHZ6RRObDjVZB6QcPUB3q9BZV
hdW8lr9wd3P69io1xr0yKNQjWbTIIuXtUSllCmnMfGgl0S9tYzUQjZy8TTyuHeANroMQ0lVikC1f
KbwXqfMvsT5dt8yr3aFKjEKlKT7dcrnDnd8lnO0HT1hk1ZfhZ5Uwpe8zV5SiHkUVT1/iKizl7JWx
k00g/nRbPdZsTuQyuZ9iCW97lWRunTFNAw/8DnOYa+fGUBwUEsc34YPtuF8TwErpsYl7J2M/Fyz3
FoRuQ477ZAACfYkfkA5A4dcAkJS8bXFUsO1OuKiSodRFdKpYmpO+ZQ49+pw4lHgHoUupFHlSgA5j
V+h4e593M2iTTlHGfWMDjHkrnpYzXTU1nTAhoR4HYQCE2Lkj6YC0N68greSaMa6Os3oeLkg5LGtI
I9DykgvU9bK2JiSvmfSpSEa2ApiP6GcdeII9MoWpnSk7Gbgu/Ai8+q+VLvpnAJRt8UGcP4wYicWA
ZUSnKefkzq0IUh1+0wcuqIbkR6itEuMsQFWOHG81dFbcumZmHBQ+por0aU1wPb32Duru/5vdHag+
GA0PP3P6hTzG6xM0yVWV1S59aKMIUtDBfiNAkb7bto2ANo+NOqHbRYogJfeyxShbGRCPnF6LHfUB
UFHYyqTTkQb7BY2simzmXmd7IAYv9xilWE1CFT9Jz/FoSzwkhvf6DMLsTPlQFKAb/L9lFOEXnq+y
mGQ9aVmczeFZyEMEnocLAabljr1qYqnu74ZJtsJ7hELYqJjm5ARRyhviSgeJgQCHAXGm5CGsusff
Mon3n3LXKSOSvHv0OWNzVDokryXWDKEIMY4Q6ZoDsC5yH5WUwXs4wYlW0Rg2jbYVfXkGicayuPyP
vcdr+k6cb1PSlv6JgcMQeO2ErgpKQmX4hGZLz9IPzt65wsQYgPVsAv50GDPEPIHaPAq+qdrCzFxU
dnJQqjx3C2JZ/Z0Hz+NoRoYwpj07YRKWkVLbNGGiOcRKI8URJCtNOrhfGCoyumbMN7I1PJs67q5K
kaacpxIU8PM8W7DywEvGCNiLnyjqGL0pmtw8idyl0WPRgnTeWytQywHWDEY01eb4iZ1YxxGXOzHj
DE86BQWWXugxqrCeB4+OVTBHW7nIxpl1x4BRKYHKUvHeyKRtdF1yPiT0BQDe/G0R+bLLAB4COdBd
rOdFLt7gYOUnAcUF2tgOUIRSwUYbrVJvck61NmSk8x15ATwZsAFsNeu6iNdWRvlIBLNd/vAKdQM0
Tv9jlkDZOkl06kt3c0ZN3CAAwur2oB1Ewc7YJ5M9WYnNiTxLmZFppVBwKMjRapHlfYFgc1dfwrcN
prrV246e9VodWeR3dB+BRm8kmp8nCvsGEkh7BZjdc4QJH9vQhKUqOOeHQpdsqQZkxzHoAsKBq/zj
c9vzuWhoGAKz7o+LmxaoEo9RQlNZ5WxOKdDa0ZitnnnW3LH40QzZ4yyuAEP3ZNH2FJJuLE76Ufhk
jnuOaTUoz7244sQvfA7ftRjK1prAPU1onxXRzKBuirNLQaObxr4VkCnlsHZVEX6+y/shOPjWhTH7
zeYOkZ41Es0x2+/nfnd4YgrLp+gZMAyf8nBle7sqw+ocjmIW1OmuMxTvEj2mR6Gk0klw1HHEHaYA
8XPNSnolRojAlu+ww43ljz1rIbqgnJwLonroTO7fpnRilECNp01mVItDFPq0xkAOmniOp8aWEHDR
VXYccmWY3NiBLiXDC9E6EKLlX86QK2OfClLv3LdtKrLzFOh7GFMbM/e+yFfbiOJmN6wNSli9vuEq
ZL2erymBA94qFiskhAj6MrmhQd3obqdzBdSyUVZLrrCZ1lx9BQMaQVcrf/yh33ug6JGtd2kROBHM
+sDkz+ibe9ljxxfEL6rDvCMMJDi6ggFjYvI5Ng5tdZW5IYLwTz6ddmOp58HcSIi1d59l8xFxfubU
6Wo/3jU7XOQmdp3FUNn5ApCUysA/UoB2UN4IWntougSFSzbqcmIjw8fHKA9XQ9Cz/1B8F3KdznT5
VKQBOyxmbEzMaUAU2HFJubecOdFgie6DBtwK7Ma5oHSRJyePjruSAjmNHe+kD1xM6oNcjW0XE7+V
Q2dSB0RpcFN8DcokFPMqx8ec6uaZobIWoOojkZu39pERwp81i8X91xeYjv8FtnJeLNELMgDyWhOM
jSdkq1jGti+A98fupqSLrHnuwc2w4xabisZuPTYG1X8YQXsYNBgvPuenzC/cKoPORknjSHGWwGis
C/Xep6H2Qkiu7qdywQPMug67pVlASzGnOSqhbwvG/xjyFQww2CaJqoVZnvgZ+UJCbiyKiAu0mszL
HPDahl+2+k4OkXWmCN39c6Y8R2k9zTCc4LPdCFlWbEsCR+btwr3+HZw3BwrQpBcVfUyqN54BroBm
RF0o++l6l8Cmg9sETE25mdQYplPn7pRb8gGBspQabamdnnIWjeZk2A2v/d8xzh2fhXW2lpOLktvn
crNAJtmgJ0nkoSnXcU+VLaLgFTKhUP+MxljKc85d7PZ7vIEgL0JDg07hALyBZyu8MaNTcBDqZQ0j
tIMWmIjUV5MUTdw/QiF4E5gGGyy/4GwOD1GFn2zaOrqLDs7dibtTO8FHIEe5OMPZSwXA9uP2pbIK
xKbiYNgWlHqZqN9MqEyZ37rIcBCEne6Nfi7j+zoPKOf7/Q9GuPz7hUNhvf0FqA2Eukv/7PpAZAl6
FRGZD6P0j8vnol6TJUjbskRRPh64m9EmXC9twd+mwm+UmEG9kk6iezTSz1FHnCvsTRgIMahNIAPr
uhN1n2gIkORlTEc4g+Q0HkMQMtajdCXpdCtJx1P6XTblYAb14CzLPanJFv0WApGOdCbFszU30Ml0
73rucesp/Dv87UfTp6luGrqV+YOuYAuSteKc13n3Jqtfrbc6fLNzH4BdB7gMRFz60bpSxLzgMhsM
NxwDBXxCjAnpRl9dEHdEGyByzBOLWuO7qMVZsxtKRiHbsSdZ978ztrkoU4g7mrWpl1PMmAFF7KGo
+uty/behUQhv43m/ngdv7t2HIASdbpjjcKjYjudPFoTb20Zeb92BtvCw05vDnawQiX/61so2bD38
K0Fs+ivyxqBYxHsr4ddrA5NxxysbsUD1eLM09a21BgpU7RenKAf6D+I6HuOdWld7K0l46MLZWzbP
5Y6SN///PBjq+AM0JFjWs6199pNyGPC1rFyHiCjnDKydRGBYpARNZb8HoZh9TgtmNNyT7DEbV0nN
CfK0n5h1URYE6JwQbGtgG29lEuW4eBj5Tcf/5rzfe9RadqE2GsqT/YZ6UhIwYh3UxaHNa6lSAfnV
6vzsTxPhaJRt/4Osu633B05ROAAQ7VihFoGWnpxYdWGl+JGmhyYtJKoe5Pw/6JB2lJV9VOCaz0Wb
ZqeltUPpNRIemSnuSOpmEttkEt9htzacC6bbqtvLr+HDjOpse6+qZsz7V/rTt9VaZ+S13gP395a1
Y3jtCJag6Ol79v0+An2DkE88/IDidNNDAT7BVtB9Bkq9vn2QfqyUCIf9wPnfCMNVDI4R8auTUcIn
TFATOuqC2J6XXurGbRxdS7ovexvjEtzr9EeZNiKjnl4bYDQmlD794ZKwtmuVXgUzWJxBREabLd7Z
SiVXHTvxNZPwXTR7ZVLyQJr4waHE8VkopeBsI7rG4zNQnVEgHyQMdjMR641BJrPe2/mIRiBglBRT
1lKD7/Rw9ZJLLrtEKq4XV+4VJhQgzYB9r0FXvRLdRzVAP8QuNrSrHBsr8xrhis8wYxi+/inR9YMA
FDDKAtVcftrbpHMU/O1XFFRFO2K2JiV1B73U0Gg4OoPsB1HAhem/kZDbwE5ZMiIBs4VGVx9iPSJm
ud1FKyEpr51hVd9WjmFRqJxAcJm7eTQ30rqD3cXbZJAZx8QFsFsAY5o8uu2OUp/YKk4IuI3g2hy2
nUF8X//i6KJRefC3T8YlzD5g5+iQdQp4mIDFnIaKIWFaWm6N7mIg8GuW0ETO0mkzNdXwtHbywE2Y
db85dcOjK6qWOWkFGkOMNxZ9iGbd3xjRbBwyhdwoCwePY4/VUVtVvdfVAdYA/KnSm4eJVAjb2QU1
iaFqdp02NQVyrRrC0Ds6FYqD4uB6YlP9ffYx+CAJurPPevcH3hE5EJLY5NytQOaQH4Y36DqYuwUT
Nt8Y80283wOgK8Rh8PvJ8rz1lrZ9rq1n+yMR2rN9JwJ9LQe+ANKAkuZCAfghdTtlnbFw0Si2YQhU
xauqKzVcWPtYxbe3UVyaOSNIFfgpohd9aWLX7rwpohukXBAM4ysIfu2GbCOYgClAN0VOx/Hwvz1t
3kBiDmFlICmI3yYtIVvD3lXfm1u9DWx3XR+gc8Fua8ZeoPCXjY/w0VPeo7Ba3LZWb7BZdcVNasWW
Qot0B2BcTzuF4q2i3ccUK9hfeNyj6WQCT3GjrTNplBJGtrpcyY0wJfZYthKFzJulQ1J95O8HK6w9
zkun+vJplvaPCLlCFr1UpW/y3r+brhcxHD0g0QJxTL+0fJ4d+CrqIi4z4JSlOkaUzu3Kh3YNHfJh
NvZAErMReoIa5XQPWDJkyDbP8bxEkHPoUVGceZ9D8G36zZrdAoZeixy/7wz5Nc9nyFUQ+S1sS0hu
XZUT2YnXLB/Y+ePAb0f5E2tOdLkwQsakFsHcT0n9nifKLlljfBoYu8y9yoqzKkTLiPETaqIRvFmU
tS3Ad0dCMrRgG80dqZP7QyRoGA6JEQw6anTw92s2udUrRd9RhJvc0xZBXZCZtXTkqjeD5/BvkKty
fhQ5tQOf2lVjzocqQfTX2W/lq3chrriUzkViq8MkYu+ZVDV4QQGB25pDyKdus7/mK0ErgeTXKTI2
jq1n5RX4KHzwCJh2yklX8vD7FMTCyN2+4V6sTwYwVDl2cIJM6iIUzCFAbsLSzAObDb7UDKdSWas0
JKbF6af7JJbyIWWxLKtwX1aXumulHeDwAGmwOB/vaLuYsPVRX7eFs6jpFToPziHIvgoPSXBZsIdY
YuuvJKPVbyGwMXEfwSLNfthfARg4HjDeLkRi/lJ6j8w4JY/IALuOxVyLLuErfUwNg23ha+GCMxBL
Mq780fwD0BeexlkCL+h+wAXDvNO1ONrcO9UW9sQ/qP6eJNqZNr1FYzbbz8P7HG7ip/oh3l6Nd8cL
B1+PICMSHdffP3T2xwoR/nxVpl3wwh9Ea5q16iL172bk+HflhTqx+dxngeemyqnX8PFtxk7MgrVp
nk6o2pyPmf+UUEJVsQRv4qJvzK7u6khGmMQAHFHBs7oMUe4nQ8Sn6gHjylQrGCpZivSDGQOIKZpf
NTU1ABgB5L8EEL9aE1glU+bNfboNopPeMB+QtjUeKo5LK0bPtCQIxOhs2MwV7abTmJZK1OLHoeaB
GVMH51+3N+rp+D+LubKcwsiZ0QVNWK4yh8bCiERi6RBAbPhHz5SDi5TLOn/lTudvPc7bz/w5ABMY
paLaNacnLt/xmSFchO33V/E+IAiUfrXDjbjwpSozQru7o3t8TaEc/bMNGkeGfiG+udMfw+QRFpAo
5qOdHDncC5QE3B7m8y9DO1RtrkX4+a0BKhrPoJRLZUdW+oohjaD5LtuvtOVi5QP8NOYQ/nwhkru0
trlNvV/36lB/QkFoOvyE7EhU/F6FDhYkFx6sO+0pRCQCv0bGscjXoodCgWb1HPP1lwne9EvIPwxf
JrQ3vD4qL07U34x7krKkQ56UKVF4NVDLRsQHiNtUhU1DSlWFdLxDxFRqda534KZ8LkHOaEUuvsw9
8NinNyq1qKtoA6ZGtjpwwsUpKtNB1sukqtaHXaDfu98z4KeEiKv8XTtehdkAqq9XwMlhn609P5Lb
cofsKRmOeYUbCnhtB1pfKrhrELTamE3xy8VVD7Tc8wDilVziAb2qiRAn6mgMSTqKNWLARmcWLnfE
jL9R6N9kYTCPxmTgcDovOxdo3eUYtnwnHRHmAZTg2JSz4Crvtr2RrcQ0DkCZnEaP/2CErbFM7xuL
sHhxBjcFpg2aUPKLuQoswDij2q26YPUTXqqGFke11z3kWL3Iz0pTu0O//2GiIAuj9Vm5GyaIRze5
ragmk133MZB6Tv320+NQWRJuER+9wCB24wRPVWNITXqiJ6tZdY2ZEkcvcj6oKMp+c6jqSU53B2fG
Mhe+ow4wd5uGgXyC4unsarUVQMYRVaqSTmj4PE/Gpek244WwcByKgHaCKKDv1FzilcK6W7pnqD6n
z6jsjMRIoepsQeYt1T/kJmDyOvWqi2ckMZ50n7CMcUtqXiy1wuo7QJLNM2Nm0qjdFwOiJs9+401U
3nH7zANbmq9oGjgII9CBhcHz6MG4cOzyKaS2HDfTRNg6GcJcnm1/5xvVocCXGC5kxiLnhcJef+JW
XcRD4WIzR8qMMPSPpkhZH/UClDzKOjgj2VKA7rcQPklByiVfJYRLe84J8n0NE2psHf0/pBLHwzbb
pT4n+J2017ckEh7QF1RpFamZCPSfgeOlM6w8HMgZJpoQQwhTdAyAAx18+Y3akYVOUo6ciXLcA3HW
HqGV1r7xjvXIKjJ9Kc8bvscglVHV8CfAcIA2EuHwHY2Jc1pJ5dkC1QBAkhlmxDCE6oM6x2v4fOYh
lkKbPEgc5a5qPWs4i94Sye29BIIBUiQ8MJe+VN97k9RUpuZHQtOUdvCACahfLD0QPkwNae0e9WNX
7zdpwoFgFfS/TdW8Nw8MQo1klCwa3wOlOuSBtQT5Y/HRQt/szeGK1pEzF7fwo3KpRredzykLqpwa
WL1m9RJg6D+sydfpEvTzb6aHXCWmK+jw5G//Zef6heBvgLYGvhkKRZ3m7VPi+7GLfBJ3KeQFAMK3
y7GtBEi1ozF+1/VVgbnxmNTKJKl2s6C0ZssIs6LO5iiTxaAJSzCtWEsOG0xm/Uo+kE7ypN99g9KY
zg55UoD9Gb+DGYEzVo15nOccpD3TF+j3TdBUho12wuDbmSRPNLdXD7nOZ/BJl48Ck5Smv1WWHDnp
N7SZnz9Y5xDTJu3O5RD3XCw3tfiU9FFe/BLXtLq0474lCw6bxA9kAp1evwImXZg9SDHNB2/mIUsS
a1StwgwnoJOyKkNtG6Ab4Xp6bie4+x2Cj8vbsfpeHEyoniaIrSjfkiXwAV+4oE41HdmWs1JHwK0s
lWXKXaeLhMnSM1Du9YtuqTy3sgdmaUuRyX//SBHoKdHzzlKQSlhKHMMKaPG8UP8RgSL5srsuoUEX
XykWrk8Klz4hmSg+UBkiEbGLNmVT+57BkLfCYXQOGkU1tPkhEnynHXjwwoMxsOMBsANfSMuYTQIi
AW8z57oBr3eyr4AmVVc4ZY+/VtA7rxqaPztwGQLm2nABKPCZtMHdmp1VNxNijfHAL9TCcBPrUpcp
p9MkiEb8qNl80uXWjExKVzXHM56EHW9OaJ+i1UaCKmsCAFvdfyWSKpkwzGUaQH0kppLlt3FkcPxf
yfCakfzstytPrQZhtLVdLVOwz9nmzxbXjLLxDnXU5IKHtKWYjw+xZN+66/naBp6tLiV2arGOTvp7
+frEe7qeqqSkNvft3FlDDkmH3JtYWIR0J9ZLyIKCMrSiE6VpM7CGoESkfevVku7YP0hmOX8xDeKs
h6FEsLebmqYvVDGOmgOqZ1OLDFH5aC17j2FKVTm7dX/8Ut4YXOkyD0LORLVK5s9GWXyby6oWiZNL
iWpMMoo7xt/FWSQIaFCOSLA/ldrHmob602f4FswcHnVaHXq/q7gKLRKjUb7Ept4jdlSVPEUJytRK
XdhWZn4IApk+0Pk9TFbLjhKS0k1GzSZhxHxtce/pnmbv+4pbqTmySQ3BJpxq8HcpbEM/N3V16ovV
h2C1yHayeVoAI2gmwFM5Ubm/ibyu+vFVtg9v47O0fXvjuQ5cqLWfIiWdCu46PI1INuxKTcatj1c0
WY2TCgQzvn68JLOMc6v+XgBSTukAWMCf/dgIsw64pycPXZksAnwswkOiX2ZkzVN8tr9VPyb25t1L
MRzlqYAAt4cNYy2E4/KN8znYZ7qpRJZqYcTteAOZKRQCErDC6wn0MoJwBDkAv09aWOPqPim3fHAb
jsM1gtJt/cLe9BNwCpG4cVqL8ycVdMZAIF4PlwG07bR1DiDabC4i41WTxoeFJIv39G9L8kuwpx/+
asNEmwqXY3dXBve07KrTIwRkhDZonVIl6pjpcV3urTxoluIZ5onq8meab27DlCKV3wQwWNa0MA4n
T/hKud2JPK9abEZnlQb6K8f3Z9wS0ujOc2arpeg8pv3UfUgsUmpqX5SbM7pIFiev0f193kIF6P1x
BcyZ0+bf5HQVvEHRZvdHddEmjCAGPXBnJ0Nh/MWImAKF8cDtipoJt3HENV4Dbxlo9KmVWweE5tAy
3DVO2CpxR8uav8EMdQsOUle5sM0e4fHedoOjCtEMDC4IS6KxsS8y/wADdyUYTU9Ij8PPfLY+eHx/
ruge4pXZ679VeM8XoQ7GIGoTu53ruk2PjESy0SxK3DAhLZwlCNfPjA+yGyUdIg3z3MKET2y+RSph
H7ZfOgFP3DK0PB2PnM/6uMeUObpyCYulyFDgeeeIk3qzTHDk2AJl80ljiZCYnlX3iM0PRl1p9Rsg
dUl0tLH5nn57S6EaJg8MgGi9d1qdJok0U/k/1aDV23Y2oqqgQHnPQ8ol73jTWVRXvf25Li1YBKM2
r7OIOaQXg+x2J+QaqXTh/cFq8FZaAkVa+TfI6bXKZAbJBqVrjrqDoF+VBvsHKWbhM7/REMFtfzh7
9/5AeTEZ3k90T2eEQdJvzNxZJ6dhaK8rVvLDBMIfQZ/qRAs7QRw5zkxhmrDPnMjsL/7+6Rodsq+3
krA0U/6/k3tQdaCufwUhGakS8n2sg71FLh94iHEkB1k0Kc8UQv484NqSpliKMyweboGV5ElxtMlg
VvZFCWe5u9rdwUwR2k05UxFKtNQzEUILkp2CX083qsUwiF9C19BG/wJFVMBDw1ckwet/Mjrr5Zfp
fmM+C6Jv5GUFxEZUh2tU35nJ9ThzpnDFDwZnxV3bUB+mcGzuqlR71EwaCupfh+59fZE+62jAcP0i
jlmz5c/5MwGzW2bzT+xM4StXStTR4reQzqzcf2aekw8EIhwat7VG5vxwAE5II+TGtPNFNqWmDAgC
T3ew4MqOykPro3gJClVM4e3O+ghEEKpuVJgDYdYtqyGm3SHrEyGN/ELiPoFmTAohfmuxU3P/gXPY
oH+IgQllQdqq/hpd4s+myq9MiIYaqgaTFT+/nlDV9aoiTSrBPxTnhF21L4C6yVL/7KbRs2FkeSmR
FZku2WwNhOiQlolPSX8/T8hnaDcQ9TGLB9TOfqHkRl7bV/O6JOjYK+f/ouFjzRR0+kIxhJ22MHXp
MwbA37yt4ViC2FThHI/DDqLGQkUs2jKfKLdUOokYePqlXGKMSHU2PIY9rD7hF6s07IOh2daj/zUj
y8fCrcLi0n1l8BwZA59+r0EfFFtQ/Fqn0utzGfqfQUrdtSfjwemCXy50FoDFD53LhXRREpo9EgJ9
MlK2d5eSl6NAp/9nyJ6ip8nokdRJcRsDMgsYmcWyYVDm7AnzLWdBVzENAA7/W/m24lzT64SPAyDt
2IcB/uHaiUmCt/BQ2MJtFkv72Dfj5anNH3tbn/9vTWkxvn1hx16dv2k6BHQ8TEDOueBiVBz+PXTY
LagVHYJEFB5POJ8wVKcu3ZiIaDDQQh2Wk6neSjRtFvkXJINtvv90jfnVFJtPx00axcRv6tWIouwT
Fjl98wIUktiJNlUz3fAZ30vX/KBxrbMV77XTwKTo3IYAcxn1CQsVQrNOoMCzuEK/v6NrZAvgdfaS
5+XpiAu/MwEjtrD2QJfYFC2j20yaCBNyhbK4FrkmyQ1nlaJ+oWQhIkQx9uMcxeTyI2HDD1jAF+/X
/CEwUax/xzI7YqJlItuttTxwLkh7hZL+C5ZfCKUGgKHdCrtYUI31VsAgfKvyCgBj/VYU821WNWN+
neVtYsDqd2NoFfCizwXXI49x+UlkDPVP4LbNraOc7AQ7457IoXu3+3REr7OjcKCP3C55WJUHitUR
9ewMbw3hr0GDoe8cbB5d+P/tFa0ZnSyYbYlg7sORfCs1hnpr5aXtPHWZkl250ifZjyjfQFg8BpR2
V+RJwVSaUwfII0pp8bieY20JZ7XRFFZH2AGfz9lTbcgC81aSpSeHQMbDxpMNQTy7tK6xrMuAOIxb
8a0u5ffNL7pIAWA7l7vGtOJfPXiE1+AHAbTtXaZIHhDcFEyR6cVTaY1hw3LkoLrmiOWxmIrCEIWT
FbMINPlASi9wSTGaKUZQ47tNpHKU9PnNFDwcPGLsCj3rH1TzS5NdYUjrhUBtj+22D79WeK0UH2Qr
MJO9kDMYtVwkXWgXTsY8f/2DaFUPzh0WTkVe+mHoD+BaPlhdMRvQYCk93HDkuctljC1+CJhXtb2B
t9ywLTDJU1Nct6Ep0MiV+MC+sgBHKMgzPnjrWqKpsWQDzDCjgUmrWQ3nxe6qkU9Sb4b7UTNNBy9y
eoiiJn9tbdQA1BCHbFW4F8OX4QtatDJrj7u/fMQEkEY9n0RwyZZFHW1vbWazB/G2opQYbZV0S/mV
xDLGH0EXn1nWbvB2jH3And3Jkiv9V3KcHSSOL+xNHQZR/g2u0GOx4dgv7hQ5PcpUFY+D9gcd4EXe
2baKq2yzy5AMz2Iou2qRXhApc1krpfbiIqF22GbtcO7uG9ZBD82tJ+cun1e3i5s8D3cTh0Km2SEf
a9Nxg0HIYAeTwJk4F4afhw2NqTsv7Qgx03NXS7MrijPf8JtNt9O7tZQPG/z3vcTupbHn+KIIwthL
Plm/wXdijB3yMVpPpymrdt1nL3WNbVv1QqQJNS9xq4t2wBv0oWKl2fVLEerXo0gqBQYC9q9GppaS
FdHnfT5YEHs3y51eDJ+XWXroxCWoeENa6TichhiOgyRdZbjtkpK+DS2hGsMCrHNO1Q+etu7x/ESD
frxm6oXlMmd4LxTRltpzarGIE2WDIFS1DM+cLNvMtm2G3l6Fa2eIEUNrjvDZhyFOZXBR1bvk7mlU
8me4kWgSl9EvmIOGND4LPRSawNuLYK4QSkcNxqkjXjf4uL8nNQaHTCI85GPzWdMJKkiAhZqTEEwZ
OBZ56y+nMc1slENf7Z/8oz0IGt+mkBtNhzq/dnluHKpa10ckZpvd3rLUNBBhQzYHT7ppGCPOQkxh
rf5a6CRtRbevvrKvxlq7vepgFhcits/syVhnnVQ4unlvDG4rUWQHZPrIv5RX1SxoFMLRwDZzNmWu
Aou68zDmeqU4V8y3fz7I2A2kY0iTsK7bcymZ1zMWOCNtS5i+/X1w2uWksHeBssxk+BCqskF3fC8Y
30RhAt7opnN8ikRLw4g0vhCC7W9WPNzIPlz24Jdp9+ygfR2GiSPeOHVTlJdf5/zmflrEKQVzX0+M
2HDXFqVY6rZJ5NqLe1pRYpPpweT3WcX45wwAWYQhY9u85gJLgxH52HVlYqGlkSOZD+/pasG5lzSg
dupiMY2zaS89f59M6HkDZTUPhTgOO1GR5QcAjsNKi7j4M4k7klwBjZ6AfkOfgZlxgywaemf49KaC
m2BrqT8huuVQIKtqTcp8HtotKo8f4xkTSKdRYpE9a9wKQDutaS6aB/cVyNSXUA4g4S1S+ABkrFqX
gfiel8WIXOLCMjRayZ9ulErzQeJiN0T3XVtliJAl30kBzzTQwJ5n2LS2m1FICf8A3xokEoaTaiJu
iU0nhvBw73ERgQ6tS3RquzmRDo7Hs53ObyqXdZIeQfK25xmI89pdvmA0Ha8LALov7ADu9+jNTJXT
PVu1hsPQ91fgEe8qyeBceAZrDSh2i+x5nh55wxZUTeeDDy5xI8KbHI5XgAF3HyozrvDg7ruJ+quW
/Z71m6aZPpu2mMFFQHuxxorb+nB8yYbfVMtE1alcHgOZs9DYdMCsTNHLlgqrqU4GXfu9a8qu/eWu
2mJTbfZyXpzIfjaplpxmggPebWvEqjGSDnfub5YjqSUtv5s1n+afvKeoOOmMYXLZF+2tkVmXrBgP
7K1S2rKMTYyHaXstE2TYC9zM3fOUiwlQHYShZVDREJ5faaOER66AmhFYr73NhXP2E6Ogvcu1NbI0
zwxytoDCR1+7zSZg5oNgh+vlwNp0pzSofg/HF8Y7MjcyxGmq3MOcNO6tRBgAjYx+FdnOwY+HZMaX
p6zMXKBGaMUkPSgGDk729dKKv73c3AE8Wi19g0V8cKKGyxaADr15QNCYDL93XRwB3W3tkB8Ou3dd
TL3jmETI2G9MKGrxCBEmsjMyESPOr2wdVDDLgp3rxiQJ0YlAW/cC6ayHmy/tj8PqIRdH81u1Cxc6
hb8QAhKIxsFstlDkZ9maIAbVRS+5gyEy2ZARr0qHFp/EoaFEvUwktmGk6mXBBcVa039S0Ee/vGh/
ZuE40I7GO9eFkoAyug5+Th4nyq5ZdrcTaeLgIXSIiuriGo1AN18lSFzKvXq30+S951lhfWQngnAP
kIMczkkhjimE+cwwdOdBwe66F/4zUQzqtvprgAP6fhWymZFJ8hHQn5iUx6X1FAbkiEd2HLzA0OcJ
Mg+CaOVbtN7yg6Ud0u62BDZXfn0jjrk4ID505srMpU3FYOh0eMIXZFu3lJgKsLNqrq0C9bCf3er6
kNE9t00x9R+lVMt1Agm+sKG8VabzSu6lTqUeV2uFB88LU6nRomj4+Asi1H/mCL+Wy8dAwWtqMAqV
9X/nz7au5b1pAXWm+hLsDgwanxJlgt0I03qQXjP4swC5eyfYQ9tKUA0C6DxPznN0zKHevicCdPv0
ruQ4G5KM8bmAP+dyl33CuNoSN6eWh0GItZ0jHynl6rIt5zPpJy+FenJbOtime3PU2XW+6hl8nJcZ
wE0k2pPqWSnM6TBUveSaiU0wtDiVYI5QrdLi4/dkP2/vMjDPx9YY6UyQW+u5IBctjAuG+bZPJiJ/
XU0ubZzHyPiF0OuKGDc7Jm29Vt2E5cAJbzg02kRjdgQV0+LalnBQfq0HwX86Pe70kYWI+psscO3T
8YZEhcz31vOehEheTp5yn7QNTNfzzBOvH0XkyrrzcZ86kBz6F16EyG/xlIegiFA/ejHrUZf19xrM
t4lMNN13VEcFCEkV+nKZrdEWzMp7HL3V/wVIUeF0+seLQ7DSnGdc85JGHt0SaMrTtWev3XzCPZE9
HYKUDX3x5gO91lW+qg10y90x2exoRD2m4n2rjCZ3GvT7N9tJ5AO3CQfznJyx/kJB7hPPa58o2vmL
DnDsVYB+siLmNrrgZYtpp18pvDqX7WWHteX24wZnM55enV/BT37wNDGqx4dKtVMzLVg6NeX62NzH
szF8W34i24O1TnzzqaZqBb8dRze3dvj1Yrk8fOgz5OEpSKZBSavDc/jL9JaBEgTGmcRGe3wJWMLW
yUGHQisNzs3BM4wKc+9xPw5sJJMdo0XIkw9JyEX6+nV1X2f5JFvedhAp6qfSl4azEYkqJE9FhkTO
eqxA8+F43ixmVRhjXedtg0qKQ00uJ7r8DpN5ZvpN5dDB5lXWHwS9aMFZiKBYB+W0qalKTQleE9Oj
U9bNBBM5/U0XekGaHWm69AWPruWV5zy5cpsAcw1GFH/7Waz8M3feJVpKV/0l+WAh1zppnjEtLWqm
rKlqwnXpj2UOBcVg6hMHknXnqrE+LFNSWoIN1NUO7OZw+QMr4ZEXVeQ4r7dRm9RM/JK/Lx+JOpGk
Y2yzUivDFtESMTeQugz/aZWXOqegFDO4/l+xah0XW8eYhGfk5hJyhbxMbkAbxrnF4jxiDOFMzUgt
IqbQyawuOxS1Twn0M8y9b0xsdida6EoOE9ZD30GMqTGKJsl+Y0HRiMK2/LNMzSxV6NWOr/ROXGgm
SzVtEh1bPrQSDSGOL3fTi80B1h2N3GHvAhx497zGQxotyZUgSvjbperjxTCqEDe50066EOZFiNcx
O2xwLEqMuvOLktLwueN+fpgkHeSc0lLAK3TvwTpsys+M1PfV4XU96lU6Oj3GrM8zvCtbu1vIWzug
rXXWNSFtfP+3onuOfFJVhQYX8JJVyxHEErP9iZXZFeib+LzT+mUSPZLzZ6jVel9xITnXb8AoEPIn
qff9ZohDguXf3XxP+7AxkaCwdg7FzmDcDuhaZgs8YTHjzW6uyt03mu9kAH1QLPSnWAOw8W3DDU5z
uznJkciPyWfpXZyY7uXNZpUu14TD0rQcaCycLMmgR4d9nMCI7K4QnsdELDeyxueFdVyfFd6DSviK
nPNOrOisLZVfh3Wdmj2lWmrkDn5YOAZLY6ha8gFrlgFjKgEZ8MO2uzp/SSQ8BjPVKyJ4Dx5YbZiR
zjlpPu1akbBUmXNlw13wqB1f1VjjYrJ/bn0xGaWuAgrzRaRqK8PtQiaTpbhuy3kRtbCnkZZ8CQ4Y
rVDhOwAC+SMjEcGI1vLgXvmsHYEfC3uVGv6fwYfrSASYOclieSgy+jnR3LOggILgEGD944Hf38oq
sItTVSXZ2P49p8/s05nVtrpm7ofptaI2jsTXxEtUEKBLD0Dzf+1APW7woJVtha7roBlJ4Xh93EzF
Vb5uRVY7COaWq/3tWT9fcSg8fYPw6WPoZ+yqU4apG6PXyl0EJWvXk9zVkkrlMEpWPIEwdYcS9L8n
j4n3SoEM7kzBh01QliNzbV5NBE09khqSDywshsMRnIIEBb0Y4tbKYnhdtWelHp5c9xdnC+0fCW3p
MmX6tJqWPOUnOXFx2WlIkYPQPPEq63DNiONWXVuzj3PFCND/oN8qPaUYlvU3SgX1JK/dNGCbEpEn
leSs4n67JqUaJJrFYjei9efKxrSEcMqyH0OaaTTqqLhIxO3TmdeDPOIqWBKzvDtjtvYCNNJJ+a22
rHuyiIXpfwZv5xmBdoema9MZRJ2E36KtHTbVnMOQ3Eb0TSvnSSzHyznQZK0/MPJxEMRSeK27qYmd
KFs9NVGRg3xF4AfR5hRkVomY4gjOAku0uN7ZRi0EClFkQKSeGz4CZRqTWB6kz4/i7pJ4HFRrwcTT
I0Dt9rekzYfSq3+u8m/Z/ScnEsaa1wUklzkhkyDZuTPZwjGSVtfATt7bdfWfRu9I8TUIvjLyUVFz
YE5lcB06orqCpYev94o/O/T21Gp3v/u4sX64C31I6WOzblz8FLEDVgpRefVSZs40UcCGxiWQA7FJ
5zww7AL5VaY4HOGDdzZha2J030PWuLPPl9PdlbeuYr4SIApkWndUsFQ7xVo1eo0WjLFD2dgFrUBY
3ozso+H3kRb7xRFdM9WgE1gDGC6DtMY50LdfTyPl/froA72x+06EM/hJswhYp6X8dQHsnLEmQTcF
USokh9wNuc7WoDMU+A132Yf7hASaUi5OC1jGArR/UTY8U6Nfhw6L8QBf7rc37rDz/5wQcGWzs6yh
mPkpyBDRCvCJ9Ep9ADzD/w3BEyHQ+0aY+ksrg9CpvQ3Iok8UDfQ68YBuxQn4dJVXwedGWn/YOu0K
1vjxzwyLYmVbtjQi43Q/GSqogqARzq5+7L1MNcFgeo3ddz5Aw7N9+NegwMA1vXgGS/cg76YDU6pZ
5cjOTe6hWbcGuv333GlnnUS1R2ZvmlLDS2+RwJLwATEnkFPN/5gBMfnU5yzONqI3Y/28eC93YESx
guWNb8ytwZxDMo2qDYkvbOfmDAlPYD5uZoZIbX7Yu7TudfhHKReKQHTXEm6m8J/TO7n/goQ6nSkp
9+Mxnfl48D8sw1btrz9DGLYlCm5JhJX3mr9aLz5llLhy0n+R+TDG4QGu4sLKbCRk5pyuL0oIu1DR
TAEWa7xiSRwqj9tdU0MFBNnSjVd1VY4wPxy2nDB3EZfIOn2rifvYEiwmu1jalUB8mvyzfAuXwEpr
nDuq3wMPUCPwsEnRbV2Gtb72SoeRQY5ywSBVn9qTV+YfC2Kx7KDjtvW7/X5rt14BKs8ruwM3SWo2
9ZPeYYMTiEmh8jP36+cbxEJJb6owFsiu7tzl+xBepSnOis/Qwedcc6UF8oUuoqWRnCC0mg44eote
66pi1qFDwba274HT8VDwFC7CxAQC2mFeipP9Wux6Zk+KG0TlXjovEXWJWSnMAOrkxmFxT2WwJFU2
bVg1L5v+H5hREW3DQRJMvNLW6Gz4mUvBa6msxhrxLedI24o9Axp5Cknjoe3encYR0bMNpdw6FHew
zYWXp5Ch8QOoT9gJDzgxV263GtvwVRZHnk33bD7d/SeicdhFteaXF3VFg55kXmnIeVOnymrLVJAL
7G3ShL8e8VZyFjrmQmeWIGWQzsbYxjdREhmr1l359QPx4OQdiES9pNc8SpG1QnAgaM08OfBYneJu
+M386B/sSUg/RdngHxa+GUT28fDt982MWOvw/UECptHDwboIFb2e1TFC/JiBvCaAmpdNPWpLT79q
dTt0d14HaTy3YJYPlkQ+lK5/dWsBr7Hvb6gjmFKveN7x5qWfN3afFdEWMgxB83lG0qxkqMwUjxxM
QqlQeksemarbHQ0v4ilsg+NHbPt4yxwvGSQS4f9DVfS5+0RgRLacfc6wgXeI3qiOPHKT+O9oZmdF
VXbln3VKRayL7z1dAKO/LEuPPbPgAkXK04VWWHIvQC8xPag6H2YBm/BJWl2lheLJzWhtHXycJWsP
JDSuLO8+tkr+M+ZchOb3GkKjInjt/uKpekE3khq9wZVGh8wT5PGMDLKwodTC4QIaOR4yvGst9Jqz
NL9QmAfZp3k2ZJCXeEW0gWyRLLs9ghE0jU7N2J7m8JCI2mvLaEKoqxCMPZS2j4rrcS1qNznFVHTn
g+jJbw91KMAMNdpwhDaLCRqOXqUp8eOvpqIRuCzCndjdwIeIUqyQTxqDCdMVeHoMnxsl0V0aprjw
G1dZayI0qwAEaQgfmo4ZZijoFUdyia1Dkmsi3Q4AKYVlBr58ok5nmpj8d97pNIsaPnvdL6VaFv8r
CfyyF5C46imMfn6hJDV5cPQyPosCI6m5JjC0XQ7Dk5TYQZA2qoDZLcOowuKm5kWyoJQ0VlpZW7hB
408MsUWMdJ4hRY+uem7QvMZvmc2mYjo6zlaQfbdI8tk2T23I++taPJp4YqrcV9tv7mYXIjJAwy+d
rrKZhBH59C4oAfI8YESOCzkHUxYW7aL5Z7puIyhOBtTFIt/NT9TaV+GsmY9hiWO0epNnNu7SzZIk
VgvixZuIdtk+Qjc/8A+SRmRC8S/6Z3TQlhbfsNi9YFgpyiK/M4XthyrYiZa9R4rT5KNE0wOwgZeL
FzJ51gZc8vM5L05o3fdtvuZinvH+1OZifC5jJHwVc1I2WLBj8umzhXqvK7e0n0BJQqSFsY5DrOQP
RhaLPKbEZFb2/JYU8CQwbXvt4XHenYx6KHdZGPdD7Y9AAqZQYnIkvARmlfz+fdSn1MPbAkjRbnyO
UMyz9hhhw6c0Uegji4wXIxq1uns6JMW7tLMmz99kqP8K79sL7o0H2+4gHQ5pJG1SnOmuXPcMGhv6
QGYKpTDoPdeDPOnDv3leILmexe/L4ee879NteFnwbVdOVcmuCXtReeDkZzZa7UxErmsl12TGJzz/
8EYbPqh/d6YHpMvJZlyRkoaKjTYOff8zWJnuVIDcz+hc44nWISKL9DgtWQEQtuU4rEVjrYis9MzP
RAp/v3WKdLo8f3WXNUJuse5yo6eRrWXHep94I6QMayaaB8cPtAYl/fnwFhOeu/aGUZZFTxlvKELa
2wSKaceZPIaLsq/cyJV42eLnNrGCVL924O9mAKMgvkCLsXLaEXt2sMKRFASs527bwh/IwB4MTbKz
ZLVzqNfftdaZmQydxqARdpXem5lRuRaqnzVBhWkcpLm75/+E5KjobFLlo9P59pdATypxhQHV9mMu
18rMUPb1+1BI6663LLvYLlhRMz4Cg8kDMURziv4YAZxLauzdnNnNt7AyOUabI+vyX3iEFg63/SrE
zVgeBdGsseaElJrTzv75mdSMHBoiJY8MxknH4/OTNuEfKdU8Jk8PSuFm5neivUFwu5ZSouadxeA+
jjHh7zcU52Kr/LSVuLRY3jSQ0PL2cju5NdFlEDq4A3Stex7FquijoC442JIML0p5h09vNHV18E3l
P8+RCukv4EC9BYtLV5FGLm61ulDbZOtmBKxBKEHXlvSkh2aMFZVaBXcdVupSOFM8ymrCsbvJqe4N
KQdScWplX052iMkosIHpA2smyZ091EDx3tI01fVv3LkzUiY5c51/+I6SacYZdy3byo+Yb9bK2Vne
BcZjtpub48BduINUUVG4p73NhUiLD2ehza8tIGj3gzmnIppFoiLN8BItSwq0uvisJo6nSNdMI9o0
1xHjXwMLv/eh5LuOmRHrKtVVuQWa8pMBuIEvlqnjCgWhUdfpKXF9wffDb36VLxKiFOoCAeBGQzY7
7VqM40MLk6SYhSQapOfhpR/svZab++es0xRhigVuEUip45Ne0uBJrLNtsSiojYl1HeHMAXmA4BRX
nqdcr3PhW3dA41pIgPE6mQYtXNSZSQLsabmVxPm1LYN0E34D3AFKk2ITBbfkfRY+vxJvGidy/S/z
MJGibGIEijRZSiH3KkQfVzEB9VudIemFedqQX6HRXxV26cbFjHgvQXUYPRUhSv8/L7od58EVoBtw
zbW9L2opsT9rYsDpQTU4X2uv2tMm2oLRm5SwMTAhY+wC77oEx7fhNeV5jrvIB9l/1NRkMvD6fUeB
uLgpPzp3GhbNFHnabsonRiET8yRV01td6PiYlCIGGf6C3QHdarcquYYJ2jeaNCj6+I/k3WoRLWqr
R1mRPCoUfRJKyUIwokP4nMzIuEIW5Nomk4lN10s6EBi9+hK+3OsvaMJZ6k06awXAvlHodvx1VDoD
S8TgFW4RhAX8NzD7B8sfKuBMnbaSfblEsKcewj/pKLnKH5UsbAiwSLQ0HoR+2XIUNyKWiXm4m6Z5
PZsNv91dB34ik9DTAxEI1PStirDOlD7LQb7O/k5lubSIF1ojAp2xJwAjDE9XiFpGv5Ya17EhDamR
4iXU6DDdGATb4V+wMeouxntdug1bJOSiM9fhXGI02ASIwdlEE8SjA0JUCAtExi+KE46sl1M4793L
I87U69y+Q3D9O8EpNOs/6jsrT1uflfF2aj1PDRKxwG6g/CM+A1LXCxHpvNJvqFZ5LtShF/RXRr6q
fasRToOo3hlT1PjHJQemSUuJ6QhAPxiXOrqg+PU/bx8FNeTwEl97xBZGmTK+QmcbDB86ESAoC6CX
If5E9DAjWjM9nCfhrsvERJb9HQ5mtAr3reiKXqJSCos3Cjqhh3N0jhT+tzGPA9koNwIxNzhrpiov
zCFLW9Am39O3Xl1XjBnqmREd6RVR7m3WdYFmSp6t9KOrBfTA2BljQEvXUkYeUsEQ2B35az+rsPOK
YVfMCTN9qpZVVpua6WdEwHaJ9jS/Pk2qik9oWGAxJjPojHvPWgiB7bBdEsheocfZmTS+PsKwOTBW
sIDuvdFVw6sgKojtUgU8g2KCpA3RVDyQTG95sXiiVA/dY79TGr4Ant4fdqVEaT5lwBWz2MDFH1ry
sZAmD1LN/IJhzi5wx9dwWIQw+Xb4JBVgtEKvVoJMdo8s2dopEIDHe7+O24hMgLLchJC9ezgNwZA/
aX+cU5btRx0H8h08Ix/u8de1wZpsp9qza7RygtnqsQy15NADQChSHWIQlhBho9nuuo76lcyAIQ8r
vuErfo4rcHDoyQiirctq/LM9sVBeLLaM1vVz4acxJmnJz/jMfEnLnTdkkKypF/9XVuLB2oeDzBoT
NFLQhydnSB47j8Cs7T2jMAAn1s08vklELvUneIvPO5js6x72BJcOT7rJ/3T8lT5UEGLrSjWJBnkU
PB9BK5us+5hb8BZuwdzcZljQm/aGToASFuM/KiA4kuGgEgDzgKMdMom9OHPOgIAD55n64jR9m9Bm
tel20Ju07KhKdtos36Bgimo4FJAtFyiri1xpwGBvHHDTHNa1AQZv+OU1BOFxNCevWqd+rLo7Lrwl
MFHNZd4BvCv0u/jdbFLpGT+8sLPvF+smN3NRgm6bFYTeoMFaCDN5KxULq7jSmeaaQc+SBgxCyQAM
ZWUmnIW9qe9JKnkV130mQgR0g0xyRHlXzdL5txv9ghkD/jZpn9oayj7Ix5+IOU5b1WfgKRoIwXC5
ZTtjCy8UUz28cd9z/w8wanL3oiS6T4lwdQqHDrq2A1/0fU6IrpC3ZRO4OjGqIJSTqlLSbTT/7Hv+
dCbYe7gCH6BzijEl5Tfq4T5+G/BlSXdRoH/GDxyoEwlykqy4kVmddQfpn1BQxjk8CawcoAPweTUG
OxoqRsanRwAxzJwTG6vMgG+gvCAVZEffzFDVr0xX6BQvY4OQLVgqn7KB8o4lw0AE57qzPLKyJa4+
CFSWtMXsV+RvLQf451EW9nWvCuGXoWvZ7GSvbE7xOiV6eQfGtjxW/xryqw9OfdhkMW9zxpJdqfMx
cq7OETG+yAdQ2MFiTGssdDTvhNyR4+DF4RyFwN2L+sl2xt3RiihI7rz84BIFaihGdUTzI6/kjn3i
COoET3ddBcm5rUV/XryS4398Yr/uSdiU6Ot60raQHnke+3XKz402Jkp05fJBGeS0tt31l1YvK01P
ws7HWOyOqddsl+IgVGTAXTvHtr/nS7HAoDpEswsqSs+LOXKCE5dalE2IXv9lpdVxyY5RaTjH2twF
7pTbLKoc2h6D2FoNEEk0/Lyxuz6K567ESLziSH0XfTwjWPrC3VOmX6utyg4wkbC0F6z65c6h/VQQ
Vv7uatOUsEqXh6L968ahfeqjSl/R1Yr2Tzlz1lGCeOHE59hNGdh33WwFqxtE6+726MQFRFaY07cU
xvyyNXTvmYJh3KWgoqJYJfl5Y95aR80nMvJD7CBtH9+voMoN9RfVEg0MDtHPLeCQiVV9xbg5WnsX
sHVSpLFvWUnxcUUjs9GErMw6NGY6l//RFaQYJzSXL8q5TRCtFBJOzUQgvG8EIK5UI4B152Z/KJyt
1Ys+MDGcA0IpsSC+X5LJYtt/mAQq3jaBoI+1qPeDTULV7DLhPm3V6zVdjDIQ+nYUsxOzq+aDBqh/
QpC72LMU9dARSbLJ4ma9d+PAb3ifz1KfRs34JprLxYrFn45EWoLN0/UHZkJEXh7bXfpGmhvamOvL
+2eR5GtFfTJloRBFvnzmpIzm4KaPIfcWLcnJyHWPd8SqukYGgF95NV3toBS7r7dhOIMjfphtgkRO
ZpoSv58F4dG5WbrK1DQ5aooRzesZg5+Qy/UfOQQ11b2ieE+RlijzRLDGCGTcj1GABZ9WTQ6fLZJ0
vcwre2Z28Ltec1OdAwCUJYKFqZELQ42UbSXa+Pap7jEwzGU+fMOsm2HvzzKUpVin85oQLu1t41F+
esotGuPk7i70H0mVb6mKRIkLLkHNMf8JWRh7wefhft9U22DTRB/c08jWu174jGLe16Qp+uCwooic
z61qPMcm9W2usuK0+M7HE/regmxMUCWIZRncjcyFDcvXdf6FJ7n4IeEPDONBLXkngYPuaxAdt7lq
lTlTy31qeFzywdcnFomKxHnTpxJK5IRmxbyJeYyuSezONZjr1Hta5aKaeIXpSwvA2A6dWvz536Hl
IfeMNCRN/K3tiJbbZtG5z6FfDyExTXrT1RBlEeXuCP7Li1Igx2/OBDet9/w3gb2lMBUJQ7QDiDUk
X9hypbQWNP4Q9DWKJxNQioTcTwq+3loEzdZ/sXWADNUznF6wR5Ut7t7Jth9EbkhpshcDpMl/xl+R
kcY3xAjCajS3wSSvJLkveQu+HRt4Bm20WpmJqWmKg/6Or441/NWKePUHM9A39aaD0rR0GYuFNaON
j4+2+kKvo42VqF9YLsPrNpK2l0TSc06kyZVg03BuNk3TDbrvqO8geoH38XjApsnszyP5Tvfwjqef
U8KlNTXWUHJ33wgtk/DJxgbRZipynxPOMp+dS43c0PHeaPSINRVvA/uDb/w5tKJquVUDkWMV2Ktl
yHqubLekrJDKZ50MPmAlzt018XevlY5kF9sOgWsu72LT8JMFGXDASdvErDpWp+Pi30VyqmrFDrRZ
rVf4yh1NqtIKuzHD1m06O8Qch2u3PFl8RJOGsM65tMJQXrqg1LBi4jmcSJEhmX3x0jmLtb39uQOe
neGQGh9zdeBPwGCdtLYJxIiY66yTf803S/lzlYzo+RfAiRUlNV8/5MMtChZ9E4nclknamoXkySIF
NG4n1hgPQFxlbJYlhem1GbNkbzOO8TIFH2wm0khemAMEpz4zL8Z7Q+Ix4vtPyrUfx6KkkDTcnUTZ
/2aj3WFLx/0QL45WmBRQMX+PreQ1awH7sRUtsFZ0rGBqzybRYp0H1aX+s+Y8nakqT/tqn4t3NlzU
0K6JruEf8G5TFaZsVXlr3ie4iDgS0QubUokSksfygB9O6GiRW1WjJpBcJil3xFubvvALj8bHsiPc
7xeax7cK1FuDvx1jtkud1X7vvlcl/HHUT6XLRikGyXslZ+Pcm0WucDBH6hZnQCxCJBFpVEqDePdF
OhALe/Vy7NhOmcLb4mFIw8IuDt1xa9sMIbh/Qk9b1cvrATbcpGgIPOkqrrXHYptVEps2b23d1gm+
qCA82nVcUpGqspBOKBLPPFew8jolyf/AhReCYgcQmTLGuhP7X8MXvIhwhZMW3x9dthMxoQgeyYKF
knAsHE3b6JkJb549Rh4fzGNbalBC+yNaLjmUbcWSfc6749x+L0VgggS8sjK8pLe7uomQyG3t3deq
Y651iYEHDdUFnvqCRnaMWwi156VI7t1JsidhyxdrM/9x7PQsCKa3bj9JUr6C5pfznOrQY49xU6+X
PK0MhyCLikPmo90L3INUYkiEf3Tc0xJTsPt87YOaBaTqCo92oouQQjVSZjmMqBut1ovLI/HDauKr
fMDPUXSPoC8Kkvt3ht1dwZ9wszmvFkiLy3Ix+4F8zp+8zvlr/3rplU78Tv7Bj3dDaC3Q7w1KAZS1
yicemyHGYczyatLRl/R/7h84oMDuIIG5+OVx99sIHZmEYgyxRb0zlQRS7Nku9XmLa4NO3O28FqjW
ad6iHIsT+XMF4/NNAJgKdhiZJHEed3i9kxs9y8MzQ8M/Kx9zeMeOjxPEr/xQjBBy82wWSub/CvcR
ck8hbY9P6m0Z2f5vf80fMYOenW95GjpHG7nQ/xdottiLds3WWObC1lvvCQIAmOhFyy7qCXW7zjt8
KctZsRUoUVq+DGvElC4GyezoTZ4R5w74EXJxZ/CvE4otJDDC3eKtNVR6dU8obGeSI6sKK0aQjDmC
ThgPNQROmxhSCzFocWrvuJ76SH41/9JvuHsF3YV4wZcjcwuYYGOAey8AwRBFC7TY+qN17xfKhXmh
YbYi0je+01jp4hKWlHj5CXC63zpX6/aH1CF/Z4fzdq5W7Z9KQV/q2ivPQd43cv5dS2ri4JX6L8mH
H8/ouPPnqoDLEY8cpsC+1R5fhB1ZGGZvi+dEh0xM0k9TjUwVqznCcb3DC++yaiuhwPNRjEI7i5TD
jOZYrqmGSebE0gaeWzA5ArM6oK4D2YgppI7YBOUZT7aVFhE+8onM/+3q3IG3KM0W977kWjf4Azd3
3LhhK9lbs7mLDF8eA5anJlX22P/SOh4tuebzhmBA/2/WHkyRFbF/4eAVw35paQHAVGwO/i8/8lqg
/sPV4t2HAefp3Qf5ZN4XI3h+yp6+gIVHRcvYt7jzJE173Nxd6e6BbMbO++cKQEDTxu3hNzo2wYzD
fhX0wiNJalnZPB0bb1zxdZFNuNz4OfME9e71f9gy3hsy/oZgaRLKk0LnOHoMfC22LdcNtX8xKYCm
DoXqJ0zjwVznCPAzBeZ6oMpFtXJn4qJVUSgyi3Y7HDrNl7WkJ41weEANB/FesEETPxiZAUqnQej0
4a3P7iRGQavrkrepJOu0ui/AUHux+cM7hVIZes84BXT6LLtEH+ra2aXtilFFcSMP2VJZl3bVdwtE
TrI+zuSe+HTJmRWjSf/iQPioFwkagRnxUIJV0426pdquE+IHIHACXWPlybqjDajekjtzIjOaQTCb
pXDmnEen5h5t1h0dOKBwenhbVcgYmvO34jkDjN74jB84vzDx+yi3Z6ZOZT3+rc5cCqPdH2hs5ixB
LFSJ8C48BNVHI0pYGYqoKmStjPI9qfjUoQ+k0+hHAB7E+tfps17uSKLuAGSgJHDYPMb2xyTVYAA8
TB3QgpTqkoIAghVfWI5f702p8qomejObpzVgma225DJn8gAD6IIDo5oPHFG3COU9SHGGjXSbSAbD
glany0lrCwSFGSddyZuZXcIMFxxYE0gqZvqYUPTQjN2kBhUbmiPNYPwdgNpYcs+5C8zPFTilulpO
1CBCfRuu0uQryvsywe2Z2Pc3PiNLGL7c4GCi3ZdvNmV/iWXbj7QcM4UsoTqWWs0T8DTbId1vP2IK
4kLE2y095z39Zxbi33PefKmXV6pHwLt9+U2xiIuckzBS4O0FjnNpzCIaiIwkfWeAnK25haFcBOBV
IFXCaHEV1YtK99vCYUiwTyb/Xs62rue+yBdc3gIvcHVNgbUKOZAm3oXnHygWmq3++VDctSmrHB+J
K6ixFGtjePFUd39O3ushJKicA6f2GeLmKyBE32suUAJgJJSEoUy6AvCeDNooan67MhXgjLbPJMo4
dbFvV4K6/xM2nQ/5woRySVh7IBT3n3ePIXfS+R1Ne1SNcbe5cQ8BIheijGJd1BIlaslFAi8hDYsM
rM0eXGcYyzxB8MQMfHyABWcdbTw4/904AQN0eHzGXH79iriNr7wV/YeXyCDA6lawu8EiqElbB9DH
5F5YfqoGJR36KkauNXIpykdrtCDRUdYWoXUC3kdCph5O0B6pqI25hPNDfY6kY6n+Oxi47oyaUbWx
ulTx+yMRtCh1710M8E366boBniqz6Y12dRIWwXWbgGLfE/PWnKjb+qDdgoFv4crPxQcKKk4IgSVE
nS6wjb42XG1SUa/i6tpHfd6z0chXicBQD/En9QNk/nHTeTHDM8C7y6GTX3MB97l3TNDWCk/gM96Q
sPmmsGJOTI+tCw67wavb0pcRwupwK0hfyOnbyWuDxWkK82rinlXVVV6/qvSRkTlMtZSF302uLRpg
7J+YO6zO7L1ukty9jwcCSuG61v0ONKvt9WYVA4Gi4CH58YCY7QkhvZd/3C4C/sBG17U0SNUMK6Gu
WpFl345EKlQxI8160hgC7gJ7KVVuQtLC7e25v7973/NDknik3iVsAEOXBDlecGCSKrqUM/XAOeYG
xVUKvnf+AoWQ/nOh831u1gDGhrnwEA3bImRD0KOomv5D2OnZngANqS9YZTF/doGibbYBnZmM85GJ
83uZLTtQkjhhlZMAqMwedBROiz0+XAMUukeVLKpXkRlQhHWKfSHeCVrkjZgS6QhpPZwqg7CwGEn4
5CPOqB7tUFo2nDt/JOHEHrA6S75FbRdjbQEP+gl3TI3KpwuGw+ulPFkpB3TPbfplyXnORDSFvtvw
kSDqo6l7rq8bavCyJnZ0VM4JihHY9CYI2nSJ2Dg8vuUDlei9IkhexdPDcmDlDBjnIMqU1XJGVsyr
kA+WucPGGdZaFYCuwkKDgnLAuELyTa3HUV/YlFWBBJmqzu8MJ/IKuxFFMfNRwk/k9eTm/iQ6LCAk
ICeSFLvrMMyjqzLMqH1HhxtuWFj0Ynu/KLYfwidxXqrvmSZtHPVkeOFYuUyOIWWwnGj3OakdptZZ
eURrp7nhdyVNe/RxSjVzh/otJn5YbMN6eVn2X7wAxw8kWuGRICdBJPb+dSp5A3H5INx0DsSTrD2l
EsR3B0Vx6nIs3nLYV6aj38ablXl0+dfEwvR1jZUSQL6NXHhswBgMoMln7/eNZSILjh/Qbdfzeai9
tZRJ5f2Y2G3syzcCQObdkUkg6q/w3olJrOKg7iLybxNVex9PX6exigSVwh9gWqNDNHiZx6tqsWJC
3P44IHN2ZSBm/DkVN6pkC6/UZ2arkMBHzKVGzJRDU9Y5u+diTUjmsUxn3iyVUpaNQ0zFW9o6K/B4
G19OXefDsL/6lN8wtqFQoxmHjXfaqcRQwTB+xoCqXw8/bOqH8/XAmBoiYSIznkp1xrd/aBoiSQV7
1W/i6yaJLrwi5wRVlRZX8jpjE/1MJTpD/VAzJ4nk+aciVpTXeklkLQmfyYtrO/Mr2j9fpzg2P8H4
E0frZdCtmrHYy5WoDZR3JPdguIN7IGswSfLCS1TBoXyWSHxFJfrDhd67YMEx7fz7WFeazqKGainb
PR16NX7eoOkTBPgwofRLUU911HHn0EkpcA4UHHhuMBRIarrrdrvP88BM7AVIFEbqKEVOuKs6cTMv
Al7ZKLwyWltGiENNNMumOY0adIgIWXnDj5t174EzpKnNJxMp3UetIWLHE5k+Xxhkrw/blfrQ6PS6
YHs/5YtMKsn74rCfOLPY7um9SK4vPiH+Zx1dcST+jwXgoY4f1fUDOP1MrVbTZq8K3X1qX7bPE1R0
G2cSo0gu/GFEl62sI+o2aWItjYvDYfEiukCzMrLijecvTncis3T8ivst0BWk2QhTjT8/+OwV5I7b
bHauYBFuAX1CBFppM+uF1bGcmaerrwMNC7Mxq2DYToSmmzeasBzZPEAh8EsD247DFzBi6BSdrygW
ezZGnD1JnPdC+2Hl8a8Hu93LMDcaz5Hx96qCv41LtKjwf9BKs/a3hbXFYltvbXDm+jyS3Nb2fKFz
jN+fqJzxldSDnVFchml1Wg/igkO100eIo3+MDkEQ5cW4lO/wktJBlgWWNltc9/gec2ctSo389bmO
QGlUvUx+M2k7JBrFpNrB0IfIL8MeXj2WpzObbZlfOnEMNGFczzb14+U/n0YLl/Za3BsbWR9ppCmm
6sFRsBEYQJsYZwxEwt4gVbHhtC3gYHg6pvTHtcMcIzBObQlnM/vak9sL3yUjxfoNkvv45BSvkxql
CkdjEB586I7rWY1qUycQEFCRxqROMqcnpxjQlqsDcipQUgQJVPzsynxxrBH8fnYvsGPyzsDANHHW
WUysUBIZ0Pp5zEQcv57zwWDw2zqBt8MFgjkOBJW03HnxwahjSDIaEcy2F47tBOE8ZxkKeO/tVcKX
17aEB+4ICd/KaqRTghVDUnNm2dF6N+npu3EkWhYwWWgIdFPyoB7M6bTPg9unQVnAUwVfIB9GwPGV
u5FxuJr3DFh2UaOB+dhcZWQF28npzo9b65zwG1BaMAWIzXHTGOw9G6Lks132BoclOlbyO/JMekNe
cLGZxf0guP8JQsQ3fWT8OG4l5G1BtPwRZyYW4T/gSFE2XiE99gY1C9r1Lml2obhecSDcjCBnsNzE
edCHQ/Llhn8eGkqL/4w1TmeZHUPOOWok4RwjeYfoX/2R4DMoz6+2ETJvId5v6xjWolD2/ynV221/
kqY/YTp7f4pWlFLF8m+nDrKq25qwukH+6kuul731B24mk2oIXihHbg6lsYbEmGX9WdDWEhPZ1fx3
zlJXO/Jds1NxP2oJOlFX0MpWLxnK9lnJ/RW8PnO35c+IBiwz/XTJwSOmaeeah8UldOQB80dykb85
n2h72Mxt5FxTDHSXlEWvl0e7HpGSEk/1svDXK07aIL9TjjFRz8p78u1/hhGpGTyH4/X6KDDB43Ui
it+tbExqUHejRXgqfZhRwcGbIYmucK61VR7WCsJcssujzsRlUCMPSFA1I6JI7ngP1UQzVjHMFSma
Jleq1hC+eOIlFNy/8cGXRXfm9g2tSCwVuhoZF4UdGQxM8oHF5dTff6iaa+boB44peKJsuzmiJYaa
WyQ28GcjyVvMwuxfbVQiGg3jB6QqK6N4s1b3CRd5EpX7Q6dmY9lSEXFvQn7siy6Kzb4JXx4Jmrzc
L+DzZvpRr46LPjtKowb/BV6vszIP4IHPnhciCVCGR0991nlpk+8ZKdsftdahYAagnN9h0qC3znOC
rn7SjR/ahlvVt6Lzik/wcbrQF9l9Xxf+d1RQbTuOep7bIeGcoKfVH1hSfLMINV/+l5ciIYlOnrhA
z0IooMthCyhKjP/x32RfAF0dh9mplwycE+LcCbrivFcKdJtxbn0lZpzfStsexXGMLpECell2Ozgu
2IM+bK99mVdhQ7uOymKF+giZhftnlUYYX1IeUyKJUqTCyPPkavcyBXwMeBwnYo3nrJPo8dlPY6lg
SVzcivpRByD3FJNpEtKeDyCIn2bVprXUo6v2cMgub0XyBNlIjNgBNPJ230HWEfqB6Kb//1UhSUul
PqPdkVRgRZ02XuasULVZXErHh/C5Fr+gdnDlrPs3aBgN2G+OmNEfXVhAOLk4U5OL/nx0yrlZXKkR
KJFR6RRPQ1nkHqXka2bze8tzDMoxaLsbNvouvv9fWVdCjucBm6YHkYy1syrySA2FMymzny3e81S8
uTOrSLBozze0I1joYgWHcOGr30CX1lh9GaiyqxvRW8K+3OUC5Sxw/0rT9ipAXCLdm54SiBh3uGJw
FKudIQtyJVzLEyrEKECcaSNaEKdHEknFBWVV9h//s11KX2gFQo7eDE/QswmsjjwR8tficGfb89hi
LLKVuOrLUc8M680iFVy42FjDdu/QGKCptiOe1D50n4L1lM4CuuiLYqfHPzPhbX1hdBNF5IgwS9fU
4Is1AV3pOsMgwBaKpxFNtAdiZdY91MnQucyQRBmyVSyGm8m1KOZvgZi9UFNu4Lho1pNeKT8WI3+H
3yCd5+YtKBxW60gj9JS1rPV8Qjaa3yp7Sx866ynePXvMB9lNe2B0GKeVG8+VT9+MnfIOeGoP+r81
o/zt/+7QV1W+KveSS/0I3t6sVOZHky5V8oX/R/v6iKN/qbpg6N8cNUa1GPXqSISU6ACXghCfsqJh
+Kvf7cLuPxlt7JEAdfoyupZRmBgTPYZDyaENT/dBmxZPHn7gB8LgBTaLUsxYKO/JFO44kX4abMQl
gf0dDrAcHjxLboxe7xn2Sb3fG+qXFcAETggQPEDw8dotOKBJ3c5X0WrE6DW/pglujt3nQcfVcZ3G
GQ4oO1s0mDTHQqZl0WmhmPrNecVGULTHRVmKxXBMcBqMBnD4Mhz9FutLeDXjdr4z1cAiYwGAtxjH
2jU69uPMH0DacKymt4tf+EirrrOA/DhgoZ+lPWSlQdp/rcot7QUYzbex+M+/wW14SGq6ittW5LRZ
U5sm7SZE8roqEw4ZCk8KdiPDb+WSkdp54/XpjNfi2arNvgsD37n+agx+JCuCrWrJ9fyTrhTtXXdD
MbdXBt/wyCELXU8nabg/jbHEZa/DpNVvShXqNb2pSfD2Ci7KiVSNvzc0q982nOatrGcvvrMf/RvQ
vnG3DpnX9x5LGA6Z29yuBA5lD6fabLhGhb7bJZoNbykTEZWFuW+VgoPnv0BOs+3m9hjLKIhpAafb
wbv2Ls3P2crw+llFnADDBXzmiMZWiYVU2UBI5hqFp1YzNVo+RRqF8T50BXyX3jIAS2uTw07KwZRR
YjaNslnHeBwt/WoVtJGMHE+7Yh3RPp7vC4v44uqWEdYQ52NM0vJiBbvJq2fLJnO8Rg5ZE5oIxYaw
REbpOoZKqSNqMpgiym9JB3fJce2JVQxto8Wr0Soam43BlJ+KLqSAhKE7xeLhmQSYfZooBlB6xrbl
FO8CYM/4XBu96FuywNOTxAhUHNnuND6sN8GQvYfoUTY7Pi8QySm97OMTJLqCoWnqifjkdHHdAedZ
EUUb8FNiWttVe/E7PtPfjJLr55HF/VYNj/NgZrePemS0qNocW86253YoZPhBuF6InUnOkZAIZmi3
1lDbi1BU3dLxWH+F4I43sChff7DD5QK4kqyjD6hoX1ZE532CMWR3ynyDfPWHZpWwECOVzkQuDQli
kk7n1yqxRdJa5RxKcHWFQHWfAPXu5eU2bNWNmfATmBurK5yfQXPuuxOidmmvrklt3OCwF6/YkYCU
xeyG8TXENskZ8gBKD9GY7Qngt3KYaw6SnIMmMQVKr4jgVkAaHa2mj+syF1n/YadQ43piGbHbhXAl
gV9XuddNOeBBLDQD5vG7kbzo1arzVIxiycLGLN6CCWw+qDIXTabQsxX/21NuVxlVzQMu4edq/ou8
fnnqAGhLhzrzOV9uUiMUHKAoQRvG1T8fhen8OSZM5W6iREumC1TGiK79ZMPCwk5Cw4e2mIYMYioZ
rkTQmZpWNX3A0B/MlxpvnDpyn89FaOW8zqPMN5cll/Jocz5Jh0bZG/4KMmrJi5XT04N5u/rqjeCY
AsxnbOwVVL/sJUpVK7CJsioZSXS3k0H6kj+7p5RTBRiCWzr2YxAjYDsiMhZxqMct/vOXu58YqSXi
ATk2B0SnSrqBJXL+d2YIkkDa0UZ3dxFqmEeJcW514MJAC3mhtN+VenpNDP4FpxOC3BD3crR3ja4r
5nfaqjqAFd5fjG9r1wYFLvygpmDT0/5y6uQ6ixFQrMcsX4/q5uIiYX5xcR29+MrZg7H/AYA746Jt
WvGlgLQUMVjErc60XT0S8tuj62wQRSy74M8g/n+w7AdF5OxUOtUL4rpFkc7SZBMb11cEn+yTbDZR
cKAMeRYeoC6zQnbyqSw7J/xUPPUvPyc+o9o8nUydbEncsgSjiUh3x5pMTBJQYB2YbiJaIz6CAVtN
+T0Ib8W3jlPi775+Z/Xk/71zR3MnwTCT70YP5OHt9+4XTmCi8fV8gp4oCsC4d3r54DUSQmRSfwqI
W3G2LiOfjKtnFcsYyHODKGHG/rg2l5bqNRJ849tNd7gfwJZTxUiZ+Q0aaNmlPlpyKq3rXzfEApn1
bLW8bdrBdmy0HgsK/RnN8snN7TsoJjWvQOXUOl20pLLZE7JI/Saw6ebLfYvRCdcDZihvC0lmdw0x
xeAmHHnkAmErcPE8wNl7JOtszbB7zIn0v29Yc1k+PXxyxz3O7IPZBxfr9lJDmULitakihS70Yc0F
lVGP516Lf2xMdeIFPCED1eKmS0aga150qU3xBY7CGE6nqaK/xfV5W4+MSreGellR5j+FjiOTvATC
7cZulqlvsziGXBfJtUyXkPaKjyqgLF8DdddDpLHhPR1TaaVH9ryCTUX7cwiDZxGVQf3y8ODqJTB9
OeH36FzrWz1NAp9z9Ir+jI4p1k9vnDNUe/jyKKhNBrPCGL0027wJyVR+96qSzIAgoPAjpEwcutpK
1hSqfiqU8hBLbFpfV3gY+JNWl7uwqoGCyMAR3JLQ/3FJLMdtohbGqclIFCgY/26+h7UI9fTCVzhu
N6u/ccL0fEfUn3pxoRfK6niqSmL41PPBKt+u+1Jt41zbIK3DsjTdQPauVuPz0Mf5r0YeJTtkutdJ
DQ77N+r7md2N37hVKvP+R4/8d6YLB5rEVhQU8+ICvUOeW08wN0PQCvmWy8+XKASrdt8rSx3d3ncL
63r1SkJzmm/BughluMOo2n0bmrTlomUFFqHFKoy2/cubZrbRquDXWH48UVDbg0cnHpA2zCAlO5uH
EKFY+zsSGJE7KZRJiBarfS6ep8tp+fsVZV6Zwpb+vPP/SkqXWGFovf9koTLO42YqrARa++9fwhRX
NQDLoA8usSH1G/VlRD6pg5jdoVShCt5WEJRQWZcUyIZ7NjXY1mouHMZ6uvLFURnD7hMcld+0Pok0
L7Lq312+Ao54XzWOHwoGann8NX3Y39HFU5Wlubps2GNCGPQA0ChyIBuIaVXqwkssOURtVZpe3idH
tbYVhZ4krT1rg6cFpcHPOkCVuyhDx3Xn1YeO78vwewH6G+84JVRWGVWJ2RORzg+4zNb+t9z7qud3
Jb8/m9pjny6xjmwcqOoeHGVofK0B30NOMcWBLTkf82x2yKrWOBeX2SjGIlZih6P/Sy1CEMk9GZj0
QjB1hQyTOzpdzAv48jbGVL7J6LV7G4SocE7msg4VppB2DX+BVgRXf275RAdinZjUOOcRTpBCTg9v
F8Di7PpfmYfdolXTne3kuV3ubdQcGFrFDjoB2ELSV6nQ86sR0jPhTZrH99yDqdjRq7glf7iqvA/E
ZgRYJVclFIUCMTmsI3UOi7IZPMkvQwgnzC28KcruwdDpiAQ7kajTWFgSRRhC+nS/Cwq7bOR/eDJO
hB64JFzu5MkmJSoJ+b4yIydLCaPIcjdWQZgWYG8uLiBCeGaVrp0fAwvbrMLHFi3/5UWOmn46INyh
z1oUbiSdfXLHCis+sn5uI4jVEPaOPniogGMKSxJHGUt3F8YYC/eR1UloWNKEZkjAmMRMeU8Ld6Zc
z/gIgKGzku1vy55Na6jSixubulLC3Tr2OHHm3u1Azk+vWPUCHIpYffpxeIUqt93T1t93n5e2g0zf
jRnrUzxlBV7hy8MGUywlRdWyjrN7kd62vqQMkXkk84bOp+Wfy7wjp1KmVNlDVWBqM3QyoeKvpWak
91QAGLkLUTNp5U+Kd8SLkPdOY3ufS+oZ/u9vfyIhEv72+1S9Rdu7bm/Fci+1/uYS3IL1OznP2q9d
KQkbZwuFpCRsdcwtjUZtq3FYUg0aNFFmRCxJxUyKAGcpXjvMlAR4pvGW/jJAJEMz0u9zDhaDqWK2
kPJ9uY0szNgTmI/CCf607nX82VzL5x2UXBiTojwMv8mf2iXCLCi5avNaVjZPvTUcostwgHb3lm8Z
NPQsbH67R0b7ni/77KVVVIMmnkCJ0opF9ihXZ1YybDa7NvzMWfDVDPnGyJVpWvUstymCDOTPSf4H
7TXQOew/Js1ZnHkYwG87KZzGHDyJdA7eNrODJRScikFBvX2Y6tSxFVRT0TxlQavqTZGQO+uRzSZt
5enlADJwoNr+aaMW2nHsNwm/NEBOaA0l3RRN871Or8eiMbopv9vR9a1CEjrSbGw3zzh79Krw4qBY
iRoQ+NkjjXr+ToQd59XHXgBYBVH/kWbQtd4jrbr0+sRDKv21qZ/k8NjTK/7jkxVndj4xykkvRvuD
FobP5RcFxmQ3o9W78s+RKKj70NJGDIQtKPOI+wRZN+mBNmuLYaf6xzChENsyV6BVr+7xrOKsxqpB
B65+hZ4KIu28NtilkptEYKpg5lmoBVjoCuqAKrCSfDpvE+ewl3tRsKjv8LeFEMoflgwxX/M9XPxz
4WPe3XZrc1EW1fLtiXDEwZeU/AUkOpinlAyqscW9y7uvrsu+H70VoA6jK2/KiXQa86VzPqncnL2Y
CGFKVPrqvjQd+AseqANfqIVJ3pCQDv7meCFbRqP7HeFQe5v4BVHNK9hj6uu6/ftM2BaVlAQVXb32
vMimTtywvRXxrawFo45c7qX6+zMip6USecReuM318HJ1//sWvt5sel9fc8Qho2+y1EjHY6GLBmAH
8amDsAFgEabMfHwjNC8NsHs+8h+wRRexspXFtbzVdZCYYhWm8fIMnkGcwvkTbAtMrW0D8sLxQEtr
tVPOL/GbK4z5SViWQuwqpURur1GjWx+T6E394KcIvpkq6IP7EeZyvbyJdpzHEjQA91BzgzjEchEc
RwFiPYIUBXLaekxfL2lnC8w1nh6Zo/SEBaW2M+14kHI0044Lom7epK3qpmSlzDCR0uzZTswze/xw
Ku9wwxTuf8dHs2nc+1ojsWlPhCKs8r9MWsTGl6YP9dSXb3z44evvvdg/0jwVJ/CVFYl3UyQ3R/BT
a2j7A5GnREiHY7vzz2ve3ailx7RKWU6gFJKtOaiKbRv2eLV81OBA7Aha9ucueyIid3UEfgKKq2X7
KycFMkalNADA2LqV3QfGbyD0jGQBffng1UuYDOXV0HKJWxd+JPxtQxU5cEbhXLYO1/7Vc7ce01Cq
ZtYXx6Ss6i/VwccVKx2IEafBXEmOJ/ZkGncmi55HqxOefd5wWFSpiUcvTEIPSAh0Ip055zEtum9w
NLNG8CWtW0+oZQmnpewR7pTqfwHnLOxCQRJ8ec8/+ZFiTC9pUj8Ua3HVNjdB1mxuw0OlkbVpfmcm
iqAX7p6e21zx92dX9DKnAdFZn7e8RxvFgfe5rbJyzJidlXUhXrUUsphzZg/+8R1u3hd5PrrFcjBy
rsIqKVwCJgIXEbCs/YItMOm2A0LqgywbTzHGEeLr3OMS6zq0kfEuoX1YhMghiwe+GQ8W6Au8YGwl
FrnPxk+lKlBDol/NHDEm3z5JxfCU3HvANyE5p0gUdbHDZFyUhyOQCzss+FDppLFFOjSTbJPgKO1b
bq1cA9d2scpYVt5QRohIjp/EQGjsBes80VQdZ/hjzPDuLmGR4n4rDdRlSPhcfX1fPwYBbxKkbWJK
+coErpND51DVFYMRq3E/jp5CKaR0rXbbm1hY0BIhOrNZPgQuUy14XkMADw4xCqnGM/XixFsMuizt
B8BWHYBIiltpw48qFeoS68QJfbZRFdtyPxw/cwWe5LS4IK1QJ697VGx5g71m1IymFvHatO+rM3Lj
wWoYLXlPGTZBbN1eeNpMCsXNIqLN0SVxPcXiFm719vnm99s9bAgu1HoYdNPFbL+FAfaJxr3TQvMw
g7NzBGqN4SGYHQZPgPswhH259Ewew9/9t1vK5eb046MeAQH7QggZm/hZpZxWy07LOgQf3Q+uZnqm
+LXThcUrvSJ7UnQxFPCbuAAtYXWhxSB8uqp6nHqSH/pVNVKI/3DZvTrVghMsw3KNHPk/oMI78SUO
U0nJBgGDg+/Mg9pXqOfnwQFwCStENU1r7BUmrY3mYOZgvpgzJbyBlNPJzuBQhJBSJnJNppbHdmhS
wAXLKBn5+zFVFP9faqlloNhZdsVuVyAip9NwJwtTNeF++O9/7rMXoxaQmyB3tqEvezsWUlrlJDnX
JRlY6r8mYIOsoRB3LL1BrDoa7bYtpCQ5X9vUs4iItxHgAfszgU7ApbdwyvNvDo/4lNBkNghK7r3N
HbcdNyCjm7pSQzPc2Gzyer69RWUcTJKeQALakSbaoTGYnVCX5FLLULyrqmRO5wEVk37PBq9wlDMG
9OGjwRSc/1YwafbrShAYTYJ51K3nA19kk6Pg2aTgQuP6bSTpdK4lS+GBRPMP4kyMnEOgWxHLDr7e
gQ6nXKvtehIM6kPf2KQnWR4jtMu5sHpxpvQ+s9IJ0rrgAedvcunkvaJEkmOH43g1En/KSW3bcCkg
IvB6M6MRsz4qYp8CuOw0U+z/+H11drPHxdJL2tQQzRlb1diteckZocrZbgKKddwTwxKhBTl/Fmif
svszuV42eS4/BzjVDSnlnsbYwBFENk2iFS7ZDIc5TUDZa5nGDxHb6P/CyS1Xgqyy8PRc/TJrIR+e
QPbEgoHFuVlleRqA2AAY4xKwJa89T0RyrTi3KxWp3h3duwEihyvk00sFF7zKOQF+kUH55Xnd7gnh
OXfEsT4Fd1Caxl/ORzspZxHcns/kl/koELD8JvGFojdXVwiiOkZ1CLPIR7xHb+MmYBORrOUXsnxU
zi4XjvldAtFEEb5/jXhwSs6uw84EDJS9D/aX/+R3LM1J3E9yXJbymeIv3erowB7g+DhfKD/M3nKA
lqcgNgJpAsCBHm3bpTNUM57cqhHhJKk36VAfEeyJ59FTIv1i6at84+2KLOkjQS4t7g+BSgvl7u8j
POyiq2uEoSIgD9WWRoP3xuND0xdFU4xxxsMbKXB6rnTNgOTHK7bX5UZTEBmhby/aqf9zg6E6tcEd
xCEPH6/rZcwjuNqmfKAjCbJpU6Q2LJorpDbVNdJEhzf7vcwxqtWyHX8LVtSE1rjpTh43NPXRuWSz
8UnhkStegF8rRiikY/K8KqNGmzaAXtqw1WYokGyZaz8THo1mhr+CiPPL6cNltUwm1+fIFTqXIXVh
4hpyXnmB2oaez08wmMXUxVtq5n9XvPcOJIQs5lISBNinfp1RWVJb5Oj/SRPbrPGc30dOKUcq4PXa
4O2gmZ9FLNNzpEakbPkSRszpPt8x2xnrVJ7ZQ2urtA76Z5qQSOWQCSCSwNyeZMjcABUeQZtBRkqx
LxdYSUcPI/X8wrs2qZM3FZK23TEiIccYHrFEVXR3jWN/2b98uIMs0hxNT8meW2UsKf8jIcfTJsYE
q8jEZWJHGUpqyuOaB6D2jCDRE5IeGb/pfuf8N354G3C/BpH3ibuufIlHy2bUX3Yv2ft89HctMCMb
j1dggxHRPXRU9K1bTeJkIzpIxjQxaeYAnhGhUCvmiajr8nxk23pYLdqeL+YRJ2Lod66Q0eBbHB4T
t8WbWo0vl1pdTEJ1M/idE8yo/EnUCSFr8qqOIJF9BNBMwNGfx3AF93g6T0JtP62IF/+gKdEzxhQD
DN4Kv7JJV7/EghWroHbPDCSyMQe9HFApZlYMh1M6x5VeOMgYgZt/UmUoCdJMcEqSsqRf7aaJ1m8l
zpml2shxo2coQvUIHQ+EebYIwCW9ZdCKzJeRx1d11Li8Dh04135N8exquoiXhkiBSQf9raAcRjjN
drIQjUVSEPAlUbPPXIHRgzHj5LSeTyxBsQzAsk0syfCT2C8dOej+dcxcPR1yIfQTgL+Tk74Ze6sJ
Su1kiOZkZXT4zIQoe8ovB7ZsRwh9J0/MsU2exxbbwpGSmFClW0aN2jk4A670DSkrfu0fI7rdSCNL
68gHKfDjQI3q9/fRmiROwc8+rlEDH7NkWktV4wOGGD2WbFAle2rgSbD/3N06rWcDQBMQM4slcK6q
+VmyEjwnmxGOh2fgk64AHJNA1NoEV3P/8vNGjo62CTVqf3RraI98b8yIkiiOhPcec//GU1J8DTAI
kukvZNGwCtffJvVhp1QLK4v5WNfuANlCoPs/o4XhbkLdc9MBpaTlIiuj5gjOhGdtTuIpKBWXRBYf
Cex+Tyap6apwD8zJYJRXxDBgB5VVDKGCfWIvuCEqKPMV13d2w9v+4vV4vCEw4A/Wd+cr4RLLLzba
f8j0Do4E1zevIJxGeVZmM7thF5Q/DFU2it25G5qr837RBJp4WjQii+jwqIYzZUyReH/DAONZv8Bv
GgaM9iFcWfxVixiMgEO8Yz3oyyzooaJaduCfBMwQExYt2gjC/tpko2VSgIwl7PSJn72b0gCnOGoq
uQHROaO6oIZghmeGODoTS/96i+lfrcnaSKc74dLxwgzERYb5eMrlodRD0NHiPCAXJB2p8KfRr7/6
2UhIJ0UclYG+uH9o3NTR3yM4vSlsoeaEnmcQufirO7QYTgf5gTlXRqghd41jb9aWi2TcXUtVck7J
oqhFNMoRql9KoKiM+WzrOi73CGf3xqeJxrUrgmFsd+6pGg+H5tloO6xDtnfiX5lmX1M6YVVfp8SC
MRbg4X5d4YGf7XS9Bvj+b4uD/OTnru4xaRiV3tLsMWG7LvIGh0VB2uzNmbfhYY1NRhpIMc9JwDPO
jI+A+4c425/x9uEyos3QYEVXKSSlPXFzaMSWQx27+Uc/XXYjk/kJHuC24TOEfEbGr+bf5vj4gfCs
MR2hJ6mtdPisXMv0MlYg0ftB3GDRxlm+lLTvSgks0xtjBOiUPmeLtLHCtDpyj3rsNwTz0aVSWILt
NDiy+AecEkPOlr57ZubRakGoBWWvq8ERgb79k9VpcXjqkVX/rHsFiLnmq0IoXaHVlJv0o25cKESN
9xkOIUTPxZPm3Jmt4ykH46DysCRsema/7Yow051zQKxvkWrvPMUXqwoeW6RLG70axFpkFMthC7Tk
Axbiy7Bf59kfv2ciIWpIq7jT3lPW1HktipU0j9kJ/DvmjKt0zfGw9eaeyyz0Q3pDfMgW1Dtq/CBk
KXMf1yRJ4vlH1jIAnKAs4sVc5XDOgjsf/o3mU2p6q8pSV638Q8r6Qq6YtKQJxP8oAitkHytJvv2J
xQ1bJi3/7Js3K6FqU4iXmeE2iOd+Pn2hRx8AUNzC+K7b0uFVajiKYrQcfJM+B2x9xt4p8TiI4XCD
A/CJBGaB94Lg4ZeDgUVHcK54z858nHZzIJUPKiZCACIBQQdLwMffdP/tTxk3swE7Vswtvme4YcYn
DkZLXHGv/on4r5EwbfDndxcHbRkf9L0SUBI4EDhL2K1sSvkVZpMNdnT4K1qWmUO23h+LCRjsfovs
EnsGkDWI1TpnP6wbYzKUfApXtouKkDThSSZQU8AX8xLFxxxnq7pXuetM77zh3gAdfaXPnEnOX+zL
UDpqTL3DAyHMaTDkiX6+QhdN/QOb6LfY8Etraem7hx0rXPTMU8tMOpDvf+L1KEwdTO3iLMhCFpuQ
zayn0BOTX39a44NR7xxHJMgiFEOteBdvXZtdpWo4AM2Nj28DXIwEsU1fCyQyQlfh51k0J4D0RDhL
9IoaS+rEQjo+9w6pdaYReNwFxHThzkDR56dBxB7dB69w3EzNOdM4/d1Ox585ihhRFJf0NdtnRgWr
xNTKac0+MwLZmiKq/Z28jn5NIaHjBei2Sk+8tcL7WseVU+a0NX0vwbCcu8A9I0VRHYu5eGCiXrOU
k5TtC2iA24v41iAhnYvSwrYfCd1KL98ouSoGzY9Wy5kHmU7XBTplddqdaG0loye/ztPA4cxBKx/V
45YnWwAaiFb1jY9bT9/j1x1vw85KdvbkRffEnJg0ez8BLmx/aRGx1vbLte73Xp3SKVsOecV3zK9C
N/1mYMC4d5pwSXu4tt4OG7p/pAAMcs/rbhVFStH4c81oY75htSHMLfPcpWq1odRVbJSnFmOHrPM3
NGYD4efcqmpEykuc5rRbBZo+hYXHtrwybMnLkVMAZPvAC0/yp8laBANu5IKwyCYHAJXr3Un11vTc
2EF3Eno/oyNq3BBSjjvbqe1De0//SSVnzUnS2VVek6UiBvI6qG60DZmVhbZgg1B0PMFsiAZyes49
fY4xGghuj/Uj1HjdlG7ZMG+jfeNrll7fihIgbS2HFx9S+4yMf/As5MK4zOiDiKQferdKS6PA3CvW
gm6zUMhCZi1qNNs5jN/vs3KxNapkJdhXwgiSsV8xBHUS2Z3CzfVyM8GvDfoo5Ey/LtiJQaxQHGvw
1kawiBDRUtGTcw9u86htYYiw8CTPPLh3rhLspMq2X/e0YeZ7GrddEJoOW2eE478wW5RtPRrpPYO7
RnDeEQlt/koViS15+83yntv1CQTea8TFTqHwGpNbd4qYst2BhmogWpdmlHVBFjGa3+yPklP0upwT
pa3miBuYf/3x1Zg0Frf09LRtDJoARVZS3IvtiUfHcr+jZtr9mKPhapJU0ItXk4AEt6yh46elyv3A
JGal3DrPNAaLTHAH1IAjs6DKZw3ERvXfCh4WJbzH+3nCcZ4kiYXiY9kFOkO6MyaUTG0SnzYqen8a
nxp0ak7AxkG6X5CU7GA8ycxWO4MdRpM/sLZhoi8brsKR88JR38ENFX+qPSdvhfT22Fuz6hiMgCZy
IgnjB80Y5BQZWHKUE7p4Ndk0Yciuh19B5prhUGk/ikPcmgAEJJyvFm0EFTxBGsLZhRz6Z1y/GoOM
n9jHyhASl/kNr0+1SKAIGgO1CsuUond4z/dnjYeSQbhmN00fgCr6vosj8YGNwZnqW3iCZevrYCRC
llGtGPMX8zoConQjJslv43qI+pyozmhEYoiH0YxzvEeNhhRWeNmOu0XmWGiAjIeoFSezZftbcTYS
w6l2Smac5TnzKPMB1mgEZa3O6ZuM+4wbuNQ9sKfRYZO9GnxI4IsJ/VD6umWYTyHgf+QZDy+zmOIT
nbA7ZB4Vpp8YwlWPMlK4uXuufTNisDIkDuAKiAd+KBcoVuAgrvieIqdlnwYwNATm4j9pBtLqDpef
N9LUs602Mfm8molt1b268aBjYhUcl6n1gpVssj5OmC4EN8uzfq5sG4BUctV/l3AoC5FT061qKvyC
01C3keYWIyErN7pDvEsy+poyZaAtnM0FcZkysSRIuKT6OOkrKVLGWGtflT3eS2fJcPSRStwoqcJ3
um+UzcYVbXuctorkXVUcT2cgx+zYtjwDDdypSaEGG+8fxVEXEUIFLL0XVetWn3BrrX08h5e3BM4Z
1ZjwaR5InPL6y8vYICG912BuuZ96gB0IdQadYWzU1S01j9ZV2HOBGt44TBk5gtCc1RROgOzdODAe
yV53ukDTe9Y2+7IvXJvyqaRCwxEM6GvSafaXdqfwET7CAJK2y2Zn91yL3ecUmffJoFcif51owXhr
WGFNQX5awDPTLqdM/SWPFOynZG1Ugf4xjVMz7e2WOWRdIiiHW4mBHfFsqFfQ/XLNDZjlXty8ptzv
8Y5vSdoHThJTyUoFnMfmuZbcZVPMX1LX3l7tTr7ONw71+O9qCyPaIOf2eS5zTMoU7Ue4kImL3Xvy
m+b7yAmQZ5b97c4yvQodYi0aGJ0Y0q9DAXDIH17H9+9lfC4R4as8z7LwfomnPZvbZBsrEdjvJRLn
XhD2AIglBqijqUVKVfEsGhTSbB4WbUsfoJLjXvzHjmQ+cOpOhDJGqPbVU7VjYOxPW+Fxh15tghym
v7l+xYxe2yzvY05J+PwOPv9sbYeJfBgoeoQiocE5ZJdds/vih4s6SfGcZKcpV9GjL1I1POcxGC6c
mPn08HbbOH/YV9XgMeAviK0SWPOefpKAFYAj4TXgGCLZ/AdyqO1vPLQ8y0Cbha/t6qBehHADO188
55KVYv7vr5DS2HnyacE2jPIuDhWefsyTtBMXhJArlSSdzgk7pKJnX/rP5UcsOOG3YSqXfyHqm0rI
01GlX5wPt4yjsvRwAZQh+v5Gv+WyDJgNSfHcJg5E5kI0A22EUrJZN8uZQA3OSzz517N5HWJNR0MG
bmn5UjWa8JPsm6RLSZK7Zbdxo4Im82MHiU9uf5NUbAlt00HT1jP3H1bes55gpp0X1SMFt5BQiFpB
H4K9S/1W9GC6CBaNwSqbFfS/99HXzpRj75IuwhHu/mgI9tX3ltK7iu1L9SpLNMriPVX977UHnkVw
2thfKOthaIkV1yfZhlEF0IS7VppLJgPaJJO7YOsJGDPwywMb0xOX17wdfQiatYxkhAUToqSTZaSx
IYkz3LQH+ViuXuuXqHvsOI06X434w3P7BQl3ZsAZoqqcGBTHE7l7CZhYrBU6FWw+YAUEWLt3mGz8
ybNjlix0SqW0UQqDvdZWZ/RpoABcex53Llw4LUNRtxG92Z3iyuah+skLBibU/biKdBFzFbzlKNNZ
I1yyCv0XYghd6j81kzrDffV8Ap+Nav9e31CMfxmv7tzij1Wd2kRkn+z0Xg0zv9jbNBaEIRuf1Z84
oaF0qaj5OTqI9PqNfhPJQsbAqMHU22wsJ4OvXkcBL49ROoc918x9bcN9hx2Wovf8tnAlvaGKxexc
7waQN073MuXmNXaRxptbLh0XdTyh2NPXhvYHQ4SbbI/ZLx5xaVsQE7UP2NFaT3Fhwa02kGfzUfDY
J8DoTzvN3hksE5iYar3DMOynsTP3YL4udHqQUhV3+70FxujxUOy+I+0l/JMT3x2T/DjvLK9l3xQD
iOUgchFaLU4wXWX4ezKMTewj6Gw3lwpkQR+NLIt9rW5V76SpZtRo08atMaPJyGyifZi5C5h1IYKG
fisfb+gE6qaRqEutFz/qHar78umJPw9xS9gE49fGGwF5AOPTv82wU1S4V0L1/dB0hjaTtnjM0ysT
H3rsTxQo8ycssq2weXADURxlDHN7ol5ODVlfRWH1E1aLO6op2ZMc61OsFgX1Ln8qoMbRS0BGRSC9
yAn+F87A7020uhLDVE1zVc9WsY5Jq59OrYvYK24I/P59WYhS8BAeyDv/iAWbWF57Izt+Sr4EQ1dW
7uLQUYZga3O89IartD8t1ojjxcxeUjtc3ek3oci5iGX6BVSsMKjVJFZ2dSHX+1t5isenuSwvSbp+
MzXYvFEFcUmrw5uycM4roT0BPsnwVWrGqAg0ilGP92P8AiDna/zJx7wrK1vfsrpA0gOBNomrJ7mn
oMnzV/DITL1vpvqpSrSCmckVB3rUem9HFA6zQgRblYe1qihlUSDK/vEkFAl5I+7ShRL0i9QJWfIf
IL3HrJjwYCG/5UjBvB84k/H9V76feoT+bYdOBbZvzYVAlcbPKRiBKN4EHRtPvW4GgYguLBYgE7Q+
RdMSfEjieu2RQbS2j3W26hXGajILUkaFxJjJcdolVnoWHiLb/PHB+VFnYD/5B5JUN/3g8GZVKwtF
Dq9JKChsbB9UOMHYjNYL5RWJ2aQNTmJd1X8+7x321Pi1e5PuuO44MbQQ8/RELOqPPxugJXphkcx7
T9MqpJhSGgOLvYorSLpEyfinnhP14rtYVjPdQu+LkQksWcRlig/HMUk/qO8UXEemVjxBXmBMsa+s
NqM8QZOGEUBQ+gMxvJr2GVNsuHCjywmxur34EDv88IKRH7BjIUkSTdnup3QfGsea340SxQxBmAb2
EYK7xBRPz1Nwy+Cq2ALKcBMtpjfNyNaIiXwx5AGdRxSdGNyw84TxCGkW8X/kB5IFG5Hmka4Mm49B
z/sE5Bg3MB3c1KKoGh9+SmIwSbGzhNAo6JYnkcmXfGhYsHXJE9hQfP5ZoeazXiykqW3ZIk7IR5Hl
JAA8e/DQw23VysS5oz1vCwKcbF0fdo4R0Il6ppGgBAhK2Sju5VKw6CfdhGdQSWuyDb9/7d9Vpk8v
3ENnipy6Kbpw8E4Ie1M0gOm9e7FQjyAvP+75T1ZeyvWKbgxWUOAWhCJWF11fIZ2pZXo4MsKvEAQv
zi1aKAtRtSn35v+RSP13vTnty4rkbdSUjFM1ja4UrkhWuBEK+Fe/CdXNQqlMTvewfX+hT+yqMLS/
pKBsl2mV0twiwmIlnA9fUsUcR0ZHwEYfNTyWtcQ7fPBo4BOKBb58KDl+Hd2XeUuE5TMNIIaqklQc
TP/scBm4mrgtwyV+x+Bt04keaadGkpWz3bXlV/ZCAj5uekY7lEktlacQoEyk9LOyGHXouJHzxNBU
qylRM90b8x8hzHE0ZXA1q9HC5wzL4LWEBHb8uYXL1DOMLnO6cEtYQNs2TDiBRtq6BGlrKixxNeHl
JGq89gWwCzLgICbfqIjIVdCpQofciy4ztzHz8NymL3Z2xoKrrUemsm9pR/HA32OS6tLmJ2Rp2vK4
MTN2jmRsKnE3hFQaWT+QN+qktEg0gXg/p1opOkqkwcfcj3ODOTjIy1C3WpEIL9oRTUqo2RVjA8rU
w3QkzYoD05Ad+uW3tgt5wn6H6LnKPjXn2F7YVSOtxKtgzzowfedQzDD1Q2Ho/mbPo2JVZn3kco5t
g6RcEaFUSig6T36klMpBGFR+Cy0gUStw6rzgu/CrdhWHwmbApBsXxvM+SN9uzENUjbssOpqj9Fe+
8Lm5CmtdFceBZnA0ecuFub9S3DsWp+SupZEoPKV5FmYVxLy9mZ6m8BukcUwIR0qozVa05JLXQEs5
EwwWuAgfGdbiYmGHb6s1k1D19+kPPe1Kj0f6fX1jc4b+kMNZgrQSGqZ/zkFbH/SNI/Ng3EjM6MHD
qSyI2Ei3tzH4umAdEsanQ1G+Uh6rvousaaVgH3t6qagFpPlDjdgewJa+tE7g0TYVgi3bvbBmSsBg
8PG5Hbi3ggqhlA8vA9j6h3cvJA9F2n1U+lHoA3YefGtOw3KJI8r04EbgAyzzK41l+nLtAil+Lu16
EIbv70TAlC+8Q7fqpUEoU+27yXvuizFSmroGMuITDWuO/IehktM95RemYbATcAfvVnn/gDqvpyQW
tVpo22yS1RWnLyltsPXfhPw7ivpcbLVIzX1eeeMu7tX+H259FRZAyg3jmIBxYTIIuODZFOmyA2oz
EXT3OUlhcD1UsLl7mxYm+n6BVdzshWTcbEEqIww0UONDZrbgd64I/FUVD2WGTiFYIFGDjIsXOefX
Pm+IAIccLIwz2gsX9BgkFj26s/YXywl0AJzWdH2PeNJ+JwdMQvMN4OEg/ZbC/DgEEWpOXyKZ9SYv
1UiFqT7LLUwe5oZRu+Hj7HbJMhMWZr1O7+H43X2UU7zfmNBpb5bb01vy0LFP1sh6+oVD90LKUgC5
sxCJIYPOR0GP2dYGR4Jngl71qLWI9luU7k4bBwCT9EyJ6GHrAZ7c0/Qfa3+dBnX+cs8do6maG4v6
qBtfJzPYUwig5rM5g+MUjR6OZTRTtWO7PMdrYJ3zJyXz2caZQSr/omVtJoZKkV7tI1niiuLIYPBY
30Q24qaq4CAnRx5al1PwO8H/YRsCoxZglvIN6imKEd4VksZYZAbsLQMawnok/9kckXWDlQT+RpFZ
L01awSfHX27kHsBzSGLaZ0n1epSy0y8PoTGyCKFrUO1tYa713J0rq9qPo6n33f7ZQRCYPrFDQ9UK
xjP49gvZ/pdeaJMltI+asDZOeHyMh90z5thdIkRtsdV3cy5igTJUtCxzNb1jQiRGjr7O46bFU7Aq
BJpiX47fHdxXv3mKNJjSPdl+OxwhdyQMdWK6MhA+O6J6bLLhhfknYp4mrUAEvYaNNhChONd4m+dN
R8PzDqsqq2f+6ymsF8xP/dqdMkLbN+yCcEXJsKfwExKuNUQwBquIDMV4pOzp5JSnfg5HJIxa5jlz
4kLe8/foZ43VS/F33s65ic1DrIClJEPGjnTlAuX+B0JgKNAjbYQ0LuCHoyi4uGDRrF6WZLeRReDl
olpaW9hHF/xRouspf80nbx23HbmSWraJAW6/8ZB3AZJm9jE+yvVxoS+leDfmt4Cnman6m+psENdT
i1by9nw0OPM3IvULjZeAPFMzJgwDb454LJfaLHRwmZSoXx1csgo8YtD09+BUHE1EeOsHEsS5IU86
sKOQGhXe9KDG4uSktJ69aeXs083yZCdbGfDe7nRmfee5sE3jeus7uoHbmVyCWDUfza1B5pl8PPYY
k2OPSt4RsLzlwG7BON5MfRDxl0zRKSCls+o75TKCPPnHLmFSZyO9yyRUxnOq+zmhM+7xdATiIh8h
MJE8omPFrmbjMeTnXVkgCRzOt5vYOxmr1QOo+wdnozlQjhX5z3ddgY5QKyUc3P/CXPMtdoBJgQN0
0IMWWnDWBBbH8yiW/l4RPXDx/OmbnahxTWTskqermSOgX2I9toqmuk1+M2OMra6MVl7Leb9f7KF3
5A6hlGifEGb1FX/S8VSBKiSa0fhNSUdLuSKxJVPePJXkAbb0hN3wgD9b+bcvJCC9rme0e1UI1zpP
1Fv3mml9GOOyJWtyzMpX8HZYoFWL96HWaHNJ51pk2QobYGZ7oMzj9eGl/NqoQWuVsMVi+cFjuJ1p
QiWlJYOYH5SAPYZk1+IDbVBps4f22/DbfUOwa9oHxynEDq2MsJ+d2LFSNk8aoxbDIHFv1cSR4y7s
axMTPiEzrVP5iBKWgcVhYI6+VCq89KSIS/xsRMvP6UH10tfxzhrtjJlnl9ajUl0j4NJdVspB93/t
x5G/5Hzh52SMpy4XlEXhlyKxkkAgUwmcZ6kXzp5640jLl8ERhOqVXqL1nKnoaSq6jLZTlVVSiNIc
6lVBUZxxrBvfXtVUQqLZuF8cUa3iOJFUGjterVfXP6vgItiLFVwsYvNjGSfsr06sq07JMaaDXY6/
uSr9Vu5R0R4Ghk8+m3uyXVizK9I/mcfWOPQuUAsp+6fyNv01AOO4aMIVRT5LdGXAEYBUOpPq0kKC
+TJLpWiL4obbuQsEo3HEQBxNPsrZdfwhUz4FvHRTqMXFjYOU5g+js4PLEajhkSt2IfJS0SBOmLxM
eZbV8i8SouaOfabIeoJZsUPZu3LtVwvYiSSH+6kEH1kyRXhTpT5ZBwacpqmSWTW2FDKmEVF3f87C
KDYM1Qq6UAd30IpEEU1rMNT0Y/1SJeSpRIBqDhqSi5rnz9bZOoRs1cyhY+0bogZf6VsvDoD1Jpmb
99hLPItVddowYlZBCrNpOf5R+hqXPUsh/YT4QEmp42AwcgJtBuwspzPLkcHE+9gV4O8nUAoHxn66
ZtrEKYz0n7gIzh9OZ1Vwv9TJZ3MMM4oZWq8TLDZjaSXvWEZA4VCFupUnRE4zB++A/Lok8cjOQpo3
HnDBtG47jWlXS3v9N3XO5LJmtwW4GkxFuqegJ7o/HJWmLcdJGbiofuBf4npzl8GasD0L2PY2+s7T
uYng2iJfTcYLKXBNYAPwexnOA8ASF+kj3c41p6jgAKT9l3abZ1A534OW+NGdkroIDNQsbBU2vwzF
wBEcIg2UZlc9gU93hxJHKmVFxfnRUfKqv1puv+ZWUrl9Z6HtvHlI5zxNGDqyjFuQOuoVUhR6EOrl
iTvEQutoVuhYPlT0Jr4K00UhZkyAJ5N6PMFlnvRvduESAwO+cUYFtPMwEf9LfupXV79EygyO6Fl+
1abFCDOzU5l7M+//LNgfVr3kSv3JXoV0EWF81YKwZs8GmOAJwTO835/8ON8R0Taf7mWbANUpm/25
IHSE2w5XHpAyZoPoPIMBxrUAxWtO01BG+SAqFG2kgpoJ6KRfRyGSSt3C8HE1e9cYGrqQdQQlh7VH
GgB86M3AVr05yDFOADstS6PKAL9XVctxnFLefLAmSTpUMB/1icH06xXMIpIq+vj2+o2ToopIa0u1
jIe142eLwFExbvqwVgI58JBh0sQFKVAJCA7o4J8SkT2Ly6H2YF0OXwDuTft9phExSZBJRetXuk/j
VUzYoz01F0NJdi7GVD/febYQieo8w463vD3nEgjJKD2BUKKZAKISypztVv15/J7evqPpXKSnMnXW
hqee+71F8f2ZDFj8gW4nHG8MNGOtfyIiopVDkqf/txbTeRAWRwaNBIaiAQ6OUh4T7J3WJpsYqKGy
pdxY22sg/plT35v/kQtJdsQZ1VM2nPVqxAIC9meYQyPjMN1rfqg/t1lL+zvRr1Rs9p3nx1RnAEWy
9aYD0ah/0E8qNrR1oR/LsS+d7LKu1zR3+DesHg0q3DGQHB3ofms1QYM2zN86Q9ztZ/hvkMypYQrL
VMD4PY4N1yRuo84zoOr93NkRPPOTFlbrTQwV9wrJsjXsihy2nsNXja4LGXLO6Q+aotHQthJSlvpf
R+Mpf7wZpwwyN0letcL99GFCA4VeYFrEca9BiP4tcoL9bLhiBuTaEebmuO9iv5e31yJCS5l3BQO4
WhA6E+xKBdiNg+UlMNfWwpo0902eJ4QTL92eqUQlv0v8mQu6HTcI16ULtX7nMoYydzedo1k6ivzb
qUNSr5SSuc9xXR03kz2SZwq4yZGBsWkbmrnAF8OTVp9+33Gw/2XxFN3thwqv2IvRQharHVFcHHw+
ykYevZrgcvhwqXATSsQh9AuB8RZqX2CUCX74WPC20oIiSRhmYbr8nBPc35VtFHllCBDtDu7OsFKl
kW41TQGdqIZYg8or2Jk5NzCEaK34YQojz0GhFvamJXCL/lMuItVaOqXsIvqE89ZH1N6OdwBfDlIO
Rszecpyxph722OZzLGtXnRINlgvHORXU0FOzNwQguuGgOMqyjSJKzBU5pc9eN1Q5UXMpCovvBxGE
cQ+CQoE3zKiZvWPXoG0UTANIwm1UhBlz83QRPANDfT4zHhFAbcB4laVcNcS3oP8SXDZnj3ixov2J
73hIga9jqRBzY6m2t7g1sIJj+8/r2/gqoE63usbAV90+8F2Oof2CRGZPh0WSkZV+7QL35dIlLN8+
9bZ8pCkHXel0V8eFnx6GxDwDRWBD2g6cqolR7qTSu+ZHcy266MpXBAqriDVQ7Ib074KB+0Ye6zqt
QEU1glJvMxU4WncRlNefsu8LABPv21pm+IL9JBh8rxdnl66MfnX9inMh3reG+lhGc8H9JymuaQ2b
//hmf6+FHgEfvuFl/7P0IdsGILG1KQxrayj7FRHI943sJTtBdQ15s2eRvoJntTOnYFP0/pZPEz9f
GYyCs+/5qZslmGEL1MLegBB0e9V2kevo7VwwKnsWeLtY+UhnJFKX6BPtXVcXy0v73bNCeRb6OMZJ
DT47Mb0zt+XQQ7ObtOjCJUUS1QXyY1ZjygigUE6TCylVhI5WpTYeyIqKub0ITwhrzp6nt64EkNRk
CCsBZxBgnmJ2p9wOKUu+iw75EKosI1ykmKKMMRmlBuC7P51MaVdtC0xyCjAjvNLvfLkulVxStmPG
fZgB5AAauc9S2cHb37fsZPjA/AzJowFNavqdCN31JINCdo8lu9M8jdQoNCg/+BiruQFqSkHDe+B1
bF3jze6prm8wBtgvDkHQ2oIa6rRpIChx2c5QpnQMen1p0Uauw6aWSRPtITzd1HPINzVZ0E+PonEB
LDc9M5ROqfCAbURbq0irmZs2qat6EI3ZhN2pMkNjbrjvo/vX779ijeRyHTHSsA6M6px9MMTp+Emt
zlWxgbeC25LjgI+FIP0fyzD41IIciykSvZbX9u4o4v4hbdFDqQmOrp6kktSTKbFhoOvX96Ic0us7
tHhHRm5Ro5OighwppamVtHjzPyNNJqjSmg+OcX4pSRTAB0bBvVQZ7aBYf/8YEEAfR40vF6O0ULPk
6Z1n6q9e9LI/WEcNGliOhvYWajnQeJNGe7uzHYXWMk+o5xM3SxqExoBXmGX9bkfD103bXDWRrpjF
FeTKG+AUK4Yk5GepJuvhZybUv+uWvGPvzlw05VdViIjOPFjTXP+3x5bXXJYqXSBgrl9wKGUDZpBb
GBHphOti4Lrtl9EThdHee/I0lZuswTzf+vSw8PpUV7RCOmF2j///cAp1Dh+i0D+spwgCQQbr5PVB
DgNWPIileaXApWlxJvwDTfJUux75zDYEDlyLbIo7AA5affWhdzhNksvUd/cO+DxydVc0JXPsUla/
sna/tsG2zMIIP/GRLVqqsjGXXanHVGlbDktzqkiT95MS7clWj1YXJThV02eoTlG5KPvraIiDOksT
uXhZrun3AoVeYBOvxIpJiRlw5cxTzs2KVqeDXugfc6aRz+3bNbIaZAp0nQ/hJikG1fqSoGLGfe9J
XRJWQZx9tc4NteD9mp0LcgC/SaW2rQ6Knx8jzU+5kJmk1qNUIObprJEHTxxyPxvmMaIscL9QNMCo
doM+fFqbPZuUQ/p7aPwEfzw83R9+njofQSoWlMXAO+1bWM6HtBJvwo4DBPDszFvhtyU2rloLkDGS
dpVECKHelEJu5E7oE9egHw9C4BDF4CgKCVQpi1zzH5alwVn7scJMvA4kl98s+TYAI7OtwqJ5ag7D
zp7cs7yhL9BZumotZaD59G16IdufryhZdKFO41ovsdl4jiyO3ffTwEXWWndoxE89KQtAN+C0icbm
SDEaEe3uwMptpZQ4kPsZc8WUTsleTWogC9Qlacau5zrttr4MtcLDRJr31b000+jXvzHBuaYjmRoJ
RObRJyrPPAyQkM1oDOKqcJY63GdOikCVy+EDSnyrKU7OgB5DoPhp3B0csKnKydq5kQfp6MwYALGr
k7etOR4zMMp8fTjKDfVBP4Mlxez4Tw0rCsCM6winjUOwJznUhvwtrfgUH95fohno31gTeBpZESCX
Fn+JoYkRgEtS8c0Xl7KVZ1ZBcKf7UcF0gQn8UJKrKF63AkI1J/dqUpg+iJSG1HFItMqVzxh4Ty1/
msint7jTpeRHQs6zdf+WyW1WKTMwx66jY8t21uAgLbxBHh6rjtG2DkYrFzz5oVo6AhBg0uc/fmEY
D7eCH0cEtrocOCj0MCngEBOkmc6ugkff7MwwaGHG980HHh1Z8VKF6A0Giz+lrfIh1/HoC3rfI5Ar
PBYs8vSRZ7Pj+lzh9EU1gYwAX2S3tGDd8hOW7YhhhW6CKwJKfipZJI2mnRrUjW4T5eKQcE1jmTc4
ML/zDlJVO96VgMeXj9NKhhDGZSy5wJ8blq0CiiFU1Zyb+BAkCMLObBRTi2fhVPs/GTue2190mIvG
6fwrTqxZT/mXB+txsLKBkWQUODJNpBxOCGiyXXxioktP4kPh+/bpMgIBwOeFxsH6OyeFrJZ0cDmJ
GhsrZC6ZI1Qmor0gbQHEasbbft38XrIfOPHxivPXD6+gDYBemqJVH6HQ9KhWnc9xrUQk41sCQYwy
Ozoqmku6MxAXxFoQD7UZ6VGFYbMaFdNflwYyDjWEcjqXhjAYxSfMkZygzmL/LcxHPCDC1bQ9+pKu
BBsXPxgyxsqPd5LDbKj3VnhAsS+fpo+ustT0+KbXXs2q6OdHJMKgjASNDEeiH8yknfiAkQR0yzbI
s/MpD8ap4MxuxcJmP+xZODX1ikAjaj1xKDnUPS98zyt1Wa6yk3R7w6xRwgyek/pnYNb/RZqa8WDT
uEVUIT1PeNmbRbghKsUu+lOgMpcWCub/j9kh9RDt25V+g0WpaA36nCxk1vADwiF9I7Too6HM93TC
RM1b9mWtLA6BoOpi++Q8xEi6/d5wkjSgQxoZQ4XBuGtzHtOyfYWazo2bRaePyhhEk3cxX9zzJJtE
xofV1Ea2tj1udcba1S6NBY65y9IHb2kIP/ul1m4IVwlwZL8iuTA82kIivPqPyO874jVsU/Ptr64s
5yIWOuZ6b3xh3AB/OpsmPEUOR7qx9VeKNQXOqS07dKRQlFYvPLObhZAehYyrpIwQ2bhbwzAdk76H
f4KwZM819VTffVXl24tGJM5uyYqcUnZCaxtbF8mjtTOfh60EcQwKVwP7I8weGvtcY36vvruaMGMN
EwC/wb0O/EGJ93OsW6uk+9Dk8E5SwC4W4PCLKK3kytVJaNXOBHQtmJhyPD0i/fzTW1xya31Ldvh0
T3yqq5w5GBzMOiKnK5hgsjOWiUtBSN3rHmu+uA882OOJkLayfOF3j8vKe1WO5bsjtaKBGIXyMNUY
qwMR9ol3WHaQCiade1yKH0CogGwJ+Tq1JG75VvwrC7CkqqJv8yrL1DzzmNqkRTgfmpJawa8CnDr7
psUhXRAVxXBUYAQoNlc9Iwvv8AmAcOk2hIetYp7JEwRnPF1nUIdA1Ib8321IyXCoFo4qaUskJlDi
wn9wqb8Fggi/QR8aMcInJGPCTj7C2FrxjY20Zstpjn+W/cge01vTloGXDDdBiQkme2tVpVriuJva
TxVg19vFYqIehwuCBAHEBwR+sbVg7wsRw35BVrgODCgcHV074HAseroIfafyv0Ll1cBBHQC0JUlA
GBvHNd3zqrCafECo1pDNtyw5eIzbCM6l9YG/jlstCZULC5xtTDEEkO7VjWs/SQUMKLDCqNNTOP+z
a/0diI0rdOtYSbMWWdAXCLmfjYi8nNGW2FZB8otcnaq/ZhcapqTyRAr9sOylGKNjEf2xsMOUBnzN
DFJ/XSXhSw1oPD/cXianP6v+AnYbfE5ho2kp1isRo+JnvbYwkp4I9bVTs39GJpm3os00wFTdM4W2
RP8zdTD+47XnQsPQKI4TcodFf2fxfLq8EPH2oagMQy6VufEAHGlrcBLGynrlgUb4nxp2EMsxFIPI
ioomEZpmfU1zOmpv6WEnjGDj+OylIiNvu3OeIgX0arCW1kT1R0gbFWx5QLAehfHWj1vCu6RJScmT
bM+3nddu6G2mAa77Ek6SXvoltZg3rTviVbLUq+7Wp6OuTmJ0yoip3dlXUltDuOvWx/DRaXmGjpKN
kAW5dq4u8UANorfmAyZhCUeBltwyoKqyaON981bculI9x1UTashFQT4orkMrqO4O4yIGI4C50h/z
UPnD6AmVzC19k/MnHliBBQGqgvk5iT3xDlROheX9MYggaCkYKKbtxsBv6WdIU+Q+a16Dsmn5MmD4
sXTbngNTZCIa8Ux9+rCS+q02g5neR8xbgF0ZO2pED+uStndTjMbhfOiD2P8TyczUWC0n0rg+1K8X
9QMggJSZ/g8eai5u67cyjKLND/MnWHXDLcdVitJKm7g+76p7YfUO6THqh+uIg0VnhlGaxF2OLvYD
LSJJEwW3HZoIQo5TNfRM2K53Fvife1rFnakmiFl1A8cO+GkWOOD8KzoL4POXBWmNtNvqt4Zp9FO6
EsZzqhduIH/COXD1WaRauAKW1+SvdewmdKF/bsxHx1MSEyZk7nAG5el6MWVOXCLYK6n7XFt2zIHk
MOUVcTAsFrwvK2kkCYUORfhPnAy4F9kCBfAWj7DUrNsw0/yXM7ECVjqVgzngA9C+xNMMocWQSJMp
s6pkb0cppB6VkFwmjeMZRnJzOeoTqINIZgBE3TM/+DVHs7SxR8jQ9WhYnU9boKYb3UWJWkyKI72B
KCMEjN20SI4F0HScqMUKJgttS22MACOiIyBRDNOpoibIhVEx8lUeU5tpBe6/PBpNnMFUaWHJudVF
oBwZ8NF0TBU4K7+jrLkYLEyVYYCpCOkjn4py/g3euEGys7F36eF4SwI1TXoPYvLYVp4N2HcocokU
43q7xTUs4G1t+qjt0CN3wC5x+VlfGibeLBgia2sa6XQ5og9lcOx9kPZ1rh9MHNupQAyGu0OKtaOi
9RmgQEO/PUBKUmSL3MomDv5ry2bs1otYnkrt8DIaTkbYsuCvWd3TeMiAu69NSqVPvAUqnilDgsZj
8jOzgGcT3PcCCD85R7EFu0YRskBedGFxzxqH6TibZQ9fv3viWfI7QybOSCyTGp26AzAGjySRk/De
JDfiBbqyJvCo3GglA40BdszNU7lD3tIUIdTQaF7Tfbdurg4okwrshtlYDI0XhlpW5Up4y8x9C03t
Sn7iZDrIO7BfTYqF4voFE7o71sPmzhrgIPm1e/FLC2arljB73+Cusu7XgS6qWj35fKHWWDQbKyBv
Yi5RunrNFhIhxLuVTpEuG5vzbwComfTJB6qHuVRPTsbXd5YaqNciboxEetIrPdpBOLHbsMXWlvXw
JtczJ3p24ujUEn1cAC15pigRbovq/YWvv9k6t5WRnSSj1/7G8x89633g/EDfzUmshOwGCgdsRz9T
2ckYeQi3Ln3DKC6nUAw8JrP1NMC3BO47PUP0BGYLfb+lU8vxyHq7YhR1vhFoZ07pWY6Nw1P6TMFB
lmkwSVbMxLerrX7dKuM1NPksmUkBPw0Lz37nrEtTqgNb9xXHAkutgMub4Sn6VbKdZfXre1HvKTsu
bvy0v7kuiS9/mTjh/g0SUiCDudU+2uJh182FVFRPLjaAa6+xthaHpYJQnVRbaRP5xxo93c32jq7X
7AhoFnfF3F5gUEV/y3v5bqL9dERnSsvghDKwGah/wZGl8AXVvVrjIhACKcU4ZECEaC5mYq648wpm
Bmm6dx/YZJvN+su6xqnOxxm5DFRDKy5TNHw2DbUUxjOdg0fZR/vfG2ZlSRR2XrX6l+STysvHP5Yg
qLUyUGzFE2Va/IFiR5L8I07jbbvVw4HY3AfOXPWmV0ItfxNZOrepN71FTREJKbbEHxfxhvy+B4iU
/UYq4wUlnExqinVX9X9jqOXiGT+t98Dbpc1m9sxVJ9B6xqMb0N8wpQX3lvlRsfpiwhfLSlnb0fbZ
HeyrHfkZCCxThqUPef3fy5tWxXzeNuj/0sHClsMHXZv2R5Lg6jodxAbeDYYrdqkdU6VD+uJKVJKn
TJsVXeW0XVAFhxkfhijpozIWjtkQN3iHkwaIonyi/DAbhY+NW7HhPjsiUq0F/ehCbptHeInXrlsI
plBE+k47Vl0hQTR/G5WaZCxnFo0iolJ/LQ/+TB6UGKfJY3MVOiGjqf40Ddkl1GZHDR4CzinY0bTx
Y1lCMHyhMXe9233KGcTJGEge4qys5cjRaLcw1tNJ/EwhtPwD6ABVPy8kbZKJ9fgFhyQHb/YGO0jz
zjH43iDYTM0QnFlKDuLV4siBy3ovFf96HBQ2HvK1ZF1BiV6BpKUoD5Cb5yRn/m/PPqbXsRUsYB/H
4mFDpdPZm5j6n4o6bnx20iQuVTd1erHlcOm/csAQ22+OGIpRG6eRkzHZ9iMSoPWj5SMHjlz3HtKy
u8h/dZz8S9vAXfNZ2faFB02yio6tsA2I/KoflWl10n9GNXLoVxHR+R4rxWqPLmBs3fZn999KF+P2
hBniFfKJmYxSHFxJ71Ao9Ond8Z648e1td22nRLVnWNYPm8bmGuPizTg/fOAQifh58MkTH2CNgd0y
b4QVQDN90CKF+dC6v+4MmAROkx746S6Iaq1RpxXnX3Qm9YGCE37rHfO/m1tg+ydODH6O2rJW5lRV
UhYk3ETCVKG8n/+WVxc3FfkOMNZdLoFEVnPMNDUSlerOy6f17J1Q0UegJG32LYwt/sfbtfRIyuwn
QsOK+6T+/JTG3CJ2eJ3zwvG7M6/N+XdkOb8FK8igmQC8L1yzFN7GZAcp7sLcjAYqOdXk50d/UsXL
WjAlksY9Ys/RJlgpiAshQ83X/D0N2UbUXDlz+SCYqXqW3YfM8FC5M45PWhzZDqY4fa0x4t6DB5qg
qNe4SsLCpGNqV3Cw29p52Q6fNWENQh9YVOgUNc+nDcDoWbIg0yYm5g9qjpIjEZCakRI/7dRCyeeb
FyYry1tk0U0yRwSItT0afz/QWeOHoDlUvEr1q3Ir6Q8TAvt/sIsSbi/8d58SA+3mu+MzC6LpbTrE
h4fRJpuhHMhQO++WAiSNQPSPN0R/dCJIwj+2UyJa7tZX61OEfKhax5IWv5XG3Trh2R48rFtCJUfc
uvaKyOdD1IHk9fgbL09mWoXDw/C0TzHo+7hZu+OawE2LVB4xBphy+wRlzan6Uyh1rvXsi1JEk25+
QGfbCF5tUoaZs45ei8tuhU3EQ6T7NFXVHftzjSfY0Bo1PhOS7uRxDBG2f7orfgg8Oy48uLXEuQXb
JDhNb9StcOp78cJ0Oz4UcwaOf7GxFoqUQ13tgspsFYZzxt1HC8fvIL5c+dI9o9UvTlOPgblXvf/p
ggeRF2scldSPjSygWQdjrJLhH3m03LHKnrRxbGCgw7COxByDVKIQ5UPpgB4YLnREZmVxesfS2S0R
iSY2f5IExZ9RGU6AkbxQohzXx3qChAL4EghyzBwHOAOcGzidXpQL3cIyO2ksSV60Ue3mO4DDo69U
UkCRwIz6HDhUVPXUsRcF63WdDrBRdfXFGLXpdappNYwsZuv4IXxmwelw0nCOpTEQUCQGsKc5Ulj+
ynv3g4hcMXTB8Ge9zee/3AuFLIbICLaXL4W3Av4JMZMj5LRw2eISZ0MHXmoIrhiERwBClYnT9nsN
CI0jRKfxerCEFPVQQ8/C4y9jse7OQI8xaD7PhxZNbDaFt+Vu38R8evKsz5g3gesNbQtyWMMSUsKB
apTWV9rBO2hxdkKXhxrFeAp34bONJmkfY00XqDcS+3w3i9gycA5mNZyiAWVuEO4kUfmz/usMtBd+
rR0subvYBMq+I/SjcXtNf6DqSXTLFyxqeOjMM+msOneRrhhnUojgHSzuRpfZlUUx8pKpU241y4SW
JV0zNl0Wbokpu/2/tlVz6fzb0FlZrw5vLBeTcSqvSTN8G9lvyzw/JVTKvOSyDOai8UFKW23q6rcf
jAajNpQE+mdoTyoEiB0peNzhh9xXTSKATpM/UflmYa6srSh3WJdrNng4k+QV2Gr3zJ4BMvp4hvoA
0Tfc9HzGqe2MgpovX5yE6AHJ22FQTRVs0kqiLYgiRvCis9+A+3QvBugfNSsBzNMzrINbq/WwIA95
aleSJl4QEf6oFiDAqwPuBJeFJN28kzXKwsy22cLa6xkmCiYhmfvIyHLVHX7T+57jRw+eB6k6upUi
W7YjuDugQ/sfq4K0ao2wj0h7VKYInAPvWgQbwzX9ipnUhsoBU5QW2+12V6c2KVD9XuWBshGAh5v2
5iGmzFff7D/S54wybtvl1gE0sZDKk5DGHcBPDoQlqo2KOHioFeDGhMqtRX4JgFsiKrnazQNKKyQL
C9fawBiQY4sV/WPNfa2/nl8+3mBaolKqsSviQiFX2PZ3eIj3heIL7GHzEYqQ51VgtH4G69bok6dm
OJ7hytB4RCXE87d85/LakPDVox2gPq7BPhHsWiZOQ8Pp69SdDI3Ah0x2/fc7xCM8Rljdf9c8y/JR
d5WO8U03mD3PCd9Hdxx4FN94CmQTcxBOAA2Ufb77uxF5DJlSkZ+z8GA2yluoe9bAe2ipy8xBguhk
0BlV+kCJTLD5MkdBnVMGhoifBQosDJEzCfO3FH1AM/YRLvBRcyfQ7kCn8RHz7yDk6Hu8lIAmlvFc
DLTl9wQAyCq1GiqeAwbDBOHN9tbyx4fAY3FPTRkLhoFxQnKvF66J1FFPcjwJS8YeYtza1ErC8/dZ
LMt7ozZCJQ0AsvT6uLVr7zn0DkxeSg5fv2ANIlayM7C0/RAuTpsM8FjFPq7jP+35MEsljEBb7Ojy
3TaO/ZXKhLYDqyMffR7FDO8EZqPMaWE5RlnJxzV+m3ioBhRMZp57+BOw8qDNcKHDtMQcNTB4Jo+i
yY6MYvvxrEhVSzYOA+T+Cp4f6OiJ/79Lx+cAjZBAOkYnf8L4oBKSP1m8H9bx+BD0KO07EErsj8Zj
gJWwUokCQAoZXJz5BoyNz1ol0Bd/MXTrBYVys6iblB+DwpAf/EZp7y6wAWpM5HOa7gniHgwCYrtM
tPbI91YAI4RS78medl5G5H8Ae71dFd+GssQgftiOrN/hEoxT9zdxgfn+xZI6jEBUc5BFgVEm63+V
RhuNWzEDIddm0Ydf+StDkeA/kqQ0hyDYIf9vFlt4qFFX5lV+JubqcGHC3gAcdm7uapYVz4oPZtM1
DaR1MjDbogjFz2noJn2dXvgx0HrL1cpWa1LCIWO9PcW66EGjwHMABOJSaoKRfglpnzx4iaChpOXX
wrbvecDUF2aXhsUWZuZBnVvBIqGwDNO19+PqPfthmTw5WFhrLWvt+7uFhZOLYFtDxSPw5Lb9++FO
fdJBx0AbKHPqqHNdZuDUf5+2x7mnMimusUKzB68F5ETWFGqRj2S/Q2qZVwoYl0rb4SJakPG+sS1l
GRPGgs4QZHrLTgVRckZA6RnKykuy/BGjLeIqFb1xmG409YLfDH9r5SAsjTt7+ehBF+3BEo9m6SU5
wyQ5I+F0l8UrN9U/iKWtxxVMwNaX7SxBTcE/gPa2y78O4Ce2T0ng5DLz/6lqWJk9N35rcTpy1KzU
bl81eVDotv8oczUJVHbnoAAyHpnek/gjg1pIGA9mYjoQq8+wKVAMxVU6e5KbAgJazZfrCOxlNBs9
HFOuLde8JcLFiyjFIsa10LVl0bJrFLJwicrr3rTvMZWdWTRYP3tjrghAbihyoFQ6lJpq5hWzMh06
tmrxc2EI/tNSaPDYeL5DujrSxQRSL3Kb6WHHKvnvGSRLTKXYqnqiUlYwUL4+/DC7gmito8w++j0g
ZByfuk+TOAEM95jWhG2/YE3TL4N3JLX64TaDEqTMGAb0mwuxn8Pm0Sb46fldyrCWb6H379wWleoE
3C2nUMXR83VLKtR2tb2bkg22u84k93dowRPYqvCPGpsQnKnPJUJCN9AhESAG7jKJ/7ihv6rHQcRY
RS7TV4dIvWuWpBWY6XRhQRm+He/J4vbMHAYW0iggOMtTRbnS47+F3pm3zxD65sC6AeDsY3JpCUOg
FtFq3UH2EKxuJHLl8WGS7KW76AhZFhUtq/oflK4He25DpbhNlSJgKk3iy7Mhy41FNDt3D1SxeRUF
dMSF7xKT161iqujZepZmJhJytUkmx38dDbwBDX4vFJNhJAsmGFMC2LoKFxl7kA/J9K//hxq+Tot4
mZweZqYF5D8R9ZmZP34/Z2KsiwMZYZG1wRWizh7Wo6Du1o7d8ua12lYNR2LbOj1WDgs7CJktyzXQ
XUeXGbxay3rBltQHnCng4FzeiLwVAR0V8MDZ88WGjWj3X89SDxfDSy0RKwAGSLJppNeU8XJeoJeM
7Sp+iQw/xds4t4nVGS+DA8A+jzJpzb0OwKFtIh7l2+NjBX305Bv/gZ1q2zQ11UWEb7Dzr0TEL6RE
D6G+Y9vE71JTL9gyoIgKrR3Z5T1DNMVpr0esMkjPjzRDtiGF8c31cWAjJ6RXKCbo+kgyJKxfRudl
6OtMml8Q3Dj6wo0x7KV+Dz1CzNmjM5yJfeR5qs3sePE0dNY6qxTakpbKrTHaXtUaxmEsC53JAcgI
gNaREIu77Df56VZhdm30UQ6h+zb3VMqzOwpMQJUIxG3+OX0YrGCSs7+lODB5EtlVC1n2un33AA81
Ef8UE4zrojuil1ix2AELoudghBlvciPoD+1AfNw9rJtk1WPpxv5axDeMnLdsm04H/+44QWkDqrjN
bhaKyV12Xy0EmXCz89Qc4Mmbl8WYYbrpJsIKF1rdN4CtWvUBi8QqHq0REj3ltM4n6YAYPx+kQg9r
WF6CxeF7+CTHESzXSz9gChnrkY8ExKGakDMVRPcBhsiz1BTwy+VRqvPvaJuuX1pQVItLPOJU3Ccz
3STSMyffg7TEJiTi4mUV8tOfvosluA8WTxBLthkLglWNUXJxX9klsWutwzqJpsi7X+YTg2tlmg6H
tp7E9UJNW/19udxebKHRizugVgQh3kuI6cySLHQJi4EyJHp22ghwrztqep74A+MVFRRZ6g4fItfy
b+yISjj7vO3ZW0jFWich3qR/vVXZWnQoHnztmb/37IG6T/a+CjfJkayLRpzgVijwcs3AR1A4t1kL
W1BFHs6LJ9ObnMxXb4xH5aBiClOI02epC9qAlsN0vQEioFGWg2qNQyxawEc5xG6LbzvYXVqY7WRb
ee0XQE05+lEZJiyL4uneQxAS8B4SUSygY9F6a8f4ekzzMyCMT+w4tkQQEyyylyZ39InBB40DmhDx
kqit7kcAKtWn0iSVbl1XZoikrjglZ8N2FWfSRUMKyhHKtm9rBMCItIVXsQo9BElf4c4/vD2IGVC6
wamUB5VPkjGtKyGWsdlySxU87bhEwg75rsifblKyc7h0v5ke/blWF9GxBdwrXRv1xRj/JEvngpI5
xZeg7UJqQ/nll+ojWg2aIqjTu9n7iG7QS/jwSsnO2Z6vKrbktbjW6mHGT2PwY3Vy9sJpIZPTfkm6
9Tl/7MYHN3ssVGi7OHWezSUtv3TgSf3yzAG2mxsacScXTQvoW2XkLjn0WFsOEQAzyiQK5CsGYp0R
/PWMK9+sZhy3fZhKoLr4Ux1b1EFK8IheaDEOcUUcVpDTLbt1lO7clPZno2xUQoj1+RA8uUi++nSn
Wug+fKhmDQAe/IIN2WjJw9QTtDSXTBiRY9ajg3ZHkTeisIt9/kxMpLPkpAMV9sUbrGgnpmpoyVGw
J8sSkNqOwxzmoR98GqEaGJ7uv4mFWM3flwjJEhD7etMho8Gj+ER2BsQyHNeIQrQvkOU4mJ6vrKZN
naFCKi5fhBl32wWGpIqeX1uAaFMKeo3s3B8r9GMTAkhgMv/9OzOVxBjnyO88FilN7GHlBBXpwqQU
v7udxZXecV3dVxnfmr9STZy5sJJkS7aQbuRSYnJt6qb2yvXqSU5P8+5n4Au4/mDbDXj/91TpM4zw
NCeovX16Y67w+D2VWxmWCQjXAqFYM0p9hV7fHUixfQTPxM6kanNYRvdnsF2sAd3uiVYn8EgyisDZ
laVX0upzRcz1vbdK7y4Sb/ZbymWLaz5DzocHzvRKSgsRX63zRQTxiiXKelmsqJcOagv0rEZKaL8f
8ahf/bqFMw1/EINfFvoaNGd+iSRnyK4ZyxCo5TYi7hVQQPGaRpOsUHTs9jvjYqZ6lB2R2+fcEF6o
qhY5IrMGRf13evScMztph2uETF+22kRh4PPLN90UpNepLbo1TAvZEBbIvPeuU0pWrapCU3N84XNS
AEepspoSvjjwBMllqGvma8Pvp0iUgVaAciE9KeNwWyqt+19ZJt3+UTXL2qO1gnIj+Ga2ZAFxzpVQ
EjsA03i4PdUqJ3XQykFjDoMMMcLV55GaHn7hVVH15zWIWHeIbBNowVNlVDJDWHzNWD9Y0h9NOTzT
kXieyVie5Oc+lvU2Oaw2V3l+v6s3a1mmG5yUm/PjPhNJxvG5p+zZ/SJonNNuhgjiGNuvZCS+VCN8
3HmTFWFuY4gCKrdHIl5b8glhxIbXeYK7IppC7NhukkzHr9xpxh9yFfS6qTTzcFnhtTAmPO5y2RVR
YHtKgvDWNqRaqoHp5o20/LdbaVs3a6ZdPnl31+9GMUafqm/C8jc4CoNEPGiRgmPwRc1rEuyiQ9Dg
WRA1EeCjkEH3x2ftvJNLjwvSvNi7dqOp0osMw5dHqoE9zgWovxkUSP/XX/vuSrCbMMjA7qSb6k06
MecfN7rM+UOIvXH9oOE2h5OpVEqbU8WHqZP0DgPwrhoAdeRPzZNDCplnH+bct0Ga/fvwwTlyW+oy
BbbDXumh8RArvdo7X6zCY0GbILgnNPBdAy9yY3AUs5RW9cmyLUzlnjf6SrAgym+So98GuBEndC3o
WAA53+l5olF5IV8p003+6cxBfPsh9GD3ZLDqqS3fqRig0ZzoUP7Pox6Hug9CNvANWHhYj4T5ikPu
jbOq9neELWyfu9Znh/beSBcgDpj8aVDv/OumHvKbifS9IqkJmt0B41M+d4LRCaDtO/LIfdTzWPYz
YSN59ejvCwoyR5ezKqMhKLmCqvsQqGzGLPYOSomUhhqEkjBHE9lGWtxt5JW5McW7HzGlY/TMbk3q
/1+8wsDSs0rYR+BMldMj/zmPf3e6uvny1mlBvV1rSUcXzx3zTtdsiy9E42AV4+K0En6DbksZvkBy
ARuSD+52l5Z/VR7YaeD8PAr34YLgMMdoTJA0FA7V79LeH9ZpMZCyn2Gt4Wo43x/W9mqICY8ZFDPa
RpB+w/RBTQyNy3KttYo/vKoFF+apsogspEYEiE9ropaHyi08t1Zik6ojs9qSzBXg7FF1t2HGjOqR
fkfEceijIBcofzSpmiX+fA141q7gOD2Mj+A2zPIdm2xppiXTzmO489FShUaNKorvPuf7/WO9fzrJ
O7CzrhIGHvdQVS4H17FP40LBcsiY4Yq+EOxjgzK9ehJmByTu6/9+33m2kIDZT6yMdTRcQ9s3AoUk
AGPzj6z1VLg/NvXmUZcfprWm3r5mURw5u4fYOvzcEc5tpsngUk6hN0xC9n8tKp3AY3ZYfc3tUOYA
4fKkNRFMO3vY8aURYRcZBXOPzUIWuvfO4l8Qq9z4qC/5dKNYg5/cLGh2rZMN2P2a3ZoAfjAknV4r
2g+VWg5w9V4d0PrlshjNVCYb5m9DpikCcWADXiJzz/JXdS/A9rxQrUv27/1harq3JOYmwSuVHhki
O6nCbqwDJNmreS5Du7u+lwISxyfygpPPEHK4y/tkjMmkP4UZpL/S6PxhGk3ja3F63PfRz+p18SYm
PwduHj5cPbrkP0OYhqORkGNJY1qpflbwhwBHhlPrVPbv6CCfhwrrGCMM84ZDSJGbSyRsZWZpGHNs
0hSJz/RWKjR4VTqeIDw1O/wkWlpCT6U+0NEeXiifSBVQsZxYKnfLh0Rdd49aTKkuYyv7RSOEAcv5
oYx3cvjlhRHQW6/8UkUVMYdQsN+aq9u2k2pWoIYQqbBYQMp3m8sMwmibebajvEC9NP2EhqEnLBTI
q9v6Nrh+h1erqjvNppX5fDjgtQ5s3FBezqZz//153l4Gdr7t9ECMujO5V8zcQXbqVCqx8PV0y8X7
CdotB05aJv1YqSL04w1YzVTS/UZCBuZSEUYB/B4rlDAeMoX8Wkm1EUzoz2coYEVr2SR+Gw2O2KG+
5pj9s6GvyD17BOUrikcJP1VmYUga+fnzuEwNOgWjax/rGzngpTi0qyFriQ3bnbIQhXACTwFxz2kf
gUKKH0fHjlx/QLBPkVvujz6lWy5Ig61/LHvypthhQ+SCOXhxspoLh81Pcb6F9N0v+26KsvM8ABDO
VNfE0Gv7m0hWxkSlB27AkWSfTgyOjKIgN5gmJvsdm2E9Rk9b7RtSoVVqSYMqMvcsAwLayfFpRNwE
YTLqfz/nZFlcNPI4kz7wE8JAVwAdkBFx7X45LQRdUT1BaqF7Uhh/8nWYkfvqd2b2OtxfAef3ITAT
UWF9NGIMVEPSd8nNuWMfTNSQ8oDD+Dg9d0iaXrwdntxdcGowyAYOrZlzGpZNnGO6Em1sdhWT4LSU
ZW50+0W9UtiT0f9+z73NHt2zVR3hIL2VwXVUl7kjFJtPQKoXm2olmz8HqycMFuDsglBNPvbYItZP
38lqzga/lKDuzH9o3/4CXKPKATobeYWV0WSvW2RXD4L2S7m28rwpo3SCPkIxP47fhHI5vjb6gCTr
1jYzrrT709k/W/bVN7u9pB7NaBidXvig77jn6G6JR9SRXyQj2/oU0NpiTBzqyu8u1T12GvS0wiIb
t48bQWliCWKPkZLw9L4DcazHap9v50FE79EvNoLVCuuWcL62UJfTocsCq48D297UeFRG2q6P+mjR
W+aE5f60cfebUDpe6a1kvgEcynUTja7cU0lqM6eo6RvawNTZuPwcrenFUSdiJu7qPEUeom2oG3ky
cWJhQzHCFwNQniqnkyNiLx6kacnmc1nce9xqO3wmS9nA0p/6Nb1EZzaTycMFhnr1UKDLx/DaHIOn
7G9WOQEMbLZdPofqQQTOMzvk60iCJJNQZiF43BLmcrG47umYRyUZAf1r6JGkPK4AX9u4KPRxO3kG
7zC6CIsWyJJgZ4hWB5bVj4PX6dsfpQHWp5d7vCLqPS9vf7XMx5UYSRv4Nd3tDbDVqvK0OwywjXoR
f3qCcX/Y39WObSkZOq3pNSCjAa8cpIeNYGcGFxEMUX/BoBg49W7NcgDuH8MQl/j813PJoEUhyu/m
VC/NSdtnEr8mtB+b8+sgTevYGfBYhLbAPGyuM5R9wb9/OaWXK20YycRhNStv97ZfrcADzlK6sj1Y
nLPmaQLOVDt8YkJ9Yeq9FnFt0DSH6PMOF/PefUo+pZLDrs1qrkQcT+2A9q0BSeSXfvt7L4x3AmW8
YReQ5H11Cl1QarrL1KxuA2CCk93jGdjPtcdAj3sJearMOlsKMVnJLAVvBlZQoLG6Po+QunWxkXGf
GtbTVFCfMUHX7m0hTTOCRCmDz3E/oVWme/mrnhF/jqovsHlw7ysyt2sy6i3noGvaSRyerdYHTDXN
z2ovUS2sM4EbFCyb6xf0Ywfd2mwC1sSOFJhG7bVcyoBd7/A1nGJKPv5Tb4PjHe4Yad0oIMDgwTfL
oAQxlidpRJjVLD7Gtc6UK6vImBN9Q8E4faF9YzM7Q3h69mHk7LFHeVdf3vFB6fQ49QQmn1BOTLZN
KlbuzljtfUrPRPkPkfCv9E28/+kdijcyhRbURZGCa5SYinQMpg7YiiI9mY+5QVVa6kODCs1M/zLR
zRSkm5Tfffroc3wKaI5ey3A07qArhyYLsmBCMlvRaa5SNHZOKv0BZancxvNcIi8Be34VtDt4Kpko
kCxJ/GTjNLSs2JS6JtkbWs51p+815hqJtOfg+f6RDHUdaYSxU5kTQIKdf0FWW8m+QFvYFHY7uDom
sIx2FY5wDB4vVp1s/AtwgHfuwyqKVD/ovXN773NoX6Jes8OG41G+6itKbKRb3WJQBzL6YwFdF1Wz
CnhZ4O7Si+BVY4yawOpIs25r3k5ZhjNhGGCSlroKeBM91s967d1nwarrO5aFG/UoWLR6FNaeJnxh
9naIBEInQTiHoW/rBYQkFmpmKt447VPkTozz5b3NeRwrEbMthtAv51E7i43svIiiGugkZMMlMcka
0/vWr6pvgBya+pXY6l7duQo2FaLzXUnvxOl+JJCuxv3bqUsATZ0VJ1XcWOzxQVUXhqw0WHrnN4o8
iK06RyjYkQxhcf39EUXdIdVmEKb/RTk1Yf14M8D+8MTCMpDmTAF5T13q/Y4HVLzFwcKcn7cmSJx+
SGXJPP4hnPmPmuFjwEtPKCiM9KDRoIdsrpm50+VZ/VBPkH3EbtG5YT3igT/0lgD8GEDGMMSS0FQs
k5WEAQNwmmEfnEyFrnJYgqJzB9TGku3kOtwJc3ppj+LP+2Q1cGtboC+LevfrQ6NLwe3YdOGofbPA
Z8MYIUA1By+lvMRfHDvpMuMnOw6ZLtNgnBxGqvYQ8BCUTvdjgC0RBhmJjMB1I2q4bOtEGMBw944M
Va1vTD0yhrte0LqzwKJgYsOi9Z/KTTk+YmbJxzU0UhuN4/P5VeWqGK6THdeYQR+KA/IWIXc8Iw51
HGl1sAcH+NEGgBQiUI8UV+Y7Vcxz0dEGO8trfYGLVcBZFHpy+kp+u6/Dmjf5G/m/rq1QjBWC9BBe
4I1lY1nbs9siK7AvkDpUZkFuZTUfkgfIERxiM/YHhS3B65hTsXKNSe4+jP4u9wadakNx/uuZsNoE
xcP5LbNXd6GgoNffWGJkkfyJ+INkqLf84Usfj3UcaDrE2P67P6yjO2GDtq3VniYCmLb1FGyveND5
DgfOTpEjhTsp/0TxbrzHWqOmO/16m3DEMnDM8duWtxH8cOBke7um44tiflQfnh3mK0umGgNLw8fS
h4Dx1T9q6Ik+97/3i5BGh+t67yn7U6beQhPtpyAfOmNLlH2j0iBP96WEaGDzl55AMB9v2nql/QQ3
uWEzzLHhZQvQDUf5QP6uc4PR4eobTs5dHHGMUEHZK1VXYZ1KTvmml8oarZrZTLRxnbSlxQQUXwEG
sUUyu0Hr9OhGvnt2/ll28OxqfeLXv7ATkfVAZt7YTTbc3HW6jOGKNhB/PPy5ftFu0P+FghU7RIsu
AuAHWI6GErrNI88/aPHCGfsTmwNX1/eZzEexQZEwsK0qzUPnhw9XBbQQj5k9ytnbb5zAgxXsc6Et
GlEuqA5lJKXqMLPs47WJVDkE5xyvf1/wExELRlrs+7F54KYfiY/IbPf6BxR95BdTcBx0Xts4iFXr
zQeXNgrixyyzaXIerge8YcfWfiTeBMS4Jpg9il+8z/h6E+fT1qcCQkb0/5DVTXzGKdPM2oO/b6Rf
584wL/1SSaKYCNwdK22r9OuWjiXMIH+uXIWFoEFHXerHv55X+PP5WjjKcqpb4wqn/KwOAQnbL9B+
gyrJdkeAUfKhGgN9T9NTWKmGWZGDchNlbKkHnFW0yRmbkDA3RJUB5SvXtVPykHl+vnPH8kItYxsB
JdmXxdl98lfgHk2Fufr342l+Efh4VedLyz172MjSZ6/54JWvplDvALpXtCeTnYjynTRkHlG2dxAN
LWYlOqKy2lgyywUFEi/NmoDnIh6WRh7MWYtmhohDsc/HQSfdeX43uAHoUTi0IZulCqbdGk+XZzxG
IBO3Qh81kQktjkFAKpbCg4+vpIK3DbNNsb+IUCIHVuQSkLJUv/lz91oSbw5baeJJRR8I7CroNAs7
Drvf+TH9mkHB4zIdZXHpxxepatmSW8YE4l07oS67Nv54vQRblSo2kyUq+OUwUgULykHofIm5oNyb
2zSOrtlAbfLOVV4o8gboEko1gSk32eaYAP2KjgYb2RAAMmSpmB1FpojuEhMQjDWiHh0Dg4lSBa+Y
n3MqeQbScT+FTgGHSCH+UhdlXN97DBkvT6QjwpJUN1iYNpYkbpTZHnWG1FENb8EH8cj6HpJRLAIy
g4x2EFsVMoATiJnynzN07CeIsB3CpJAfXWGgRHSXCd/WhVXKiubLYvGcs9y78S8P3O+Qja/sg3Uo
pCK5S5oHj2dFhGr7SeUu9L8SpJD6OxIhG7tk3KR+F5kzEjou7Yq7un8LFmJAsOdby5w2/QYqEtvM
0uWnt0AStzluh1CPIt1X9vhU0fN6YdxRZ3SM41CivUpOFYM0dKx2OTpCT9TugPcxmj9bYeXeFWLI
icCg8z8zmhRaSondSUPfUdtXhcREUHlppH9II/bgvBLCFksZlpSnZc/RD5RQ98m2goTVv/yiEGfR
iOFe2I0zhBKWlgGKrUoSCL4kvxGLlLQ/foh/TLtQZCJTm3u2sSRwsVXgVitpJ+z0FLvv9KdNlvn5
ygha8wtLR94vpDaA/RFol5t9j9xX5p3BhDeGy+MYr5LfKlGJQ2QArpnfNIjUZOOCTPPXWJaCzYh/
6vtBm1hSrSccfGPgGcFHZ76t1hwItxl1dMu0pQjBkShQHbRKG89nGKObgEJ9B1i9GbcS9QgjgFKg
jW1/hxxphfQCbF0UD6ZhjGQy2M2Nt0QxhgjHVYrN5CpmUvCt6qNGAWAhqHSqu1iiyE3jj7232g9W
KqjfXlJjE5bR4DiQRemdJduxWBqoDrzNxeL9XigHog4heyne3QmkVzkVGX3VKh5ULRCKij1AzB8x
IXRdEcEgcdlFW9NCdsQonpN1+D6Koj902XPHlNF8yAy3LF+tlrhBUZbji2BeSZvWpIaBd9YJuQBX
wVcUdq1ISL+3D3U3b+4v88micTCmnUdxr4vW9Qm0xVUyxB0GFCVZJJbKil8IwBXmg0hHP8pwBbuA
Wp7wLb9YhcZwBmzZhi23EBUMUbsnIDqYzUEzuWsuCI5pBYsOApf/pkGacc2DdIFQ7oGwMPD8ZcKq
csKHFo/jcDJRm3lAnHulDG2qERzAFdHWUmgstRj09hDChFZWsL0x2boaiwR4+tnbP0fA4kWTGV9z
g8sOhJkD3DnMLJaVyCj5bjOYG/tlCooCXCU+euas/e8Clmw6ElAFtZSFyPMAuSZxcjGMk/T3HpdA
fI4TOvBkVP/7MpkQcKg0ZKHYn+T0TWckV6Gsl9B0mnjaA67aJmRhQlQUWlK0vnRk8PEF6FAMLxIg
0fVCIGpQfQd7oSkK4ZFh7dZKfhlEiU6TxnLxdxDddfTG9eUWS+RCMODcxm97P02i3qr8/DLjvmL1
W+b73Qi7Y9rqW140lZwZBFRO1kChOqBq8/MQAS/UTEqfbJ1/cLqeNkFmsghHwNwi7/G1VLvgLhYF
w4owD9WudHxVVievlJDjCBWclCQPcp8kzlsCZTRYzB/JTAxX8u5HgfYiNeuHpLMAKvczeaq/5pmF
wHr2rb7KkXsAtcWogv684jkgnzdBGQKKJGHUUZGb70/0sML1NVi5wup1GQOg6q0H6bNSLZPKmrPS
W8XC7W99lk7N15X1ZP4AqH6vTWIT8TSFx28wpALN8+rsdaAAIK/Iipg4Hv0AVPrbfxKaOx+ugrHJ
XGyIBBk2Qde+IOuNnRed7uQkHEZ1k37c9hMp4cIC34nHTX/x3Bf8iqdUbfpMi8Q0jFMrPJGzsEZT
4HlEvQOaF+FJo7H73hbcERfiYihmfN3Vz8/L/HShker5F1tUdWj0QxLPypAZJDukX3+F66I4kesS
9dU0MU4M2rZrtHMZzn0y+5SeK0Y4kaYLIjTD7KAMC4axA3HsY/jNyLNmWdeMx7pFz5gloPgRzGNo
NpAm4NuBDW7yIJxyqS7PNbTipDvKEw5lH3int+jNRMQm9qqUvJxLmHTO7nR7zufWczHKNa5i9lxs
XOLqDYfOCk3vFnLaTEzFixtVDC7Py2WaE73cf79YUEwPYYDd0d6TtBvDx1PBwQC6NaE41It+4SiS
NMK+wUGuUEoznIG5MlPYTxtdutpOKcHpzPUdiTwAguSOwnnBh4TTLp/wUouKqF5+RcQ56n9Op3az
0rNGmloSQOGC1j7nqHbYHockRncEI5T5IV8PvGZAmvFN6ml1h8amg3qmAiucnsKyMaRTIS56P+Yg
D02lO3RwIvyoconGBtBRfB5xqQeAbKTyt7H7x2HidPt+qXQiw6QBbmDVZGeRxEDAA0k9/e0nULeL
2Z/wGLgMV2pvrwqHfWMqPO4o8HBY2BgRlVwJQcNGAAzzOKDm+F6UreTrd9HX+o+SakgvR2Df/F5N
B5+r08xs2f8PEsMWLVpZKuTfwfeQnQ3R6j+r45QUpZ8Nn3ucFCO/qoht7+rPjPGM8jcKQ5HK5HuM
jj9ryeLJP3kK9COL4UROrdXXa5YatqLrmcX9Vd9ze51M4d4q8BmE+QcJU275xNsU3O7bvJy+qY/6
GxA591irffDBXHpwMb22q23jmaKXwGhjIoqCVSIHhUb4HKrZe2rdGKpeEZKo20d8xVDqn6+RjUxb
8HJb2pw+uMbjf3N5s8rG9L+EWdO626qp/vi0/RlaclkcuFANzPICH2hn7qPFmzcbz+CFnTK451Et
mMUQ0tNWv6Bvpu1km+GT2jNOEmGyDEupzk5eqaB+zVxCPCY+HH60uL4+Za/B/4FFnXWIyizbk4Yg
h5l5lwGHA1sWVwSlHhzGg1lYxz3dvMf+dyEDnW/NNomw30Qxcw98tlq+4YNP8hKppBE+riJWjpY9
+l+S57fJH2FQuv/eHX/RnI6v/O8YbSrmjxy1+xxWMT3Rmc3v4gWfQUL1wJrf1Uqytgh8o9qoDb4o
lctN3HKrJxVaCCgCa16DzXTHPnoxbMN3ciYdT6b4eVXPpFRV/LWLQCXF1AjblD//MrFProdbYeHH
NKrNCNRLCV7ZQ5pGJd0QbO9RkXJacyEI6jnDOQcUmCLpsgjS6+GQ5UyS21L5RhYWlqBciZjk4+SE
jA16fUr/1nobAmffbVnV/RoC9vyfsWyPFTpWT25HAfFvW7tr957LdTwCoggOhZr9IMi0Q79gERT8
jH+/SmVKsJCcIaI/sv19QR19Gt+Tutnmn8X3AUhHddGuyne+OK+537nZN23NoMSkm7bMaxqFE0Br
tBk5SBrd7yO48/A42Y9DgBPAjuOmoQhDVEt64yHzhQG8/+K2MvMOE+/34wC9qVWuZxsw96F9XNFP
wC9aJ9/qKFpieFXKtbY2AlQYw3kf4YFBbxXr0NVlZAsYnyzPdetAaSHNsgBokmx2ZI3ACEpVV+0H
mFBvUdooh8Q8qLg7S59SQ/CRqcMxth4e1fEKitZsBvHsKxtcAMvM+HRt5IDISAn/V2AID71gvJ1D
Hh3K9Kscf+0TAm+3b2yKwAACqkg+rtG5MJ0RTlth2PWcLKtI4mvoGluftTT5yran0cMm73rZJBpV
IqXwQAfajX47HpCLiXb8+JH+OTIEu/6oSC2Qb/h6N0fE8kWI9Jeue7gBmA/uArbKcuzZXxc4Ad0K
udnW0fPRmVUJMq1SPx09fsV+gyHFfbjHyznMOZDezN2DwxULvB5LpuOKXhhf338MdPfOwPqjWBVX
1nHUwnEAHI8PnkSPUFVDgzx4Gf5Dp20vvfXRvvS6kJGS8vPsN1yilm6XxTeUVn5kozDmCB3vgVTG
nuYUPZOeXyF4b8oPrIgqLrd4pyU7HKHPJsL3Ht43JA/0liG8gL2qDjjKEaXM7yGEOJbj4JIdCbgt
iN+iOZCkrcE5tWm/P01/B51busYs8h5kjl2vM8wIIu8WzWEBVMtQnjPWnkXcAuxc8FHNndLxDJ5X
OWuAjDNEAn70+h0Z3t68D3f3LnjimCtp/xeDLPo9p0/Va5JzSlWkxO0Zjfo4FiHNcOKdfJWfnERV
UQOl/noSwMZOy+0zZaXP08nmXy2bDUAwXgNW7OxAFuAoU8osDhOG4utKM7PVxoUR/p2qhCKhFpX0
uT+Gezs4IzZdJWHiT3IJspwl3PRqfM80iMTJARrnxNLdDuLXE9QLxgbOzHMXcpwd1o2jbH+uBV+L
afnrBvk5Jw2qvBWmK+mF4BltV2CZB6oAed2mDF9EOcpMDmsIxhUmZ5OPm2MrCc2VEz120ZVlQFvt
M4+uLs65Te8I0TM16Juf8nYW/emtujs6OeF6jUTYQbT2ySB3RPPq9zllcEbDvdy21S9SzO5GMnTA
Gs1SCDsQ574vE9hw88AoUNa671lYw8GLIdPI24BnIIxJ6a01xJ4pIGCdtSl8S+O9hhPiO8g4cXU3
ngXyJXXbmXLsXGdC0fgCG5uosoU/tiO2X67saBfQsWx8OrwGT0BDQbDgMJIWI4O6mBfqr3RtLGSO
vDQjaf1FmND8iUL4UOHg27WCYkwXskooZ9Wp8Q2GVN0m1ZzsP7mp8zmfe0A6kmLCA2IyaT251lJU
sDiBrqXxwFRcU0CtprGfV0Kc7Ias0nViAsuRJWf3OwqAB9JCOD8rg5ntZFoh9WYjH0Ug+8kAwiUx
f0s+WUdHwxzxp4teSjAGBKeGwm3ib3dpfrd2Fu4lafrVnByjvOXvsthJeS8ArnnMX9e7x+/y7dI0
6mZQ4Gt2t9/r8U2J/bGaCFxaPtG/eHfh70yb/SBfuADcK1GVSTM4e8ZZWPPocItveR+kLGbRrijC
Pv7bCZc3telhFgwoO3LUK+yzpmtbRmXeOUTG12CIMNfrRc5uQWj5dVDud22wYkmERjmYeJ/ibYwi
7+CmO8zEBuHlun5fMK7aSzxKN0FFGqHhXsRmqmfeZa6LWjkzvM5PSQvovH55fPDMYCB21i13bbjT
AS1BJQfX0pFyAzDRI59V2goNjIa60O8vzQtHSoPGtatf0vmE9rwXNIGAKYcADIVXCKIYOx+80K7d
MZsMfEox5jSh1EL7S5rgMHxxYCcZhly5MtokDjfoGtZjEuz2jnBMpS22scgI5esVo9onQwjZPXK6
ypSFzxmU3k6uX/oX9e+egvdOtAo17Cw37uz9IMOF4y9C2pqDx1VmIUkKeadtBoeYILGxnAmb1m2g
mwnYO0KZyZV7MbYDlx+vIqLt6IXUikZzbx+QCNmZVU8w7P04dHbLMihrDTrS13JPeBniKCxSMe0U
b3j4Qi6l+3dnw2NCZ+3t7TM1rAIZZBEa9KMTK7ySwHW4IsnlD5g3iKJRHjigjqr5YUDmkxVSZDxo
mZjaVnemGDAFlr3FP9GgYcfoFco2cLXybVOL0osjvo91J9tfRn6Wjg+qwpU+ctkbNBFkIg7bfROm
ILK3Lx44gyxAYw6e587cTgAW0sEWtloRvNydz82QJnWJPfo4v2nyeGjz6tcBbI+qm3crhAxeJsrl
Ivs7sl+5YyfZtnxJFW3Yi62n/sWpi5OU/tZByrfQIf5TPBzasZbnYe4dsHNDc00fYxmfE9Xkf4MJ
cxDjlMwV+3cIvMrvW8GFjY0TA96wStsRqBJYDRmT8YMNndSd61h2X8941uRR/cVOOF25nDKa8Y45
oM8+FS48IAze1Ky94lYZm6M6gmXH4504eIVX1yiDtPRI5mCYo/XEpXNnLcjNbh8DCXZtuQ1jecFC
aceXHbtvUlcsIM28SPcSajIYl4UkQMX4zULma5iUBP9PLhfVuzGM1lZc2yavpMQXNXRaPQJXRd+7
m9uQGcgMEy5Rvb4widKUoqcxCTnFSLoSiTnjSXB4nj0SywLP/fZkQp4Zvy3q22QUxOciln3xII7d
5biYywuLizH+SP40scrkwTSEIo4DNTqj2nd0y3Mt9vDz7ThJX5XpuPJj5S0FW6sbrFbFuHBpvfoz
BYjC/J0kj3SqVahV+6n/8m/Ww20VZm/EJBHuPnxXp27RjUzniq2qkjZm/EPNL44uSFAbuK9jXvXw
I3zW9KNXdF7S+73waN2+cvJ1H2E0t5DOpA7UH3q/sw0ZS8Uu2OdMBczpg8uG3RAzTLNZ/FmfGXIp
S0bTTMFkHIt070n7sWAoBrfIHqOwmC5zf2tSfN2zKEPfD8GUlALBYq6ZXtUsTJxffhiFi2odK2nD
3lTd/k0xaGwuNl53AykwwuNnO26Um2DeI6Mak+WZf3M5mnXeExtsjiinityzmiQ3u6RTadEG8++/
rHeDmkOHhuLqh2JGSqpLpF00jXL5evkXnrkV0aSyY2TVDPZelaJ1pg8GnNJttckhq4lxWadu9f/o
MrXO27Amot6SGyBWaSWaPodzkW2RfKSLlXfLbEi27rbzcDSJwCoTwSUGtZSuHTqkqXMO0ovaxV1B
ICFKlCh1DQb3lNZ6E8jF4ItxC09HB7sgd3tGgasz72xxaJXloEdzNg/gKUPDAeEb77nnAdl4B2oE
SA/y8viizr5Hqe6tmHedC9jOBHJ1k40CA4y1wkKWh5Tdo5QZUvOC3UxpjHUKU6t4n9Za4nr2iBzB
XniZwASxM0hLfwUgq7p2olax4tqX5dmtdAseEeaI2MWZHjt4ehNIPNXBgWyq5v9YyRG2GKeLya4C
MychO4xdS/UNbHiNG529Z2PJ2M5IjN0uKNptnYGhlcpTcGEFM7umyZe/Nq+QVWa0QGs0/EmUNDwq
nemfca1pwp8EH2rW0oKL8T6dMFGqLaeNmIEishv5AoiNjTzCZa6P6TLHDC3pL9UxAvsYqPaKEo2X
/RlUHqO29PwGBgHoS0b4vbeLmTIEWlNqhd8b36+lJV1JhWdDdDtONGr+m0OEi+6zk42xW6jZ10BG
mMdX4764b9aQzodrVlWPxD2aXOjC69ICUHDAt6I8OXJstcspFfMvCfzHmRjgoLkzb47njmnSb1/V
dNIw1k3p2e/Hsp4nwgVvDYrKclO9cN5LHvaHh/yR8xP+GToUGHXxl3y+Q4mBOQVzh22cWjKVI/Aq
thdpNkFhzcLIhaFeu0fzre+sqmQfnxMJOFQU8ryeqCWiA9dclG9I3te1DX02xWJBDVKf514vjojl
RFfRsEQI/4aa9lCa42S8KbsUYrIaw4tIBS+POUfLuuCpZxqivmXYsCTvkoQSVdQUs5QlWJqBuhNk
++Udc1yrTzj2eKQDbsjpQ0RMqtQBofYMEUKFrbfi5VWQk9wuESlAC/eGE1tLLdRmqs2Y4EcD1bIP
Uq3DvAwSluMSc59JFs4VEh1bQakpGxbzZaU06xJIfHhe8ntrGXWmrTlmAbIRdv6MKc3/iYX/6MZO
qEELPOhnIJYitLJ8BRonqopQ8CA4tFvlLw4UTKLVa1XU+lp8tw4kBla96kDBGirb3RFxDICLZDBP
Oz0DaVl7sO5B1AbV3UoHUFwon3U+qebW1U5dJBjgUJeQEaOjyHXk9S73Xic4gt0XI2eg1jX+vu9V
Fvbngf0hWm8ntjHkG0xix8Uo1a5pIE0bQ4XyByq1fu0Jk9lRSHZcTuiXsryJX+99LEP7YQZzpW/D
NCNZlIX/oL6ZtdSCUTy6cQIfmIx1ejXucPjN9rn8zyvPDPiSgEtFtDA1OpsepG0Io9N99xFT+KQ7
HgelUrYZGvGwhhVxZHvLtiNgePMOgZZpl4iTzBby4yf2XX23M+QDPSjSCtI8+7BN5it5M9PSslKx
cD3OWLQBOujBJY4UQZ+HkmqKykCQm450Xs/Y3ibstZpxnbhid7WSOg+5ofij6ChdOCYenASbP2Uw
n05hswrogSuMvELrs35+iOp8G77+hHIh8S80edMod6ATcWa4et0S8JA5xMrJ96reK+fzN/Fpsr8a
ZKfq6TJc3E4gJrh3nNAPfQlxI9VSxlqQ7I44czjhzOHyl3ASHv6vR2FFajzFwkYe3rtxuUIOtON+
Euar052VO2YeGepgqhbHw2fr7Km44ccfZMXXx0NZDHlz4ng/vtqFKbXIBlbweh4dINhsE4UQyp23
wl8rOCliPRRrfyyIBdkotA8nHwE0kwCIrhHaWj/WTVVi6UgBhxhpndAY8Vo4AiI+H4+sjvZJDRVt
XULiJFk/f/B0DFkrWjYSQHHXpt+WTYY1WAnRA7QFWkAM0G26IPORN54cyxrXhf28iOLJx0aMhsE7
zn4l3+nfpYFa3FWISEMSTSn+ZvXNJi4f5vcmRY5XMD+bWu/8cDW1Is3nGAq7R4b1FUm92eKiaUZN
MLs0NMTkWOcupMDCfIV/A8Afu2Wfm/dzRnTP9v5hBNqO6x7I4cYvM9knFVi65Ok5MoTBADSJX/5Z
1jNU+1vmTOVwjQ8mNTzs751qmVgEt8+XbNx2TZjp9ArUnduLu4Tj7z2xHMkO6fTuwQ0XYGyjBCs1
Bif1Zyrr9vamvL/M9Zt8VFZjrVuyooWZMyGuGspLKXUVb5WJpuVhb3hnEr5y7WHJQAhKjTqhnlxg
CzpO/x0P4u9I0f2AqXeOGpBIaxB6V4htxcj3L4T0vZfGXpuFaVa01KhlEc4iIBsN2a/AlmEsxa+S
ZX+WA4qVnwZrxandcl0b9+abT6R/JbdIczYLYd0k9SNLcQxYh0+8hy9U9CIKG+3wwcV8h/2Y6fUd
7ezTwYX0MFqrc2XNwl2LUsR+Y/FSX6G3ZKRFxYkHNcdRqs/H2qn7dzbo3H9MNCUDKRoYFJram8je
/AL2/LuqgUoPA1pB9hhK4U+njZr7QIfMmE33zqB4618sVZfjSbRqEChSNq070kQM3KY3gmRMnhKF
HhS0OXOp1wlXUTiMlJO6TUZWU6pMSyGavNtBy+uR7TJUGaiY7NDkrCNvu+LiU81MUbRYhrXXYs+v
YGY7bryEyFO5BcTvrzQJLkei0xFzj0v3N7Yhg23Mxd2W7Dd2ow2r/Ij8pW1jqMCZJv9hcCLXDKJq
RVwtD2BZ1GwetDomP0HcDdYV5V8/18l/9Nx0Y2CjWGZNg0Usl/4S5qOrGYffNgC9y3lqhc+dU4vN
+E1QtgjLivX6Np2p47SBVCSVnreYEuB7Xz6Gj4nrrvJtrvlAe3y+RDPHWxRMeMqI6SBR6gFjFccS
K6BJY7a1gubhKrgLV4MSCAH7keEEq5gMI5SnDKjKFxygNAOSZQKEx8+MHW2RQESfbaBLYI3ylAc6
7ZuM/2T/QWEvEqmMXStBu15fbkspC8ydz5TamVwM2vnI5DPs2FosPT3tsdlc9xLkDrTY8T7/er9b
RldoGUjnYuVEJYDj9o2HRyfS3YaV8qjilV97sd+tLiKhf3c8Avsk/1EynlJ9GZdhDDnwoL5s1xuJ
zj6jh8iTiFV4coMyHmQOfCfPkHikB8/SSyyj3zMXWa0lGXVux1q+JIZxqZ2QgTR/OXjpHnEUveZu
rgrfQrPvoOuDjR3Hht62kOVTCkB6s5uuCK2lfms+qhKTi2BV3Do7g+wEOMOTdw1TOYJKFNpOa57c
BKdmJmZTdQOZjCZuSTKVoPgYy4D05R4yGsxcRL47MPI/jw3039CvMK+3yYBzKhSO+Z4HtKRHbndo
r045ngweSnkzmImdsID57FracUC0N1oqJq4AyccwB6zXQg8WPYg35UftNSFVuo/2AJx+6+rSmAPD
OLtn3r3WfXybukobiR1lTh2BtVS6Zkp2hldGQ99vH0p1oSGUpIPI9wz4n7i3NWNJ8AsiS8TqDcf+
k+YzLwn+xWkxcMMMVrtYAx0ydIq0Z7STaAETFj3gCvOND+m/ZeKze8yuw7UgCstP8BWxlWU4mjZi
YvGJoGTtlUO/DiE9gUa/AODMoF9QUOIxacSLwTlB655UGr0wG8gA0snQioxfKRt/nLxZdvkyoBcm
rgU1upF7vWQj1B5stbakvrDAVrO1m6dSYbn0Uay8VxUUk6hgBWjGZ9txgSLCAYHucXJG5E0HF/Ej
wZoZ/ht9Bz0N7Z7ywDTM5ym7WegUN4wix3oPEjSHCHBFwBMTWdptLKLnhHLrUjXs0DBJdXfXGGVU
ZklUbx/j9OZBpyAmbM8KA2krFLa6meZF6FCMee7iuYm5w71NmqXnWo3Me4ys6PtPPPyX5+7UAZSB
G5Gayh76ajXIEGz50ypL57KYAf2Dqn7hgMbi36arvlhVgAPFRtaaj2H1KRpsYPVcS5Ug9dNCC+vu
zwk2CoVgOcL6UyqfguwmkyMNkTFj6yKFV9YtXASCKEyuqKS9xAKfvhimDk33re4sr7SmPBda+XFx
PqCmpUOHyLE7GnqaxQmYTo0m9QFu99Bfka5x+0dnPtlZiMdspL/QFkSJjUP+Y8u802PkOkyh1P1P
mAQMw9kR+tMuBOblGEjf5oeqy9CHhbYqmek02yoFSniSq4XqLj5/9a5/UmDvcNQv9YvlSL2RPJCm
PUEcT+S9M4zr4U3IUUwizlMKpCszKxTzn6mcmz7gdm3++t6WBIPwHY3zStWD1D26xI42ldsLJPTi
YHOwSNptX/RAD/WqNQtKp3ODboBrONarpKKNkxPHbLrNcf7CHosi+BJWY1VFacH7blUxzBI1F4Yw
v+TS8FlrJDGeyZvLNUgddSn4SOPhSAt6k3ViNi0BqAa8l7g24Ywp8St5TfeITKOHo42dSd5cKWiQ
TUEPnDJ7E8KMRGoN/u0d8IHlXj0NCmaJkbjM1+JJoymUvLJ6V4O4PS+9NELVSK83qCWKBPvUgaXV
DkXWZ2jVFiNcJjHyPoO4A8TVzBnEQ1cjkiHDxaHgRZZtnkgpMsuoc5gMzQw8NblTOYlZge4mm6a6
KmH3Ts3ceLAcmaRNdSwji9mRfnvwWU9O4UXVJsKRwCuB2kQkVS9gyVDTcaq/2UDpPA2qLoEPvWjN
Y4bQ4iwN1R6zRPjb/H5YhRihTaQ2SRSSAsUPmEnDwW6QFWaoC/krl9dwekxDYN+57i3scDgj4oPw
XV9chTHz/Y73nVl/WRmBO8eg1MW4uC1eWnIN3NFVBjwPK9bJPpLZTPI4DIGbMp/wy+ttOv/+3ehW
uAsGJTvIzA+yEmilXah75NOBqWslraxOCrn7k4/kwqeq9gC4mMix+TblwIxZd5rDSFvFyR3Lr+Sv
TpXrLav4YboqAviKMqVhs12V/nSI9l4jloIVdXCrBFN2ndhPvoqAo2tG98SsD/dsGkyMVX/HP28L
7rGuZuHPoEufynD+hNfZtMjQ9gbToevLzI3dg62ye0TcWmB5Mnd1zmEQr45TUA72K2V5OTxLbivh
rnrbbOmhJIdBAVKQIxICLDnTpmbkcvAA49YnfGTcQ6qqAQ1XB9Q7gsGZogmzmQzl4qSO9u5Cpn+E
nj6qa4V8X8xcLyW8cRtNEmWbNhZ33uSjOcbCrljMxiZf85QY+KrpzTdwzxMgwQ/J92SBW3Kkzopu
Z7xz8S5FgEDbR5VTOqYsxwXiyJW12n3pWprRM8jdIpI8+x0vq3GD+8Nuj8XtgtdiC9RjExxDavPb
mI/g+vUO2o91n0pKhYoXkr+PexT/T3oqFAwWrTmaYMa2Cpa8D5ToF0LrsJmcGtlCvybUD6ITLtVr
TqXjGZdFP+LRbRSdEadrURk8tWFfIoVZ62jxAAM6XSNPHjU4l85ei8I/pexRoAtahBRl23hJw34C
0XAl2Lv5NtTcvJTRt1oboqQiWE3/flChnkcfCwQlpYU7XF4m/cDkJMkI2c9KEZ6wweAAccwy1Ii2
66JrrvOu8+a5sr7acsVsKf3DHnio6xGhvLR0jkNLTWJZuAY9KQEDM/VMyCl56m5nv+T5j+erD97f
8EeYpRy8sT+51reNxHgjSSXCU4brse3g00Wmb0MrcuktkavfgEeiLdyYj+YcCJ6E14MNY4bqNM8q
1ea2aYzrgk+w/vVONH2Ah88P8b0CHp1QCfsfHw741rnzeeBfIq17pUlE/uSjD3OJCEbuoPb4hZaK
m3dkSBh7uHUo988HV4t1NN1f57WXAMY7kBo2VPnYrixxSDyac9jQSP1tdHCBfKkPmKB+4HEN8LVp
Pdn5WIRpeBIlmjwFm71b2EY6gdnUC6cwyi7rAZ/eitu2H7cXSryCJYxt+/WQ/t8mPwBZz6qqc9lT
/w8g/vqUIA1n0g+DH1dqSFXmJ9eCCUE0h3XuH+/kuVDX5Y3u9Q0fUdz4zK4ZXvhapF5BPYDHzbyP
Inxf4OCHHZyuA2Cv4352Oj/dCm4TIqTHv1n5rerQ7CrzFK6KWuJ+0EOJvJyep7lyKZNJll2oITt4
MbIBzoZUnN7wYIR2yYQ7MUlRdGuqrslX8WkxEO9oZDMhJIzf1ozjDcgvmJObG7hFWQiR1D2F+ulZ
pWBvrOwZQVe6Kt4Yb88vinPAKJUACGVKvfmQM/DLk30nBvH5aArH/+4luHd8+bX0N7NZTFXw/jPd
QgWpJ+6w7Tf0ETlxOooj6Lx+atOPiZiREO0lRBKgSR9C5UVKXrdr/Ri+zTuM6LJCM/zjuO1BHzhO
aWdPbKQ8Lv54lFI5ycSZ269ETeRfhFezed/Jmn9eRFMAe92fXNrKaQyml2a25IKxfI8gLrCfA6fq
zyBPLqZE4mWHFKFKfz0fvBv7r0PKsB5ZRC1oi+mmCeI2hTvykPc/1I+i1y0wVO7f+rWD4ErFosK8
3jX1bSeg6UrUmSVgAyfYseu1c1kwOTNT+gUEK/QV3XBcCFmTWtOsOa2G9G4OWVaJMwkctv6VQmL/
MjpehR1W9+nEMebnG/DbP+bbZ0n1k9oItYvVMajTA1rpzu52VK7EZch7WZpHvd6masnTPrpRuKEX
ocJM/5YQtJOiZW5U3ZJP2BC2JX+zN8ns5M0KJVHJA2ekzGhNr3naSy6i06qnMU3T77zaSwVIgHDW
tbblZvNUvoZGap/G/DchWC5+JoH7PIUh8hRc5DCB112cJ05hrZWVGm6vUQiIZdB3lR8h2MVXN8LQ
7ZKKw7B+PzqEkw+b1MNzFIXo4ByosLatiorkp8az1B1yq3BBSPLxOGOLb0LwfUzlZtKcOfE5k5qG
niA7NT0eqvoVcX6GS2/5mfhwNZd3kIIdaR+6Vu4p17S2hkH+ZLAkvubQ33LnGxLuTNKiqrOBgXq5
c6gzBlxx7rooDPU+WK4Ei2NeHNF+xdXGiyXqXVy9T/gCm+uONWSOrG/JVXAe9WZ/9wYeGgdhlXtm
S4eAP6xviIwNaz+OoFfVM+ZAWr2cGod2hsdpiy7LhPSRQjtLfO3ZXpSQlCyi6TPIqRLiEVnlaFyh
jOPQAUyAG9ZnoGRzs0/as90K+/PCf+x1jRqZ4F5WXZCquMxjV5As05AZYbN1ILGTiL9/zob6QYd0
Oi6VHop8JC+glR/OgoCN/Qc4F3AUs/LY/QZpvag8DeHnLofmhN/1WJ5QJMpEgY5kEpwK0YNfHTI7
Z3SDAGINukohV2lDjnWYjrhhpT08qvQ8FU8PM8h6+K9TL0SQur6OV061zBVmkxFYQ7tixlhzN84n
H7sVcBKsyG7g9LN9kH2VWu9eo+kPfErjxMzrkPAVcDrO1iKEYZZVBIPzJyfYNKK7TiRATX2IV3Fh
GFea784FZs4678U+5munKlHQRJpzfMtgiNQBF/NXSIRvmq1Ia/nvm3hAPwNeMNW2k6fxkjnQeCJt
H0flaacL2VHZU8EWr8ezB6ewuqGwsdERzCHohHqVpg5YhkKxlFdkydNwPOkFgS3ijbregJazyKRS
Vs1W6gOvAsfhcQ7GFP9gUVCmlegGCh3r4rit0/p+StbLKrkdefEUsA/Z42tVyPtTgpNeC2fuDwvI
MekyALRpMEaq3Ze1ywBC1k9jam1HeEwjvfsk6IXEeFXbOsrDyO8GKCf7d2TZyNvtgebQsGrq9Gx7
/FqVqgHlS6WqJ2w6I7y5VMYJjI85DoS9p9m3W57yxldOkyP0ALV+/MDAWNC72GEPpPCN18enzhcB
HJSa4tQrUxkoW1GP2B7ZfLJD1AnvtJlDpUnvjQP96pnxrQdjGT6jVTAPJW8jwk/mNKJPk+6wd9+C
JKnYMY6kKoyImBmW8Ji9TqDG17hCXLCF9vttjtanHQID+mZ+mKuylC7Reh1FX7UymtmJNvT/5mDf
6VLDvgO0LsYqZZgnlD5Y70UosB2KMXs4XQZmw6yl/ghqXC/BZMBVBsVHvT3KnbQGYhg05RIgRYAh
8XSBzibAp2Te46wY4zkXFgTC/KSK+X4rSSbjsWUwOpwBiMDkosael1ar7W64so1K2FVp7bAlacbQ
C8/lSIGY9iZTD2Fk2PgwMZdEkTcxGmH1VAomqVAljU0UqIAWdSoB5PA3CsIleyJwxkjWs7r6sjmG
DfDXfl2rUbE2HSCzadG3dxkZWsFLDXknottPO31Br8n2a5SC3mhCKaHuIPYUFbSXvWyyDZYk+C3f
VxljA11nsG1d9z2uuynkdpRzpxI8+7aFHVjoKbJ9ZQtcxOW9TQSmxw4tqyYSvfYcj27Wex9TiN5o
zj7fjAGT3iievq60z4plyGjefOe9Ltfgn98I/F35bipEmEOZgtz9eAMzqyqwM6xCOXCSprhiiIPw
mpN56XH4sg0pEGLDdE/lDkYz2PQYl9W8Qde8dUhWAuEldmH2q9yLgazir8qvIR6sZMCfdy0KnaRQ
uaiqHmvpSrtmL1a6V+4nCiy91m3Sj6XUYSaFEvh8oxEjYilEt03u7SIcDwMUKIi9h8hJ8HdqfnZi
zzaD0VO6GjIJlrLb+FVq8sfmacekkw78W3eee3UMs10hpph/Q6n8MoCBu3cRiQ6kKtWmr1zKpfxl
DXsJ+goKaD6V4TqKi4OlG0z/VJxU/5knsPxrXgArMp4nnBUnrzvKryGbpL+fJUy9AbHp/P/ERcMm
1IPVkbjTYgSZVWbswbWPPUat3pBkBdKusgNHC8XxMaiTvoB09RpmQilp8Q9LLG5b/M2TvbvRO3uw
VAvUoYssYhWxYF1aZ0CuSJgTNH00MfzHpY/lNYTq9Yw3hAKJ24Sqzw5dFN1+X3dC5orP3ApUbwBB
0Td0jgetCmldlOhedb4OesbjyF7wBehN5F+N01T8yENUXw+x0tvzy1WEG/Z+UHBgJPOgoyotrdZw
FDCKGi8GBML5ekSuFuaSJXfmvj9AOe8sHuZAGf6pYyChlSG8aFSDC9EHI4OgecZzNgula/QmxDI2
w5kP/zQ08CIotwamxBfqlkz9PTPJaqtatT1WaGNIg8W8v+ZEe9wWjZhEEqKOjryjXf36mBliFmz5
EVtHqNc3HK7MGn+ZuobmeC2S/7vwoOkU772JeerBnicHpWwAqP/acVExZDw6rKL3osHyQUPo1bpb
d3KcXTg7O/x51KDvzIVScuhUOYbkp1s4ipZpbXiq6GIzRJVVrY9WAf/CA6/fDrrXlrbDnVyHfCLr
U+i9JZvODbWsXP3jKcr9VYzgKKVD9p52BufHXqwdF8JBUcOP7Bt056/m1dDMAXhKTBwT8f8LWgkH
3HV+iv3gi2kBDBA0jvpT7B4vuJtgXcVsiuvg0UqsQdtmoh7yEyeD8mBdKZI/5c2u2+XQT2p6ykRi
d9sMe5kP1SakocPz7Ad2+zZQJCerVcJkIxdFUUO2re+K+K9yfnpu33g3aM1Rq7rHOkGHpoNJXfGm
3ENqkgxTazkAms4RMJoqTc8ZNhG/f9+0KjuTYQ/3QHE1qRLnk/yKdj6we09KTotOII98Vk+95yqn
Z6unS7JCcJzJ7SBUPnTkar3L05KvKQp358BAw8j3JjJRdK6jtMMVNCACInqKMR4wxn78rzdOBOOt
r+HZLAbSVjo4koFvwlxLCkELe0KG62MFtvCnWKqxBqZogUpHHRfjjEkUu2/CNrRwaR99F7cYQBZh
RHO8mN21z7XOxUkB5jz9HaDBzxWnfsTci0NLwSVmHkvkC1IJ+vH4gi5YMj52NDNyY6QxWthc9w8j
ln2vkaTQSghK/otV9T016NodrCkLiajKxd/McPZ4NcDiX78J3c45MgCaiB5WTeatPHu9wnCx3Qk/
VUuVPH0lM1EKivk9utNDjw1tgWXD2GseTIrMI/OaH9eyEWYGqxWh9VGjvF5XQGb0P+6ODeuVTdmv
pgtHGGE0S2HddCxXSVopegieFwhC7KwVR8ZBHLWcY5bhwsAjkMUNvjE+zXa6pm6JIcEbpsfJl2KY
ETSmNTTMY0uoS+88aoRxc96DCDDCrzfc8+89lPRZZjYLAYqu6IoT8gYI35ZozljxbYzN9iQO0PKU
9xaVdZ7dgF2gMWGZ0djlfErdLRiybzJnr2im+a+UcFbdiGJjxG0xH26ykxryksIn2VwA4uRXj5TO
9xFNySU8WbYH7qO2EXdAoY8kLcHAPb+39jklfHmiYOS6mOaAy4wn7qfAwR8zzUhjUREnvA7a5Phq
3Kaug9B7xSUQgBZhUhyncMU40K5IKKemJIkTqATKz1yPT+Yrm5E3fA1Pg8MoDzGZDKZgGXF+U7H/
5/1cDucrM/sb7imhzI+plUN6F+lKRi72oKsqyNP/zejwI7aSVxcMK459WTA/bEL6VL1ifF7v4ZjX
OYPYBNHJCrXablJT03eHgKKJ2hzN0qJDGhefkQ6tybVesBb7Ly4sEdVHYlv7J3WhMZX6E9EG5MqH
YJPyzQHQe2sZYtUO0mE2UN0w9HcqkdyoyfdKATIjxvgtLMv5UaasEWdg4ymGLvFFHNqgxe8J84zd
FPMn7FJw9TzLClIBAq2NYwQbhqAVTYGWB5opy1eU3+Wga0QxwBsW/IIj57NgOedxchEOI7woIJD1
cVJki5bRl9xa6NbY0w2g0LZR4ku+5GSejK5lTYUjDcogx9xFE82xLy+lWWhaR47dpkjjvOjzK4QU
FVwa8V7jC0Kelh0nKaNIPwJ5uvauiGi8vPzV6iFyIhzhmPurXQjZGPZ9BNhsesWtYwZUdOOzxzzd
QcDcOoNOhPpbVwZorPkT7qXjN7U5epDyRwO9veuc/L+BzlJb9ELVXtckGy6fWzBQaW81dzolS/q2
KfD2Nblbg1FKGmdju92K71sWF9CDeLGAPAXaH87g4rlxMUi38FQclVntORus9Y39AFVa4hXQGL09
EOHiIE1A9bp4WOMFSYVJI3nMwXjxgZ4Derpdh/PXRF0VVNW59vC2W20Nn6HC/rPqtnnbdQaVSici
3ixZdqSPDl//GkHM8sNVOP+AvA36BihLF7TRyHk/wRlt5jHcLgwqATdr/Ky+LhQrW5i+7Fk2x9pz
l0VC4YhcNrSwd6z1mBITCDtR0N/S9TAgAMz4aawzSlyFDomw2/K95EFkeOFxe3eIbCWVXlvJQcro
KHi7w8tYnktSKuc1gjen1JoLg/Vr1k4udJnTF4Dugq09GBYUIalG3TJjQkmsmkkNIrYow38Jz+Zb
tlqMg5oKrKVTB4Zu8gXFxyBBesvmjqB3Ek4IsP0YrNs+lZ42PRNYr0PjceIOHp6CzSupdUnJ7/EJ
WRtnA0U2NUIwAt43SOcj4fmzeN+n8hWOhxBer31yN7Tk4CyNMxqOX2eO7M4YE4xPv39v6Gj9fdA8
8dUUScUMOP2xf2zPi5A5Gyix1L5WJJO1yIGR80BaLoermI8YkWU6OfhAApy+K2Yslzioymw5A0Gx
KPFP8XeCG6hcT9mg96zXzPiJMXOwSfFNDSuhAoohrflTtdtQMHa2CmP75hwiP5jRA1exZtqwXz+C
SiqwG7tQpJ/o9bg5P3nef6X9T8rD+vcPmFaBZDG3GieGhsNeK8EWxoJA7MFPFOdC0LV+w9j/drBZ
JBLCF3nv9Tf5QwXi/kPGmbQAHhemWj+EqE3eGouuSh6K/U4wbiqE0nBsiU24TrmyBmu5fcVmkd4f
MdmtXEhubi3hZqktnZZaerIPjXvdwxJzDPuhZjKiy2+k5epjff8j2WSsTwp42Sbz10uayrXc3Zge
sJJChtJiPco85HvOkCgqANduGC35muj2dWKaZewbq7BoFAzQ2LjYoJq6yNQVOTf/BKqZ2bTNx6eB
/qmEl6pnJoautzuSmMOfqcnDY7IUwPXjvLsEh2WmBdT3R3DipNJrfEVqQIi53TwtJr/W5uU0Ha39
InZSu54fah+s6g5tE2U056RNCVcmZY0IBaG4JlxeQBmxgncFPUv927ME5ei/pJG4s40l/7CbPnvR
YjQK2LYD9mkQnHL0NB2PjRwKgUDCGD+U2xdyNpCQK1oAe5lU6OxExKN9LMIr5AzoLDoKMlAihEPf
gVQf+ijdg83Zoxv195J3x7tpS6uChA4E/qudmGtqd5yujACiIUcuHZN4X3cOaMnp0JckF/Tx236r
qhNz7CDdw5ryElghZzjYVWKEcXSI8taEn/ucNkFzL5XS2ot9wFHt8acl3pKpNLzX0JZm1fU3SjXz
uxroyo0C8LTXHkZSb1wcPiPbXwAsGyJRDZukiTswWgaprFyfI61c1/r4ToOv3IwdkAJDzKkQDA+e
tUWmCpdohtD4eeRHxNN2GuUVF6ZKZFuLhmKDKl+6ESC9DilGXcvlZ4/h5cD+MEj2EBrM6eXHhEMz
U8pN1rXQcX5fgyKJzOFG5+URJvYLLRLyjVXyx+g7bnpl+7a9O1e23vF09jiCToMqt2LGfvoA986H
KKtqjhSEqJzdj4uOCq+Ge3phc7IwkbyD0F7ZZgjhODcORTNlmnutg/qgtNPy9Q4nc7YiGPhP08t9
bymmoZKiQm8BMIBZmx1ukAHE9AV987AjEBg70SGXZpbuS7AN0qUMmcVEOu7faZY4iokHJRLZ+ZhC
R6goSKWn1AK50XnjloYLbkXiNY2Eq/DxTlA9JVV6tJ21pm/LTTwh+4HaX2FQj39u7Qb3Px5UIIUe
OGdvAI47nYkOm8yRJ9Z5HXPD44IavesqNV5P7tmvHa5k8rOLrVArvov+jla4h+Io3lCB84s2vvSe
/bpxmJmjXIXnhHRM/ekeFCMkFSaAMzL/XzQ2LrEHUqthRKCaQovmkng5KAM+KgdtxM9+/eoKgBpW
/F3M5YX3YAUuFqzJpAGe8qOrCfIP0eE4T8Ya2VEnDSDCn9IhOI/WwVdfv9DqhAtzcyXtVjPwpbAv
itXCSRep+CPrp9X2QoJpHxsVuhcE/vy8MOOMPC24z9COBhBYrF4QlCB74LL7cRgZpDyBrOdI+Vrd
xKYe40fh9WsP+ucWL4YKonultUzsVgfJITFQZDiMSTwL83RVnSF4zZyWRSFJT5LMpo3qDzSYu6Lj
P9A7fse23uZD9azHkXHq+fw8YM2sP95Uht+q/6NWVFOFSXTpL8JcgByRFVBDrzsEhkgn6m75/pr9
scwrsdbA8pm2W2GadXnvJVRn2RX2Keb6SDqDREGoZix8RuoLhbAOqpwxPnI7F6i0r4Oj8mVTPWr2
8aLLiMwU4uEGuUostXVveo46/Lx70bWl29gkLgSKzTOj2cWRGi+ba0ZHlPItsPMVALAjsuynUe/S
53596VT5nkx1ICnocsUvunNPPsG0EMlw3VnErrXBKGx30WAKh/qz0P/mYu7BjxU0UAJd9sGVSKby
KeQ/tiB+aaz8QB5K1YpBe7mL4cRHVTqbSXiJmmYC7C6Lm60pVTnXym3UhhRUp/T23jkXA4quZF1y
OvWPZjFBIJMfKTewVgL/H3x9SwUgPzWSr6bSurpSAQuVjpOgg0jeN+WfULNOwHlsITinbkD0I76m
rg+Qk3U+F4DPM2CUM0UubgHnmHg7x1iFJJWbxXvZjjnpOPT/f6AuWOtciW24LDkMFIFtTnyjVoKU
28OJ2FYC/7UGUGDWObazE2mv756GOgPlSomBYczVJ6m/WZvD7B7c+5iAD+t4ePwuR0yFpkescx39
GB0Pz8L2n9NncUi+vqlBScsiIpjmZzzqIAZ3r0Q50S60tNkM0FsbghhAT5TYBpxqbNAjkxWOSNFa
ZtWqn47pQga19ULP1hP+u8uA9FpQ9AmEw9GWMUxCWq1SPLIi8FD3gf+Ry0cyD+JEcszAuFkIoI4g
0gaYT52OGki3MMPIcpZzkZjERhelEXoKTlypu5u36qpA/axYHsRrLJmAD+CRFnHghOBCxHbPapf0
wiWH2MgdqrVcEekWCiRhWuhgrz5ZI4pSTdz/RYA1n1IamXvodSCL6jklEiCaiijaEthj0u57OSE3
wnHkUtdZqvRhq32nE+tFY7F2tlJL2hYpbmSClqeDyTXfwbUcWolQK6MDH0lXKEtSlfPqT6g7L7Yr
XueIxse0FmMo/LUajuoVSRKLRAZky4A+CfLmq9e9fxWHx53RRH+S4N7/7XmMQYTvA4r44MtBqKKI
WyTABOcGXFSYyXg7PglNusIiHYGi/GmT6+KojgBUmBttTUWp2TBG4E6cCXymQgVxVcC0Z0N/IS3X
/baMB6TZbOdE21tnwtOLUWPxhiEVk9k7jAdrGeHso0BecqDgRfXYkq8J+QrAo5QSNnMmCu736yi5
uLh0VcPc/tbO2GKFkN+Qb+PUvmXvUN/IE6wHglFX4Ih50fo1sEna5/3Fops9btWjYjwk91mCjCuk
IJM1TerMl2KytC/s//dZTUKKBoFcbufHHekY90NKu2HSnbHJ1DkBuYb0Xbp3nVEOK1nDECoGk4NR
BDEkHPOcWl6NY5WPFmlJblsAMITfcWboC8rfQhAOpZnRRJ0Yi6GdztXqxvOVW1jRqkvFpjadfoiu
yfbHE/q6s0YyHrpolVflSETyrFvN7XqjfwxrEr81Df9c0fqkRNLJIRgPHPMnmtrn+xqu/RlpzITr
H+Pva96onaD5ZT+E/MFS4RRyEk1bBWjlqk+UcVrS+rT86ElVHSoD4++NkI6sDqnqgC6dlR8tSWGs
Qh+T9XdxpNrFJtJCdXw7GXbAfbsJBXVEwyPZl1ap5N+akBgsnld/NHh8rq2gjfRbTaAKASNn+QGA
zwd1lBH3xql391AVtgH+39a651N11FrfVfI9iDqJtWmyH/69pjjvR0FDNzsGpK3PUf0da6oqtS+P
PY2tlyWpg/7AL8MExwB4SE7/FUxddERGcaeZB6gIzrOQyXfyagu7iaUXHLZ9MuIFBwh/Dqq8DAUx
I/KoSXjq5EjIzjHdf0k2xC4MvVw5R7QRplV/5tbCaO5UNQV+7gSQq6lJ9cf5y93YceWL2QdbiqXP
COTX3ctChrjagnz1pXivh+lO4gTQNmLqN2v2NjH50HmxugkwES4poFPhhzEj23wfGTp5hTmQW5+D
nGZJPLxDeY5vy2Rt+qgri0pTl2eaxqID2u/O49/cu4M7CIBiUdK2nmqMrv/DRbj3l1mUL2AbUAp/
2Hzjjk4Oo/XfBAtoxpi1TrT9luhqxM0yksE0cC1AtyY0hniUzce90FPmsObrgrFdsv7jnRvM/smY
BfuM9UTsrR4HaONC+xOmsZJ0Mb6eCJMrkD8KBHebDZ7UAYxdFDX1vJMzlBWdXhCfKdJfe6v4UHCi
HNNBEvQ595YxmjhqmGnwGPVXhzp1DR44ZqKsZzRbxImYfQ5OMA5DhpFEWlyd0PX0Kgsh04gxL+ui
FMNCOSZF06D/ooZYiBvryhWJUebim/8CyKrqKGBaJeS3QhMbQaDvheUmr91l5Rjc3f1jdarAwGrE
mMpmeL1MpUZOXx3HqNgjquERGDLSf/wExAPXKWRqn+bSZpHm2t51Xpye/5SEQPkPVYAo6K1Ax8w+
fhdTD2Hnqt+KbxnGXbSvnis7R8dmbdDX5damHtvzcWtLcDRFve6eq712+3qtWMhrNj+Cy4OP+aIw
uZ6g0aFTbE5UAYGvotX+U9q2qsU6v9Df3p8Ia+DBwm10R+LkSDFwKeGtGMdI1fXQei3Gq6vfxpKh
jesquZWxMaqBUtlKOrgnBAxkDOKJUhgbIh3TrZSSY5DxN7snvilJzJHqbnERhMjrx/NtkEY2w31f
BgVANEe8eQYqH5FOXTZIxVwwgNdCXfv1uxskmqgu8lqwzLaBa5QY3PFRUUucLeUp1AYpxEpNRNOH
zK6/zE/17KARWwirYXs5kahd9Lsq678eBIPsRb5pZ9mjUnfIaZ12atsBTtapwgbbxILWxUxYaIJK
B0Gz4Ehcmn4DVfnDph8okxd3ZQPWQRxs8bOnIjX5h//Kjbs2+IGW7Wx2G2dsK3v8AaUYjrTqLY3a
7+x5NBHz78J3RiwAnVEyPKy2C3AxVLUZ5jhFnLju2eFa1LIt3MlrC9regJpNC0eDU4V5O10PAJ6O
xptedtA9ayXSwAATJLhFkKcfXc7fQ1yJ8YC4zG8VIv8zjMspz9mwhNOaHvcZdVDHLzfJujK/msoL
OVGsne0B50TvkUeOgSw/qY5ZMaeOGbtLEW49+VXp2FOs80qnQsC3LtxzUL7063CS8xMkhgsA0KJH
ApMJa1wd4WcP3CALWUwH8Gqsq+90+LE7gSdv45y4YEN9nI+j+qoI1HeFNetg13L3wxFJp2tkMT5C
4rmGiivxqXsyDA/9c9dOlan5O3uFayApSC/yYJAnrVmuPXOo61r3aEW8EiArTXiB3lTBo7p0mzd3
k7N5t2k4SQqPAcx6TiXFl6oEEwq8APBgPPDslJUXy7jQkHEEZY92TM9b6XkSS4lCUlkk/eX8REhU
sMAH4ZWvi6cT4ToBeUO7C8rhfxM4MhdPN/G13pecukbWNe1bh+SUg3v8SRI+wzPOCbwd4/8kQ0Vp
w0D6WuOPg2IASZYFPazMzjAVwNTO8wRieX62A2PDIGl1OPhjhAc2gL0Ys+4HcraNFisQ/naoT50W
nNhX/XiJ3vEv98CLpXN3Coay1hu6jQumZTXh27dy8MZ6ROQV1JQ2u9lCfZuR9IVCBVt2vgSn8tnV
IGJadj7T+5bX7g7fsS1SDHTJ92qwVzS8rv0dBB/DUd0Sb+qhqPiKEzT+b2Oq1NcA/Sp8xYNmCqXa
+KaCMf+ZEVU81QWU0VjfEOjK57F+2dmKpbHiauwGH/eFUe17ADvLMHWX9ixKdiV6Lh4JgkBKMwzW
uQEnvQDPb43Ln/kICzTfvs7LiJFwS2S3LBPgXCjU2PZIF9g8rql15ZsSdQJMh/N/5mLZSunwdf3C
/cLSXRt4w9/agpRVp1kOHaK+mhwNqudDndNhfugv6zFJLE5nZiZTfVqzW2xJe6polZjpajOL4hq5
9W+NIaRLXyRqgEq7/XTLFIlDuHbYvkUcPC1wG43Hn8sfWDiDrD7/M/h36Fe1+cHO/2dKqdQeQzxF
x7wiKn9XbeMlvMn4JeG2DcMdDxtLLohCIWwdtYGHCRwuUBh3DX67XkFQ2YAAGju4LSVFcb2iN9Lc
VTm15Ltq2g/ntT8xEgH2A5jY5wH+GQtiZC+IRQzm8G0Cv9RNeA7FNPysGGjoUAF6tbjpa+qYcX15
wx98n94ZH24T4AY+uphClUKZKd0ehvb3XVT6nhZR98bQnPOsdJHJV2uogArGLb88uShBMAYzb2fq
111VVB776lCDZaNmhk1d7rYLMAlVyE8SAizzLHRe+iJgM0AI2Fgpp14tBZqCunh279H28QM5628h
azjl4bTT0PeNse5pF6GuEpkNGz598Am+Qza8/hqUx4EBm5lVYlJYc+ld7j/MdlUpYQgwUN+UINgr
WhbSfbk1Pp962q7hmEiwGfkNfm0S6jMMS4dZX5rlQntbBfGOPJIMOrfLcCLHx424lM8QoTHCLpKU
kiD+1eLRLu7S52H2t29fJCwok3/+KzJcOdlV9hJGxa2uScWkUNrdryKHfAGzvjWTvYiGK0CFGET1
oYzp9AvWlRDNCDAV0qv8bDaC8a4roPgAXQHrJGErEgpKrDyUfK11eN6pwwmRpQJfLDz+Zlj08iKj
KpdGK79rdI9S5fOWspHgiloH7PRhQWeKuXj3xUYSEGnH0e5r1/e0N9ufsIsnSS5Rnb1psyHStnCL
YLRJpU4FEHTV/1bbvP3/8oP4GKC/hLdCAGzHX9Zbmg8qrxQVkSrLK7h8WI/VtdlaDBy732nm/STi
N85LckN1He/iFJQJzelB8BAB+T/M4PhPetJu/yk9aa6ed/E5F89yWxmL5m2EtGM3L1PAWz3Cp9z6
koKQ0edz9CeFfAvJJna+OxoQ+sIoZwbSPNdmpoUsAQwy2DvHM2MZxdUwjwuLSUGYRqvtuOrCks12
q84p+jxIHVO7J3cf1+0nxvrX0xz3QZlkS+sBI1FVLzFcNP7FmyhZBAPPkPyiktNYv1qgS1YxDF6t
3tsvslu6UitIEuev1bn6ekcp1uVutL8GgXnO5j2zq43jQBd85rinGmU7CYnIeHdwEEwn1I1XpfLE
sVYWeVYsPmTe08oTlcy0AfdOD6Tq7NVR5xMMPeflNeIkWu98HH+BeU2IJS1C9+wnG1lD7QZS+qwl
wOLBHFAB760H6KV8PB1OAbCwOeR7NDPfJAIKrzarHkn7ppMWFryyZuBLiASGTqmsWtgamZn1mwNw
lcSpMXR/ucy74xWdkJXMuXsH4qd3eORFYz9GvTwqUTRoc9CyPtgDMnxHFM4bG3H5pBbiR6iZy68d
2n9bvR48ue9uorVSQUfe1BH4Q4u9K2Ong5m0cs756xV/vYhHejaWKIXP+tn03Y6qQQv5NhdYG30z
QeKw/ka8UWAsEJOmcPipO2Jxz6wYGXwz4vnWAv1JeVnF63NfLHLFx6AZFqE7AOAAqQ1mmJrPuNKo
eFN9uCItX31dHgLmHNBlby7R7gwJTAVrPxo53sElXHv2gaQu2OZvD8HzW1zjQ2TycwoyIRfx1f28
4Gtr0nUge2kKNWXqTnwkcTD89HqzKLn1jtB43OOO08L01cp54yJ1vs4mbpB9PbEw3KGItyUDPyof
74wCazdAq+sH5o+wcgDs/lDuc9iXHeaVZ6O06AuIVjmccG0Oyt2zjHIXU8L9hEsNFX2lFwwyBpN9
RpRbJ5rlavVEQsu2DxS9S9Xh5JUMRhxnXS2iKvRoiEWqBCnb4St36PP5UWADjH8k4q3+xjmxrJl7
E+siEmvxJfO8Bs+Hb6K34jI/fBmi152iay5zHgnNxowuvbIbFIOE5PvaBE3AAt48rLiXjZt6hdba
C/D3ouP4Mdy2bM6GK7r5oexDAKNDhi67AsDYrh+L72fjZBNpPJFu9epnhJCVwp168b5zG1g/sT2C
ST4q7Jw7qz1YNKEXa2gQAyx2GgZI25LG2VTv9L491RLmlfJB93+Gu3huL1a1QZI6b1p6PjHlZqmw
8NiStFaiir20t7nC+KyBmp7hs4aJ9SykopDxL86VcN++fYkFRMTamMLHueDs8akDMwx2hItxhRBA
cdGWnat7+fxQONWnlcI2/HMYd0Ela30kers+FGztvAzAbO52pJidpw3td/+1S2KZvc9wNwoJVICz
TOVeGfst5Wm0w33MiTRojZHNef0kKZRcQ+P+fShxg3UGzuYX2bPrqortyB6r09Nb/uVoBe7+hX9n
BOJQ2IfGpi9HRN9adzLKdMZzqVHQYjy+NHCuLDfX41a0NXaMLyYqEKRF7X/tYF43EnmLQ4Jz/iRG
ZJIy/zxZMpwM5OvWolovrLZ4O+fFR61D7H82ItwNyfgGgTld/Eyf7+INlHSBlo7Ybsr3jm/4+znO
ekOOvllSXGwP0CbcBs+KO85TXV/3Bwaio8pIb3KQy4TTIeC+RrHsDRlZKjZsuWnGLNLCTTfasr+Y
DlroA6PYQDv57eSbdd6U89wBxtdX9Or5xFZXcL6DTvLTuFkYbfiSIPbMwHyhB1nngB0UoxmhDwLm
NvVRFJLzPLaNBbQxistQTkBY6//Py08EJd9Ie/nqi38SGbVNUTDEXfEm3svviUZ7QOCXCXn9u1iX
njcrdhVr02D3w0jDQ+jFkrdKLO0uMh2gmlFpg2TevAweZ9Ne5HqRg2kONjGZqdrsVQPqc7/Q6kBA
Ky5im44wII1L27ub4Dx2DujYhjLaTee6gLNfaNO70kQC5uIws1OmASn2SeqZ225KhUF7qSbgu3tX
bG7Zi3jggzKduCUNlSJ3hrwSvND1w5eWzGtVX2q2lbfYRSo7xBc/+4cDBKeb95r9Z5du9vT/qSC8
Gr38t8dR6mQuU7xN0fl8juVpDqpzip321sTvX5/3EvFgGkD2udcwjmJ7OInnI1pGLusCsLAmVT2H
Gh2vuxMK4ycW5C5sSkMonjJV6acNyhkvjRODv4HR1wPCSO4tzZtY/t3l01zjrkY0O/Qqf3YW21I2
djOFDSZUeLRlzxJa1NS8N4ZsNokX3wbs7+r4SptmU2u69IYDgyhKac9eB0AxoddZiACiMnR+D0Ql
3tC1SHJUzA+k5FWoI9aUannoDWOSH7On12PeTZ7p6ppT+iZGQQ86wMb909Jx/d0iU9O4uMql5aWp
yR8C9NQawT8qbyKl9s/igvmwfMN4L8xni7tl9TszrziJuqjiDgLm8RyMvLsXlFbvy6R1Ajn/exjN
BLh3QeL3hWM5LB6EE08FF9V5Om6UuwuXQe/MCXT2sEWXkssm23h6W4Ra5XunRPUcf21FkBu9inUr
XzVducqrfWQgFvbYSiWcZCOG3aYwdSugGekDTz8CPJfNMl7ArzrpI6tF0wjcigpcBtjKOdTlriXp
8D1Onz1jFxAiglrWqHL6gf/iUixFYlIeyIxWY7jP9TbDovODzi0UKTiBqVDmT71X/ujL89KJ/1bV
dQ+xBl9Y2RpJv1e+H2Qs6i5vLwBgDNk98K84whLpj1nvQM/2nLA9xPeOz9Qzg640b8dkgquTyBK9
SDaAzK2UGEoAnfJYuNOdov7Iew1iMwnNCg+qgJUUvR/STLAJ+Bw3Sw5XbKuA3Zp1q/vq4wsBvWCs
CA4oySpFo+0zzwdKp2xVe0ijhYteGcMoVThuNgHaLD/PwdB+86ca1+MS2TZhG4NvAZZg2IRVsCTp
ImXSUAD+E5haO65SwUqC9IbI6HemVM/jf2Yfd9T4qYWfXCsU49sO7wcbc6oVPhJhPHBf0GP4R38o
IllsK8cMAuxdVBENklmutWtR6wYg3Oj7EN4oJ1VaNdfkvwicSAS9xZ18fZJU0a+rpIyBTy95CrJp
5E8yLjBBlO5sG/Of/hM065SdFIsYVj+Dka0nsKc2lOkPIRO8Ft3muZbwB23TzNy6SrmEEfZvvpBt
vqCBxCE22iHkZTfhEsQxptLB88t4h5ZcMoIDIEtqKuKSIevKEYhuSN6XMwXsceL9vM+HhtoTgI7E
5DD8qGfpeRqUcuiLsIU/+NfIbzC568clVZpLlDRjQaKy1tJZSic72f1ll33P240zYYPUe7BAJaym
Zt1sMSyMb5foZ7HezLOXuiyNedOo4lAHFooEcZSahFBh56stl6cZ09OXsWjGF1TEPz1JI35Qgi5c
dNDflQf/P5Y3uaisxGN646d3FaIFR0Yq/jYhDmaLLmVgAO/BS2rgo7k8LE8U54c6W75KNRCnOeD8
QrjZorvknC3wp9aAxzPOakpXUmXezAONZmmq7tfgRRRXkG7cHUqHdAu06PHNttZ5IXmk81YqqTQz
gHSTXk3ewIAI7OfYTqAQuJDp2mtQQvznnAmvO3sr1+m15WooGkIM3bTcFIKi2OcbHPQ8QIcKg+kn
zG8So79uz7Nn1hNa9kK+cZ/3EvvnBV6OHnTScSfG1e0w1MG58Er7Z81zicFVFC1USHbY2QWlz7fe
WT+E50DPJWxnTFV0Juk0D54pLBiSgNevbeeDydPMlexGFsQQVVDX3dz5/qje7upX4aw4Sw8l3Vch
tyBlioWUwR9jXuKoFwxZd7q7UtSCsz0NTfn/onJh+eOjnZWYRgFwrWx1NRwqa7z0grEHJuL2Y/dv
Gs4HIinxJAwEfyf+NeM87hXqeGIDrWGB+xQIXbueCrGFWPXG1O7zatWs/oeNka20Qz4Vw0RStwjR
PSBEc6YBDqfSjU0/RmcdH5fxljao1wpVgbTwAIEKi9NlC5wRc/HUABTHiULzmjCV47m4RtDXJqZe
5GcibovZQ1NKxfB4oJtXVRDfEmXw+lRWugqW5PAS6Tw9e9+rxLpT2oiAgUz7TmmVQFY4Q2Jx/sit
Oyeua+UFw5YiIZxWzF6oravKMl8sHcMIpaZ8W2h1pkxpV4N/2Ey3W4HXu3t4qjTHJZ4YbIrPy0sK
fVde6WN2vwEwify7jpg3aCfmH9pxu8grO5T21oY4YGXQw/qPZR9+9tFN5oKSYP3pL6jioohkxmVY
OsOOaPoV6lwk2bStVYSFWwau24065S02xHCT80u+YaAQo0596pssIGfSMSX2GHZNvYc+V86vPiuD
Rpok4CPiZlT+3ViLeuCDw5DqZVDwfApDLfjcOPDfqnE4V8YpwdCjYcNPC3W49KWsyMt1rv4JPk5j
xLFNBlpuGpzERRuEvEW43kvnh4Mu50mGAdpi4Ds3zKemktHqVKn2I05vhsPEbOkKzOndU9+9Cyq/
awGlyDkw/mO5eVlxZZyD9qYfRDAnhMoVrufREeez3VTxmRzaUXxN7ocvMELjXKfs7WClBQteUwKv
c/up/p450NzO7MBtL0fQV1lOVwL8xxflRsM6KJwYl4i3N1I5RskthqVtgqPCBR+UMK6iOqNUj8U2
3bQPX4fuEThFELw31y04CLzzAkzjxBQ8F8lFZkFCGeX1qXZYK9VzRy+YGgUcI8S3zG7azSLy+vjF
cYv976EXnSN7/5pdEw4ZsddmYcH/bLGpx/Eny7z6GLpTtVSeb80X21JeRPa/xjeQMw6T3PIwmc4l
vq9BXPrAcAhMSl47Qllly2CUkS9+6jGdzv60LQkIYE4MkPYfjaGGay3YnUAqspDfUpeNtFHTv2Bd
6ID0fZggdlQdPPjw+hnoPWjKoNgjiGpoPGQyoEq7Hm/qMq98HjGOjAoIflPQjGEt86LDf+aiXfgL
oKNtlFPo35uPn5MUn4e0nnxy5ToItN162XMJnUHtxI2W6NCaiMRmDcEgtV8xfrCDqoxjHNIzfbXr
D+IComNQbizuInSnLehZFAfOBah92BNA1QDrlSHlaLQklXrEpwvLwnfuc2VquDbjqgzkD2SLJh5M
8j5iewRbhtmR4S+Ctnj19KJH9SzFKftoYSLT5Ttqr6YkqvEQ891tGha+I97s5kd1bwkCPVywWbPB
svdQ1YCeeSsIQmGZNd2SWBSn+E0rC7ZPO1mDt5L3WlaKKpoNnz7pMh1fMrk/Tr+D+Js76acqk0Uh
rUnHM8q9pVMx5Tp3P6CJBytuPVq64yVRah/gUoL8tPi1UXnUbQMMT/FYL8god3eYbYLT9tPy2MwD
l6+2EHv4HiB5CH82nprkdjH1nM8D5rHd3XvoMLHxHXAVIQKDvie3LYXpJnSjGir//Za0bXp8c20X
1EQKV7+/U0FhEDaDBD3AjuJJqpwIEpv7ehIvUFSEc2aEujVJZ0//TFT2xZqs+tNFnusPb2ekAx2w
NnMpDB9+YSK6/dzmvuiVinhi59/W7ye3lgmUtr4E0e+bEMT6orN/n4Y4QoNiJZVLQ35I7sk1tg90
531YNCR5XGqVSP2IqSyMMWCapm/GKkQP4ZztjuNe9Wm61yJCDBnUJ1BM7v1S3eZlhBecX+tH8U2w
BCPvQulCShUjPSb09KYO5ESrU7oXK5XI8eSPUBmoPdmPx7hhXObVcMX6YTQHH/Wrbd2g1rna2zoo
WuirevFOKiJvY6LvMrjYiwVGx1E/Ks08Uu8dQTf3Dc7EEy5m6P7+kHYkZ0L7dAs+10Nf3SwTRKcr
vZhl3CVmULEO/yQX6z7zihm2YBlAh7vRAfacjbY+nosF36Mp6AJUYmh/lEqiGy4fLioCi9QXhdcb
L3jwD2IcMRJkJ2da/mWdtkihghh94TxSmRlkGiR6/IvkuBdvyvMuC6TAJcXm9t0MNGhoBvh4gmuK
BMLs/RLd5FmZQshMvgcn80/oNlh/DgpojDR33C7DAIDU9AEPKqWYgkkGGuamMVN/L4FkOPS5n0gn
A+9k0iT4UAa6KnPPOBLBAsJjtPjV9L8wlGmAStIV2ost+nX2j2G66fT7lN3z22e7OynbG2tC+u4U
9Q2W0Mne1wsDRF69uh5R/FLjeyzcDpIgekcJQqFp9WYxqAAzkHhfB89AcYlMIPV67HxUHcFasnZ2
j/O00q475rKZwIrkMpX4qvqL3iSG8CGQ2NWgdK0xBwPPI+9XA7XfAy4ZGOtz35y3WPapHBNrq2vo
d3iuMxDLBqKR6dzDOLhNr5GyP/Gr9hwCXxFagivbnUXQXvq5C9dwkkh9jVXrOEJYJA3Bw+pbr1xw
+zVCOFx7H84+botW9As3pAArRTCa4FawUX1BiNvVcRQO+pcag+l+Wb0qCaLydsh5AFyCHSZ90tkX
u7ZvzHSuM9JAyuolWdGQK74jMb+9FOBAChMVzJgeneK+MbXV9DpMKkdKLn2B4tUr4T+FC+KNUl+r
8SW/VSmyfILOYYANRwlChqH0WBM8bNIOiEGAZSXagdpTzaFxmnB76P6BA8byPWt0WnW/tqqUOul6
28MPHabC7vAKv8JMJ5Uh2y3oIlfnynxH0hI66VWFcnr6XADU0rlVETt3EEhoePmDmDVdfssQt74m
/J75w82f/a5enCkRwz059NRHLoQUCH58jVlymm46sXVSt7zDh5hdmQx+rMWEt5P183hfQ2beWCBc
VR/qTsnHgwkSKxKqfec2ZDxYVZdlxjpa3kBE9vN2ncTqgDpsdnnTjJPtryF2Rcrv7M0NkgeIUpQj
78dE6QK+OUfKCBe5j/x8UnTkxthuWibEEMmf/lYpu5lkitHGh3fEy2YiB3ijNaTbQ9b8WqnYXcKw
k+2juuNmTd0P4LP/NuqBvI9sWFdUhRJjIRdLOuZnn5WoZUqzxdNWwacff8mGhtr12L1jsoAD8jRo
Sbg2k0PES6NQAQYptMtCefP9Bz8OXb/Y7RzdRJn3lMhmDjQ4a4mFCDudD3X6idOfPVdOquU8mcwm
vS741U98j5Zi6GW/3w9gA5VtIsryOwbqRddJMm3/KA/5Yw11vBlNH6voEqBBaqITJfliUtxeT1NE
cRC21Z8Vx/zSZBPqyxAtFMGPlSB2338hPdeor08A0KypWmq9NNSG5irHBkYaFjHfavmdBwHETCj9
dxwRR7CnHhUNP4sUVgEPDsxyusEvpOfkAv6shuBmmP0qsuoyEJK94tj2caIZHnB/kJEGgLPsT/84
5YBP/HswtawQ/XuUsj7VprDzgv1IXjx/qZOfaSnHYF0ESF76mNxEj1Lo0gcHteUGVD58H9WeJev6
4tq/AF+eEMRLr3+FPZoBLwo4AfL0l5qRwR5ubv6JrYSK1Mriq+L2e4PtvQ4Ipxw/yqzd3N91qloz
UlXiwUk8zL6BwanU+AJc3hWqA2iz1hlspURORLq8MaZ1iPLaX+YQKWsfWKs4Lk1LgzfJM0hqRbrA
JDFf9OGFdQRCfCxzEZXFkgR961Pf2EzAy3Rw/DXjy13Y5cQrm1qKKxLJbzgjVqAB0T5ck8U5UJOE
hgcIOvI+HPBU4vbR0XQr6JZoFVigZ3zJrpiM4vYK/FID8Ort0sg71j/HwKTtgTu5vtiXorVsgPfA
EnYGXXVz1MtO9sofXMdk/bH5AFheiYcDFb0JlcKs3OwOCbMKL+5ljbIvdqKgbFXij9o3npFfGjdH
gzOxVt7Cvavjv6ZyfF6Q5x8Jzt0dzM28YGWS5cooOU1mfWeh01AZZVQdzJp1uQVNiwAj7Tsyxt1B
XvtUgxHhn/mesMmLk/2Ps5ou/yNm/n8p3KhDDbRdK5R6Rh+zj2lfiOhNNGRwZiP23yaj8ewRbG98
Tx0Cvo1QPU8XmuXZR1Hb2+9wC3KJeiB+WyLYdvUIDTMX3JFS0dOlyzpMpR22bIYh2AQB234SFYQA
d9BPistOPjD0OVJPup5A2J1PP4dDBMbQlDC1RM9F3wWwi4N/4N0L2VONkihkQW8D+o7QpeR2Ryvd
X9kODklfTEN1b/sK/Es+qu1iy/tnlEGBdY+Enie0Uho7gn6zkfOeOFYAFI7C5nrWscuesTEqPVYG
Sq7KJ9rDR2oVcPBj4Wb/Ji3haiYUCMjSfSyy/pjafnCWf6Yh1uTI1GsbZCcSMBhVdpuptcudlFw7
iMbGqGu4JCbuE4FP2bKAr2WDdIdLricyEg5sAqjVwnXaUd9ItHa8/opg5EPOf2p2+wB1AlTWpjpX
ZOeQmmYqQAL7O7ZIAPCDf/FDGbygdd+GyKJ7iFj7nTirM27FjcVnbaQ7JFwEwH9giPHg4dt3TpJS
w9ozS56N+yuE+Ru2Lho9UsdGfQKAu5zNSORR1AWqQpez2O1mm+bWg3dUjoPZo8fsQv8ijbQPyn/p
rauPxuM5CC7sDZiVvPAHqiDci3Pl6WE4Wpz83Hh5nWHdIiz3cf6u+BoKkFNHDLtlaXKrpidrzT5U
iPqBOEtBEKZzUmOHJRWBxxn21vdoDm8g7jFu/KM1AW/xIZZwkAq2uaEkQG4gD2DAjsX/zLYJpn3r
nN3P5L7WCbpWnV2hOPAqnkQm3oW1K4vJKWv+nbEjWy/sJH+hJ1PBV50MYjbRdeIN0kV7Ea9KQP4U
nVrUdX8uID7DH19SCKPjenY4gRt/1hIkdsGTCMENnYkEvIgUAhwtibaohfg8S9uLb2RbCw/M3oYR
s7GvusBGR8xabxej4Mq1d6sHCdf170eoE9wJR3u8KNFAcwUQIkwY84KVQfPiyifi1YBcByo113Y6
LY49z/pWWdIiPQq09pc8NVxUVjdCbhXQOx/ghMYrrkV5CpXg47cx4iGdt+XfXqNknYZDaKJr83I+
IaGUgPXZBJvqcZdkXsFmCwDjroNwkIexNNLIxaepvA0+oo9ZK9hQR4UVxSkOnPCq2zpTxemV7TFy
ZsQfMBfoqpC6gxE2K2JMsU8RSJyezwiIxr1czUcoAUcbLwy3nVVzE9cPxv7gSkTictOqFW3Eyg5Q
jJfxa/pd4q0qWGkR/RlpwtaEgdvB7FNJP+LVQDgdGgdjPslHFtL9tUlUSf5uJtJa82htHRX301v+
ZxAz6B/N61xLyoieJzHkK5KaMG6mGLxDDjg5tGEDEL72H04mIYslFFii9fkzo872qWXZNgFFDUg0
0ujm+ln6nC2lzbIRGv8NPBeQFGkuS486A7SfxuHUC2KggJw1EJvdrVVzk4FQBVxA8rcT3NXbzv5W
BxRokKsNpGO82dMIy9A3BDUpG7w1KQPXzaAHVux/GGJtatl7ZMOlTX+vNQHZi4uselKVv+aMU5of
2kYuixrcKNGM0AAxZpTFtpAlK51+/dPGWADh5t+IaI0tZ44yt9Z0IIXHnWJHswV8nVtaHVJGdSPN
Ebi2LYhNtai+u5Mv4L/JFLxRmaO4ruK0ALtdkVMmmPDmcx41oVTzYUwlxL8rd86gHbBjEYAvnsif
vV6q7KD/lJMW7GdKU99/nuH7fc4yKCrs0SnfA1Yx9AjVC6lWpdeUtnbqNeF+PrdXTFDT6rkOJtK2
CgyhPwJkf7rIqHDPsiyOcaMaTcLE/Lq5u38Mo/tQ+y6922AAeTlvzyPiN4I0WDtommhLTa9j8XLa
aIxTOu4DMwE4odeV/MHu6n2lh1WLvOQ10x0nmDtWAdfXULHbquM+xlHWGUsqRJXeaERfFaKzrjyM
BlDnn5kglc+p9MnkMfSC68QjJiK+8KAOhRFQjO66OhGo/WNbUe7hB4sFuMSBq5lU10NrhUzaIr0R
FfK1SF/wk92lPanvVLH8KCci9HYlGWFg5mqs9kCDm7ii9rsuUwUvqye7JsNpT8n0oqFTAa4Mp5qm
E4FRBnhyc1erqudSlKWRI8eYd79Zf3V/0TdoRQ2vmWOWeTxI6TG89pPMWOoT3zwvyP8BqZquHK/D
AqMu4nIQv+FWXC1BFXGA4GAhTY6YUGnyDZDpF39ChVsQQckk9gaxLm0AjrmJKA89l4O8WvZVA7qH
gg1MfGJrobP3MD/tlLJ4/RYTsAfMXDHLzqUEL4T0bNq1gXURw7aqo3w+/TfGNwfMHlyvoAP5YQy9
vs27tkLDhBdrFeJ/sWNXJuSPwbGykAjU1HBg0cX9vxtxOeFaf7gV0L7oqIxMDFq7RG7WxuclRGYd
cAgjrL5SGuvNSF9dAVa2PO8dKr8m0Mapt20ta41yOrpmJKu+9/RS7+s/P3OO5uORZ9/G8arTjezC
KIvKmAMfAkGpZ5fBa1GsOWADpkSk4VIM2akNxfmedQWX5qRz2KJzVva0a5ivABXUSjr+I5/+XljK
iNeCuAWtLQR9YL4Txl6L0zlDitbO3+KnHM1OUFtOknK8GjnjrUKG6Xdy6qHrEqwiNAdRHMLHCe31
C2D7gMEc6TrP4IjX5AU8pctM1v6LBF9QeAishlZmUBPPYnkQmOGLsfhrcmWyn9CK0MbpHDVRkCO9
e7nqRXO0U86+e2IrCjGqVDAfcyeZoFdAszKTpQiwcvaYc9VxOs2sdhCllnunI0HvtZIP08QpEFT0
11Paqe/kbuasbqk6F765ziuBRd4SGmPNOcBaJsAPTpt5fVA5vVzv+zlPPZGSXA8AZ333tRg87rUa
0yJwHzX7eUvAMsFpZJBV34r02ZmH9wWvRPX/NZqtJRMvWi9HoEsd4HxDHgLSK8S4EJSxvBAuGQ2M
7cskPsWyi6cdhS35Ea9PQIpIMbTK9XT0gpeoONQWLbWB2IuPw0iG09luxOZhR7pExuwEdczg0act
lMewnmSAAEl6X8l9uWQJDKM1gIiF4HYKH64WBLWHVuJb9+rCRVsBUlo+BMtdHynFtP9IaHlsaLXy
+u3S8akFXmh9zkE5H9OIkezrS3+/NWz4PTRYUp+w7rwvIQqX0ZGeYOj5XNivRkMijsoDMQ7vddzq
RJmFMOhpF4RtTtNmfGCyMm6p98k9TAJUQftT3zYos2/OBRmY1Hqsuvg3EOPKjUUHnaba8BcqWmUf
1fNbcoxzmisbCDG2hgOMUe8IkSp2UKinlfD627RDWkNr8DKy41tabtfm63b0j2ODtlSRfywYUVVr
hunI8vzq+wUUdrR0n/kUH8gv14AYEChN7B7IrYeYr2y7f3i0bdcwyOlmIzEdAxwMFhqd6zDCfcvx
hlRxe/29WOT34I2UurG7rvGNe+6vhK8A5JHlYLY2O8wqWBRfRYYgCpuOV/fa96iyRRjjXOQRcaQH
EYIVri4+W9+FjVvu195P2TrTE++oC/29vbSk15NJ4eK1pcaMfZaOFL4z7t+RzjnXzqszePhsZgg8
zzib9JWaJr2ieL6ni7bvsOQ/FHjgcDFaMqiYW1ju1AInsLh0aswVbFLqWDs9I6QVnsz30kW4bC2O
xHLVQcTiajH1mxSIgWLZqu8W86Bi8UvsHilVUNIWVfJg0FJ6cSayYc2hMxQ+ktOdXixd4XtFE/Kv
2GGmh2fmGwdnr/vn1Ad4akK+FBreQWMe+TJ50e5aMfDudkwVr1v/LOUyvbiQc2q5M3qHi0hEINFJ
xIT6nnQAxWfWPHkEDAhxdiZaWoYzMyazS9g4dacfXu63HJ0thYhCaqX+mvQZ1IvKb/1FN5GBMaX0
amZfkV+vb/+4MdvPt6EFoh8Yzj+hbXWd8QUpEnyNL0qBLwUIutoTSvitVLOHDK2t+fyoxLcaqqPw
RZnDg7pVSlxecBwZFKo2rZ4Y2GntxnawFsImZZRkvEy5m1LD1jkLaywRHXmrcQSbCvdTGd3re09G
xIIgyfyKXuvU8bZEANGOofDK73FsfvXAWOLz0par2MpmgEpHLK8o8xeNDJ8rNjJXWtMYJ6UiU+HS
eRnT5aWCnqFF6xd2P/AuhTcKgO7Om8zlX6Vr4i0xravfZHGD9hg+wGB7L9OJz0IZ2Mn68PK3JdV/
oeFox25RL/ByhL0qDzJ2kcBF9bXRF5LqDJxMbydKntZ9xjNQ865Y5ufBfIsdpv+4cAv/Zu5bsS3N
qKPxVA/N96KTSzsq0mk5xhVSUusuRv7mGnfheZ4aEa/TdvrUkgi4N7j1vvwEXDoyu0dZRIFTU/Jo
1KvDA9YgNp6RYQDtz2+BjMy0ZaVhNEWOLG/cCF4tHHeD0YvsMQ8OfyIEbSWOXSzO/v7z9y7GeSz6
uV3Q9E1KPB4LLXqQQti2ZAjBYE0QP67BbOlKSMrpRhWjHOTxXymPSyshEuK+EijzqmCurE8xGe+k
PcM2MgjnEVfj4riCor0hRAfQLgHuJA6Z+hXZFnRsf4Kz3kp6gNcHfKlWooA4pRLJouseSEHg498v
A1ECML88OUfQCmPcLOCE0p+45nf1xbhCTT6ORBAycLsADGYLs22psDIZ9giCnSl/DOCouOjBpliM
Lug/yj5M0Fku8C7h04tLxqoRnN7A3+31yIDC9sMtIcOnpmPGxXjbGyPhhomED+SQV83AAVQzra0k
ANUvwqshc/WZ9pfpIvfo4hY1bRDVw3Hf/8YeRX5FBlxhCBvWwXGH+GCgWwssPJjmaCvZ9LvzIq2K
8gxkGa5HzMQ6MaOYwT8/9u0oK7jjtmBKpIuMiFLOo7jPDFkQFyUcvZoPsDSlmuQO+5dbKC+n0IEU
TeT3uAJEb1NeQxQj1PlYOvEKETFTX04zHkHTeZxGG8XJMTQZIyqiy1chxsiZWL+d8Ot46CcFtt7k
FEhQmvRHFEqDkkvwusWysZrMB6YeSoNpMS+zSPJO4LT5QoQAU/wDhcyacbwGl73/1+YH0hOHthCi
WoUmRXdx4BdfA1geGZGGo0N5ZsheIHHtS2IlmQhlGVE1b+dqYesWkrq5rhczE2+c9OUrir8pV2/v
r7lQho8swBjtB707t2pFOvZfVGNi+AZa42rpxSyxOy1T6pCMn9lwC/YX8/D3lLLq4bc8QeA5qM6T
phwbjA5QtBalitq89KyJiW+FHbrX8twMkJIq+tSPEXWEbSVpSGIWH305ZaRXNenhR+aYfKAZLVh+
UjnAAthd/nZnB3NVLXUQCYj3sHJH5j/ggN90oZmJzlCbSRqrw+ZuTZO1IXtniqE3w3er620QBu7j
E9eCA4NvgUWuLvhb74MSiW6FqJSiy6rNLnL0iRbxKqviEv+nWin1GAaX1ExgpsUs/dhPr54At506
n6+kTWpdQOYX1OBMUdbH9oMOLXo9b/g5FniIXAlUCMXxB0MhDfCEzE6+iXSo3rZwA6uJ4+SqUisY
rxRWsqk+W12lKbv1KZc7+hXz7QLfCZaml+KW+m0socE8iASYy5N+pgqCP321Sk0aCBBnjxZq2Q9R
Lurxn+qSk+hPW0xTYyLj0K7DD7blFIABErg59kA8YtqxZnWPQFknk2jylewZXk2qpSfQ7+fB9jCM
+7zK5/Tjr2/MLBQ3gpy5skXYcgiNVo8XCGURqAJkyq2uOZCEJyiIq7an2m+xTb030jfXdeoLq9gb
wR5Zg7I73V8NkwTvvZEGIcnQeSeex6fm0kIAISFNrtQaHVNVdX0phSoIC5kANcjbceKn2Sv3wvxN
vWl8WeZ4wyunL0jhqRdU6ZbM//BJQnzWmqum0nDphHHWv0dPyWLg4JC1AQhaJU/51pj2gC20J6eJ
DGfrbqYym6xLvRtAuubd7eaYboqtybyY/SlF0yMA2Ei6ALM2Qn8LZqYrmO98uZGVBoGwhY/kpJA1
L6njQvqPxtLrcsYiVVEytl71MWhiupBej9hbu5rZm1dn0Vojsik3qbk7b2u4oxeRlhKGC1ovOj9h
v7AJ51WZSa0HKR7cDQjhSyvs1yvE2ZtRqZwHNK2JiLcD3yOK+pg9laSt52t5tfdUVWouanmFOvT6
A7YPiuk1lYBBdvwFez9tDR1NMFMQGsZPmmDmwI12XwcaEHVAWahOIpnRilzDCA1nTPqTtt9G8zvC
+ikXa8jaGp2GQbCOw2gkfxEmrbfhgCIdFAAU4p94gyg9+Ux8JnLHWFCTQXRVijUlIydYqT9W7m5o
55f6Whw/mCcFh49TAN/JAeMx/CIke4KOJNYQFeZ58LVwlLt7MrBk98/bKKVyDdssB6IfbN5VnnOo
lfkpAV+w5XLwOOlA9i+wzf/hKvl+pR+RlI/wT7DKakJ0cNSgHNaIbjGu0XVIhl/BdowuCVXLopM1
WtDX4qV8QQGfU8KDs3NHGRvEgeSjLHiBjEhG0FZp0KB4gNYp4fUnkN0jcoWhg4SLg21x7QAlkYcf
BWmqw0y9S2+V4uFSqsBUz824UtrVcFRgPhi4Zd35At5z3cLajM3cirwxp0cwQLHuPGpQ357tKNpi
50I5ooDa1aQrTskx4K4EjvE4dJmHJToa8l5LhSJHcgx5HowC2M3I3389+WjVF1W20imBXWDPO0E0
360yJD2qaqArsjTRgmR5AEnl0v0CE5x+FHQLjRXWVsby7G2BT1V95O8h4koKVvNSh0YmhrdEpz+W
3mMjuPHE6hEpmfbmvPo1DPH7p1NjMIlrEsde3ABU1u32DS0k9mtvAGx6m6aXKFo0XvAp5QkeFjg7
pAXJFQPkiDWGPYW0aN/+RyMR8xzbTefrcKcxUelQ2i/QwfVMTu1nUVY/iVjCmwhda5VF7ECtbTAs
dvJsVmaRO0raM3RhsWSTSNg9BHiW0ZUiv1uWtWhkLLBWPbEhB8K6Ax/VXcunxxWWTPqkfKweybiU
mqmXgY4EBBy6CXo0lTYyhux9CYJgA/hWTriLWndUlj3v0S/5jXdJghjD8q9V7gu5vbDqmW4Favgx
7iW62ncM01zuFWfKkiyOwL84BA3M4e6B0s2YbTwIU0eia7c4SFHlJqZ/owrAcwxOQfQ/q9EJ8q9w
QpQwvlry8Ce9JimeSNVYaLEdTJVjUdU39Ff9RR9Gike94ah7cL/r0R1mQEeeYekMnaSZzTudyEJP
Kx8DPgrIq6zazPJJBHDKfa4AX6sVVNijRYRxLEopNZkbsaJZ0LsiGIvHIUJcX0h5OxWJ/5ffHvAo
Ry7u4izIFUov0b/p5pDGFPGyv/EBVI0DxVLoqdbeW0kCkltc3pvNizN06JrZPdqP5s1kndA0CPi4
oQ9eEAJ9sY3F+M6KEicG6AVylQLu5p750NofPviLACPd6JvqLD7GyBcnV7XwaAqEo2ru2Fr8RSy5
gBq/8BRPtmpgtpFy5vdi+2aohM7OhkGlqIYin3Rn3bRUT0ibNdsu/VVk47Kk+VOTt3Odt5d0KwQI
05Zj9Sl7WP6nYe1yBA0qhq3AaF1kYGfMp4HG27kwNcZrLd1SnoYO0Q2WrlN0vyqBimBi1t/t/VPS
Yi+tJzbwCx/WbV6iS9FQsU5jJsiTjHvJL/aVMBlGU0sfzppNj5oFvzikwy4VaAC99Z6MQZKCvLKR
VXlEuW6BRLw5VKj1by+QZzId9W1UEG687BSsLm7j4rPBIW4wm2ZZqXufD47uzQmRZ3bj/cXw1WBT
Oj7v1ue7u4Im0XkuWrk4vMbqd3OsaA5C5YYo12ELMTyOWmk4pNGxoq/5vJIUzg0IAV0xkDcGjLI3
41hopodQvhu/TTTr2X6oLUAugKlVvyPbNZv6FkEglqCOsiXyNbYiNbaEbKZxHI9yLjdiRirEPibr
NBgGYG6YFNtFQXDBCpj1YoDMu5ApOXbsqxfYPfexV1TWaRtnLpfht7HiNOstkCSOm4siQg0oQ0/1
+R3UGEc4OQfpe7556UqN84DQs1HpLXZw25+1SV3olbjAcxh1AwPZ2qghqxq4DuixOVZtvF3FL8JI
cn4SQsTA6H4002eamOZJJ16+D1hiegOMKbMHi5m28/skrXxmN3qdB6orWjIg/ZnS9937hSqFyGSl
4USYI2IXeOh+IRU9e+yJKxDrqi09iV2bfuyRr2vnI2aK22irhL7K1jZCsQkqTkFRpBV4iShgl5+T
Sbbm/MpqySjWvlzDV92k5jZDxRb/Qhh20psltOoWW49Su9JipYeGOpbG+i6WxkfrNIbmJkOnKw4K
JiRQfGrheNd4AEYzlDMQrFxpX1DvvAJYOT87mvKSmroHJc/HPKx98ZdJyHuTdyK0K5PY7/QhKCku
Tqkzd4khFU/6eu0kPNaIXi29XDR4otONkQqaptPPPmIDbvWL94kzYqvpdqLYoRjOv4c/pqwh5fLg
QH5xlw9z5Z6b5i+qMT4DdTQYkeXaOPpwtQ8Txp+h65NllhRXhFW9UM7XPTi34yXNBfeKcUnhNtTy
MVcIs8MTDvj3zDDKGoK5fA01EKZgGFGD8qLJy68fNkBkFhiHZx8NFlYFJ/bNneLPJfIRONGHlgfT
XCFOXoEHU8NOG7NJCaDndhkqeBcaHwwsB3duKOdU2Tz23bLXqMtCdFrj5Ni+20xbs2EYlXcHcqA2
jmFiZ+Y0V46rNOxKtuEONlMcq7ziTV86jtQf6Do2z+pcjwZ0l96sKCqbIzoEUigmXXVrLA2+II34
eFya9DNoNoEssCYz5jqUXZJzpqBHDJ2Vz1kKrU79Elv9qeuR5U88FmuQOk/EQKs0bjbWuBJhPoiN
giEsyht8XT8xQjlTjfL3tX/Ln/wk5/543V+GGC8A1wjF+vK2yIRJ4hJ1XLIZgDO87sMq/theokW7
C9XDU4fzrNUEG3sbv4iv5a2UjPWR50MOhh2t71otcw1CvdQ5tSX0dPCWWEDx2O5yqLyPFMXpFpbu
NXYJyOQCYajiQ6ypkW2HSPO1Cm7+8xIBFO/JcQn4Pw+knifSh5UArWcRbw+UQDwJN3A+xj1Dt/b+
EvXSJtlZ8gY7aD/gb36rUOH/eB6FtJLqSaX3szyKQWwGGkEIDn05bRDiUtFD87DRMQSZWNXdCC83
/RDqdufrS8m30UE60ZJHYm5N4F6UrhcGUI7OWq1Dtc1w1O46gF9o79sna+EA2CEP8Ud37LwOchbL
A78C9TG0vOKupjIC1YO6z5SWrP3TAH2Un3WFbQ8/g3qPJVGpNB76wwx0pRzWm7x4eLCumCZsoz/i
w9C4c46a6ug9Sx8GTUPK/N9w0NrgqFI7kg2iNwUwu67Izx3vmFXYRq8XNMnumjNBzw5pva0cXcaq
uhGKOfgs9XRwYmo5a0ny+AJQ1VymHKejKbdAZITfjg5wFDsevlABX0OjYQG++bbIPx1vmWbJWr9k
EJq1JPz/RylxRELNli2MDwIZtQUioF1+vgSuz6bndhjVT9kb2o6IqCWocI20WcddXv+xAoTEC6pm
L0/boeIbN6/0F2swOdNJcZHwEkxP6IQqxqw7L0vpMW0EfveBeAYUsmwEJhed5d+zRTmkjCyb5etT
L6rDht41NGhgcLxzGnr5nLkTWkTTy2YIkGXYsmr23/rmabfLJm7of30t957ncgEBYbiGYE8zMo6F
9GrCaWAmFJX7Yfxwc8KMnzjkQMP+WUEzmCZyC4OONQAdoPT0393Ylbo/gI0G9BH++zn6Ux5nxSm7
7eyWco79xTjKNsdxFOuudhPvo+oXcYFp7aGFqKO0aCJ4XniYI5u44B96vOBaxzM81IYcOgSYXVQh
CMhFz85EKADrQdiD1+fOjyk4If0GGGaDhyuUrBp+aYQieKyH36EwD54mECGAgOTCDyOJMF2BU5Rr
tNGoeRH8M1DWmyathwx7o8iaTAIsHUKTAQZ1pHg9/F4zgOT+wrDL/LgUy1DMdKUvXvc+OMd/zreS
S94cSEPA5WixH+pBvdbCvScHNfPIZbeR72HKqpP0FlIEXJsQJZpbMHCLksC/eq6mjmvWvQ/lHAig
dSmHtiL+UrfUz9HqMH4lfT7cfuRJj1a7Lxuk3+XrFAl4aCGIibiKDsDAlUDExmKwKbUKyOLC5/BO
7BT1KHFuWfYYpsG5KmILUX4q+k0r6aO8ByQjIbeHKwdHAEIhf60OiRoomy36GM5BwWiYKVHtdzPU
xQpLPlsP+RklAhJJ09wj3foY3XphjIo/MXnVuEq4CrvsKJcNcwkQp0t50mRZcfRAYQJM8qemOQCw
2JJfz1BuT+lAils2IKENwVX9jQWTwRrbCRvmHVY8Lxz4o38J9Z6DJSjEvr2rYVYRZWB8v9DnbZGF
m7IX4Er202QAvOWAFztIP31y3+s0jd+av3SaqFgVuoCFALL2DQsf8UOD4ar72WtrfJthRAsLEKxG
oS6Q77kRaFTYX8NgnlADDLGj45dY7WbRUeuOekNJnGqOEXPTCvQ9KE2sL+bEJCrhlcvNTHg12lyN
pNvv88zmL/XQgGsNPbuuRT+LUA4IL0+5xsMC4kN6mx6zGExeaR99TKbx9/NAFCJCJsLPhFIl94fK
OM02vRqKwryjihDxTdYmDbJ++TPcRkLgFxwLlF7zZMXVIUIG7Cy0RmroB8KjOdeMbESG2SRF320Z
6rKGFP7wBDuH7qYdPB4wfZCy+BVoTUsq+wIqd0Heu36uJm80v0c6gSeltOKQxtsBAoyC7RQMd11+
B6TYVUfkIuLO6Fc6izVg7ng8rDi3Kzpd1F1kQx5xMekZtquCX7IqzA23zNmm4pKzCVA3fFP4NJxX
n/aFhN/qgxe+SZay8cz+ofhk7jiYDnhkYQKYArDP1SsLMUoV3pqUNH8XxsQp1bnuPMG0Gi4inQSh
MmT6QQ9zxz8yQ4LNRXDi5kuo5Z+yWcF4DQS9/zSukYhja0QcqPL+XMS3ihpL+UKtC4TfVxEjFlH0
kywkSbCq5za1C2qENN22enQ1pCI6wWJ5oXOQh3mrDatuL3Ug5JUs8QNRStZ1Ev4/YkfCA71xz/i6
HeDkEbUXkCuUR3+pqBmGYhl2kb9uOYy6slyzU0pJa+jWCHMZuToGhFj2haiHeLQ9Auis8qwrmupU
fki2YWQp7vCjjsbc+tAz+spWHkiAwEuP4mxq84DXQHEsT9KeVIWQlCV+4F/cUnAVobbD0V7dgGSU
EGhaFUiDfLDpL4OezIbv8rRHndLxHiHFHvXHywHoEN8ZQGr8yCu/lQ78itkxsRF3IDUVMmchTZGZ
c4fugVfX/wNc/mxXcbBc9K8ywqU34F9o/HcfZd5rqrCCYcrT/TaizfxhWDn+9KnQ+die6Jo+bLzG
P9/8CCGGkNC4m1zG6Tfbeepj77zm4oOOP3SqRrC3NyQmvUc8lzVfAmCitXddnCGsDbc5vD0T/I0Q
QVRLD2tIe4U1ukAMimjMsS5IhpA9CcSOvTEcZ6GcDQIgfwYJSeMXNuyGwRXth5nhy0e5i4W4nVcU
LBEO2GrtoAAdmHwjdK+dR2FbKGlkm77OyQ3AEnRnVIGHznhcHiHjdUT0/worcASQH9yzk+23cR9k
Qz6qTtvDFR8PF/9sQG9JxTE2P+qarGIEBvKadqH2WRmGB8Pcof97Jdr+QCiRQ6CPuTSj+eWNTQUN
R5j0zfRi6GPGwhOtSmjaiPWvcgvT954wah/wRa0t4LwSUUuLTjl8B4LW83e6C92RW3XHMf8jxjuN
yBXOCBP8arddDXOzKKH2zCEQQ8021Up4Kz5J0sP26Jx1wzZMy17y3fdDsGYawkZbTSskKqcm4UYo
rNvTODa/uX2Jx8aA67AV61aTDF+fyzS2HhWpdmZTFGiu7+P27Usd7Oc19YaHh6X5wWsHeM8IWJqJ
yRf/s2JhmXOMZIlBfCs8fQ9FzY/f56wqkBvLdUv0TJsOQ/JXYqb2p5+4L8oErQmImZpIihmUHwWj
maHONA8kXcQrkeYAqI4ntNuDSnVcuakyNqBV0teFaUqhwtlEHZNW2btLMhIBlMSoTCJqHX0KkhZp
EfR/iXGhVZnwSNTLAu/hyajrVdOVVbNwnbCcVG32orrGH98DiDX0vQAQaihPSf5xaGgPAj7YSVcN
ehWVGMt8af85hyMjzsgh+s9INgwzHkZUhbiI9e+sRBz/GayMTO7B+sDn66AsSuQm2Gg2AVlhSEDb
Jw4tWr+XzNqtDzcjrBeeqx7XA5iTRGTUbbI9iQ6U4QYwan5nod1mKxR9DGHeLJZy6f6Wry+mpqXk
YSNFn3b/B3zjBqWOM4K7wIDvEIPkfgbVsdgMsNfjnAJSJTgeHrQlKY49lUj3z4tbz9BHkZtNtOk3
/qJTIOXJtSpqLXNhqfFIov0jy5OgaG9dqky6nz+p8yDELp0ZSw8c5tCnn2NtpiW15Bcv1kIUwO3Y
atio5+PD51Y4pHaxyQSf5OOFVZ/XSxr+r3sR8YfFFDc2iMLmFa7Wq4psB6KmCJIjCXChyFZ/CAhe
tnd8AgATHs1/OhzZkhQLcXp9YHRK/TBtooFHoSbULGynW6zzxnKbsVy6j7cgpgLdx49FivOqt8aT
D+VH6vUy+EO+5DjVY4e2XkEsHH//xzqkwtL+ypkudzT4pPucTqo1TczZqIoSbP+8QSWYqxdy8Ay/
2cPfbBjR9MP6fY7i7dahKZ/v42MuH03uMoHyEM4319SMore0nP3kLvH8VimKrLuSyppp11j3Eowa
TiM2/iYLP3dT+0PWSANzPiRh5YspHo75vJQRJoz43oMPAGmvQaB+q7evyCjfDyGV6UiLu/C6bjX0
+qezUu9MOIhqPDF7Q1cdBYCBYEQfPtiMwdgAXO750bUvRoA32sLTHkeojIhEOktQigR113nk3B3s
NTpMEcrD/TIi/T5VCYV5Yna13gJKlKiW0WQatJvxn8voe8iuCDgfQkvtv1f3ineamDQhIV1aTC2C
GzOi2YSfP8LekgtQVQ2MPnHW+3vCe/TiTfH1ny+IE5XT7dEDHLRi9NQuN3rI3c/wa1YYEbl3SMal
uuI6Nsu8ebE2TTLLHc2f9ZgQ6+XImcLJ9HxLMZLYMKwNZOE89iM1wj529e/ALgwO57SxVxjRVBxF
OyNvVbrwcBD2jORDxGnaHsmWT3mcYz2sYh7OAxlpWj8GOn5KQO/XKmybjjwOjq4Jw7nnL39vNNtE
PaWQOVEN20QwuMgQwotG6Ou9fMZB5Pt7VLZL+DTNyppy5TBL7qg3Nwo08vUIyk6GZwLSt5/qPhjP
tyknpAx3kwzCmSkbRCUJyQCmw6rBD+0R1OYE6pWy/t6ZJ3YM3FDw6twpkZwUs7YheLG157O9WuvA
WNYdOVtzKhrnOsveggD0+oFDKrv2ig6mL9qKydaXpz8++yOzq6F9IlM90uDkQjEWJX5ivaTfAi9/
9uduh+qDRt/binyMjMW9UfM7ccaj+TxNxOTItcL9XuIdHft0414EqyXVECTotZ/F4AjHtyQuFJtJ
d3SkAefb67fcY4YJCEr2q7p40hCHGFXCzEFFwOAAfsLn9I8t0nQ0sr7AEXH0aLFWY4sZm33a456R
U19WE5WswJ65L20XMipwaLDVGjJCJW+wcCG3sZPh+dyqI1VKbvHPh1wf5xdbpJnxwnsEDDB+ofsE
6AuJ0Hks4YEVXlsHDlmWs57W+/jde8Ru/6jE7TUIQv0HkkU95jv7qLz0iYR6ti6ptAbAX3WloFi+
4ru+VOnzt6YD7YmaijDHFjx9yLK/GPjgvN01amIR70c1pp2mNZLhXFhJpaETXmYlCSOUm9QTCaLb
M/qrH5BScruPm7xcMpGsU0v0YciggUNWRa0vx9ozL1+/Ku+AZHcUgVfGtiy7mXd4Km8yWw5oo83p
YGvYRDzSpeoH+H5ScMG0PYSznUvHtullsjklUMc+aQGmoJ7IebWQBlhFibA1eIaOycOQCnheNKEs
Z7CPCWjqlBenSD6ovzkhnMkrIvY+hCRENv5f33nhM0t6+5AHjs4Gs38cZKjGYQYhwK9YEXy9LXuC
hGfs0gKNQ+3rq5ZEPCypXK3KRYX3P9dm6cyvUrgTl3b8RDlwK23OH1H1c4pIjlzt18GQeLNDKXku
2THYGjPaiu/EcFlM/oO1j6WxXnhQx6NtWdfwrpI4mUp44CcM06/Onikoer77P0rPQav/7vL0+A77
ogAmu4tWIXACeUynhmW0y2zmYb0Z52T/mHQm5kwFjO99rIaxI5yD1QvxdHNOOm7Tard5s/3S6As4
5/llpUoEv6pGnqVuz0+8vCj1sABGapu94+/c3/2E6DjqnLxsOvYTiWCm5qpzRpxV9ynR0efleZS2
TrxshxWnd3iwQ9U2X2pYjhHNPcinV9FakmMXPHLCEkI3ymE2ghEVIetBr8xjRk2sj4hZrFj4SJxu
0OLuDh4Zl+dwgz4NpwZ6J/WcsjLRe3YczgqAivt3lNk9bljls1ZSJJD7FkjsKCGOjIrw79ZiVtj9
MaoRLub3F4yK2AGG/tGZ6Y4KQ/RH+L+npTGdVteh2mp9NIyAADUEVZWvyepF6rRhybufbt7PJC3y
g8q0nqqamyTnW0CiajhBWh8qUtZ6MqMPq+40Rd3Y7UCT4CT+wnTFueKOiRTvJbddPsQF8gvQFehi
cN8UCHxcH65n0bv1X6mGpyoS4hQy7zqPjrXLJcwIH+bc0E3o7vfrl40T4GOdtxX3eenmo06kHg51
+c+krRE3cKe9JN/9UVWA4WurN5itJStumhsuOsCDmLceKsGto4XS1lJp6dKNdawPFYjX4qwPewvQ
YEI0cvcUgv5caOeJgT1sptS9w3cwbBzyjPZTanYjMw0UntcB6ESYFSkIHSUtj8dxNSuWnlvq899x
3QfsJPv83UX7IqVGpFnJ3HFs12qt0T+HFnjkho9vpoLcrhA82m3c5p5XkdLAM5dPtVINBkQoXcXk
QRh5w5q4IyhO6aivXwNwAKgMXh0xoV2XQsKZ+qJnQX+0FBfp5wGkSUWMXhKCEvidxksQhX89s7nZ
JdhCdXs4uis4Xt/gTi4rLD8rJKi7G2Wg0dcjd5w4NFdl0zlqdEwsmqa7Yo9UAcII6tKbjWvzh/Q1
DktNSWuXL/O20YvMn374lwv+yP2pUTTEt92MVzbz2xLPRsbE9e2WPjfUeCijaAjBv0wmnSuZfvFD
tF12nsBZk+aMwf/V0ZEtpgdskml98jw3U/bRh2NBxm/BQ1ZR7GS0Skj9ftD7tjQStogPdAv3nii7
3fTjsZ8ldxeMsI1WDn9wEE3mHi1ulO8LfFDifoaLWrLuC94uNCefHaOGTgYnWbMKtZ/zUM+QUUMB
pnNf058P75NPYwhwxIg0+p8p4DyENh9wn2XEhIumspcZnEab7960izDkrmgUb6kjtOWETsM8wllu
FTty321FZ+R8jQzrKc72kowx/XfW+4Y0gONIJNFzMVRpK9eZ9RbxrRO253UOGg5Gg+DGOC0QaUpB
uEzRbMxaSL328RBkZHwQJk0aYDhmMmkocR2WU4Up25A7GsoxMWtisfhewJB35039ERmgdj983JHv
9ppw64V5YUym4u0VAsn2blhozWW8JKzez2MJVk8CqRAXSauLOMSA7mFug7h/xIAE7ttyYrIJzy5/
9R8G/dz2zaRl+tKRlNxux/fhCrcsnsxVFTPepiUlPXw11qu+ugjJWajwstjapeiAGd/9w9vCQYRB
vwv6+TXi1AFt44cFaEFYdQGbZWj3RJ9Sqe8yL5be5zw+m7MGoTJa3JM6sTtXKsj+iVpKhtw/chAK
/0f2KNePPxaVE8VPt/rHcIeWxvTd7cR4EtT0fNEeHDhtX+cH8WkSO+RYAtPpKshps8MFBb7iwM/S
g3uObSDORbQ78WV3YGpxnz8HUQ8hyeJENaqUN/917lb/9RRq4HqCsyA8q6ES1KmTrRyC/jqM0OX+
57zrXDTg6cA98/IhRXJfebnIo0WKeU2+kiOcppbx/K7co5W327ZvfGXsSBhLN/5COr5vMTSAAB0U
me1O39IOtaX/hEBTgMy2MvrUFb1FdYV6GuVFzBO7pNm5H/fDo1tuN9uaWclSqA5R/d85ss10zNy7
4PDC2EG6742gPPbeZb/OEfehoATAb1zm45ubSs27u9ypNVAYu81uh4cEV56WDNl7U+8+HpJuhEhy
/X7hbTMi6ndO+5WSkpBq8ojGk6C0SJ3D8UnVfGiZZfWnBaoCymuJ1iUwFYGy8d2zhSt/xPuwTZfL
75fjPXwiq/KC6/6s+wA6AUWdRPfKJjid3CDjQh4ULAXPpV9X7e/DCcx2gwFFMBZKi99I64rmU7+Y
pLEpObSAMU+WCjkoVmBGs9cm6xd8FPpGAI4n721xntIyhxdOGvYANIj7QCqp2rg0rZbgcNz0B79j
9WbStEsExYNxAfSJMRoZMAhVqFPqea0PtcjSnNPSyJvnIV2zM8ZLTnUIEYlmucSBwiKaqjPImo9z
FnLEayuGJHfeIjsrvIiJ4ca0dQABJ/2nOTQRo8pHt59G3xsCe55HedRbHAzU4uv059MeD80as/a+
5ZgOcQu2ekkujND6YpgHRQUjGOuF1SQ6EZIcyn5x8nFigiC1bwjsy+OlsX50Dt834hkNiPq0Srtj
grCT8lCGo7vPBa/zbdESGsKu46oA2d7BoH/QFsHs4XVb2mVegkuIAr3JH+IIZb0p/41LXspIQ9Xl
X2WHSZk6hc27lPF+5Jcbrhm9bZ2HLPC833nBTYpK9Dz1WWOpLcMt+UdeIPyAMwFypNCkb2m5Buqf
dLyOXndnBoxCAShGYIiZcjld7E1C69y+3kCMT3xFdKAVnTaDDCpQLD8Qz/KKGPoEG2j9KdRYThc8
W5rcFO+5Y16kxmJhTjuIfmNLYWPMAlnthNpCHv0hKJZxAMBkWrmevhQy2iQF9y9ikp0s9wNMq4QQ
1Qx66o0iucTmSfIZH5tDW71pFDQo9EZzPzqOOEKkRvj+42tFSDvFgnQqYBVVIOTUU8g3Ik0Xb8kn
NomSPBtv0yJVBin4HNfuo+DtexWjo6s6bjOPxw8MHKm6pSCPlQi8tup4FtcgWdISNvu6K7oUwJGu
Y189nFKWHpg6fknbE0FvlTvvI+pdMw2l69ZjUhHPHArYW9fxRlCG0J5/38keVN/LAQHb9gl+sC6z
3EU6FuaQISEFt1x2Ob1nmI3dro/4241Mub02FSuyYVFYQEJTSJi+p99CBErF9QhAeA8MTdaBbFm9
R2NFVD+v3DOdZb+RTQno+q1AfG8Wl2HRClvXxOxBRyC3t08Gsg0taYlt9kRx8D8dUUcuazyp01IF
sizmKJX8OdSv3K5bWKX/N+0yb6y/c6JigC238mhqDjIPWL3Pl1rptIrpFIfRPKC38CYJ2WecJDGI
Zyf1NUR5BQQsvIGevZc58JL78WrU8MZ/WCdkux2+RfCRlyIpeRMbvnrko876gwWvJfJHSJAw6ARd
1oTPZgdMxBn/dafv8t3nZ3Ad+mV+APKo4Q+ttu7mokCRB+Ecgai9goCgXf5Az2l9F9IBQu5cCMyu
Zegux1SU8XAVgLWqlgiLjZVEc8R4F6pUWY8fdjIwgosaffYBakY9h35YBWbFIx3j6Yu4EWPFDCpH
148PyiR5NEeD7eYcjfT88qDpQ/BW9rS4MyCV+6CB2ICMoIPyJLzxKwFgzdrArh8xNIhsJkcIhRpr
t+/YTun4bV3uBbyeu9d7qNivSmQ1I9O8M+ri379zLqBzasj5+HLUcDmrbG2g2arYN6CODgh/MaVC
702Lj6cA/QdUJoQv5TUd0YkcM4PjbyGvAvVYw+0g2GIwFU/8NhmLhksvN4vE1W4+d1bVOruzH/9W
ec4UZ5Di3Os+8U5MSc0dDKBrugej5piJPrxvmykR6xHvGHQOVKf14D8PdGlhi2tOytnfgYePGObq
1R0XCZOg7VQniZ7ptdmdVGB4E7TSmvk3mS+IaGd8uoyBnn3PcrlUtO/xF+e97rA9Cw425aam5kvb
LeKdGkxCAQRdjhJ1ARJezOS1x39fQ+Gz4aS34sjP9ax7gO2lwRS92E+2kDby605gpP8wmpBBwU2n
kvjGreY2z2LKjzcnX45lLVnD5lNUIEmL7VzW1cA2uICb7mHpdBWgJjPV/N8MZ8uUjMFtVtsTBvxB
0foD2NhwhazGT+FfWKKKWqKFSbkKYYknv+aDeAkcVD9+EsOAfQfinDpZQLkaW3y41VtS68K8LbMf
9ySH4vjNTfDXu5fqTI8+Cy76tdV/R72sf/BMLlcNtWozn31e8kaHzv7WcP54cFZPT2oh0MttoCF2
xGHTRvF659mc25hywUo8LjYJwDkoKZCen6rkCJ80qxnIAZuIyQfl1DVgrzFn2ttNZe+uw+wjm6qv
Le2N8hd2qaLGwPwTaoHKL9bNiuekcVrzOquzG0tjr7f1h9HOknqNMb2ZWq9h+0xA1J33Q6cb3uOY
g318SqzZBweKZnQZNV/ksb7DkQDHKBnaNcdgFNtnIjP0TIbNPxqMsvghjEdhs/pPDXPOFOOvxulx
u5EQ4iUS6Bn9Yqu6VlL4vdueaRyk16Ro496e6xHNl/nEWRXvcY+9tnJFsK8fFl+NzHh1kczaXRi0
BtfLybLYPkHFyAqVUq7BmaLh4s7WTVKM9Flagt1gf1YXx281sFbLK/GnUtT/qMMFGbSLfKdSI05K
lXRrOIYS2I8MktvU4YxOGjZgLmBOZAhvGDCE5mn/oorQ+pP8ncTdbFAC+K/LVJdCaO9Gt3tTTMEU
TCjj0k/qr4U/mEGZs6Kbl/4vtun1FR+zzFnAx6IRzS6PtIiRbqKW7oNTuQn3GTxCRzj1UaGpiQFS
RxZlsNdE+pdFd3u211kZwoOSDdy+wE1uf+XM7twNEuMVtAVLRbujuQXhWsfm8fOyEQziiaeRmqMh
XSPsBtsXXf4kpMlRSR1KkmPOIBWTIOBbCqB9YAehc5+0RvFfolRQFCzf6U9wu9/MM/kWzhtCEp1E
QvCr1z/uaahW/5yDiTlJGAPq8d48qPJPJjVx0zvLdAiGKUBIVQBkZZeHAPfc9ffSb3/yt11Dwkj4
joxREdJIxbIAuIaeoLRPyRAswVEaPefoBTGUCU7RFoY624BF+Dsc32/Wupg98I5DFbvvuqOge6RM
nAIaKxFfJgmmbrH9v9t8uotqqn3u3770t00pLKlfRPOWvFMD1zw6BGZJcnI2tXIrJUzP2mCoUnwK
ihpHv9MSYsWtIoDoGXMq8isxCj0omoMWkOrQcI9TnRvpEioyHHIhXp9hMYeCAFxyJGY1wlAtpick
XFi7a7ysdJrInRARWmshGjI4lQd9xCuyABKJELrY94cMgdqGuuqly9YVRPnKa0s2+BujcY0SU6sP
FASwRgr5fW8SYsRvh1xW3bboAkWK0liufIkgd5ph5xk3P8fygm6KFDNkZb1cQbdjpbn8+64YFv9t
TvvRYRRi6YRIFJKctWKP47eT5WC8Oy93xIhoQm4Sr1OQdaipzTVKrfz9JMH9Fjg9oJaNi4t2dY5h
UPja0OZqowRv0Kf6zuQ4LdZYH6Frri2Z9c9WAKDhNohyfHJnm7doE/rI0TCrrdvZ3Sc3ku8KaCYd
k94gNC9Hg5GlWT0nruhQy3kwOfHENXkNJ257L+BNuWzMnho6QWH7a99mrolmuA3TIqyWDqiuWqHs
wZbR2DhFnydb6Ypww0OCFkm7I/hdN6FNmlCDZzYA7E186atFxGseSn2poCzmcgER0lsIWIS3BENU
9S6Wezm47gCgDv6ku4nqLCbhLEhRBQ41AO/O0yozpsepMVg/ViNCq8PgXwoDkE4tNaaI6qfqCAcK
rm26WxHaJWvCxwLl07REvzOa60NE/opdkOhisQ3dpUKOSRLDarx/AihuFNXZ8axHvGTGEbQx7OVb
3E/nRhDF4ZDlgijq8p8oqeZagx6AWXTXt1vyGSlMfODtX6MdtGFB8FGBBV6ONLL8Rnxn4AqLE3+m
bZRtuUYNaZW8lSE7Ik93iI2HiJMEttIm3N0sz55EbKXGTOjcf9MNOQeoEvI+B4PHHG//iVCShU2P
g4jjJe8Ykpcv0ZGEwEN1wioXPpql1mudwJfsmSyOpmZuXXVYneBDyUQ2qKtERzv7Rb8vjOSVt3w1
IIu2xj8hxdm+WolK9uc1DO/VABIGU0h2bkjcOjLuJiDxKqTCxsPrckSk1ybitRbX1RNtANbCEscU
BqToatfo2wiR5nyCQ8VSgB7Pi5cOQPWybd/iH4bziX2W/EcSsqCXa7TCxcynVvpk0TkLEdcpvKWn
x9XQBKmaNoAuMmiqHs6ifJYkimtbjsSdHD+ThZZj/plAYyY47/GpF3uAdOK3bap2z6gbs5lowr1N
tFhsncz4cjmMUrAdvMGKdzyxV/EW1HiWdXSFFAMeY3F1fRkMAV1QbHzGm5HQmkWb173xN2M1wbDc
sJBHf6j8EjxrMQK1osDdm7Cijt+5bjpxXeWlRlJdEi9AYZvZC1lczLbPebMAToUmi3dgGqK+t5KV
cgcngl3/EhSQ93DqljQdE20gpGRFnl+MPdJ5BiKCc3Oy0F9Y/xLbwgraY/7RkpiejdcHMWJzDw4O
u3JKgeFQyJhmaDDbK4f4Ikwz2/Cb93NAgPsrv/EZnextpfUn3xocHipmdIsLQBSgzfG5r8im8Y/5
gvGenRcDG+U6laMBQAKjR/T6GEUtE/sYCNmZ1gAUxKxPf/UwDKgTe9zBcuJRewQFc9s3nJTueKMG
edMmrcXLDEXubINS/QlpjUDwKT2GdExgihsz/cK7/OSnsjku/CDGLDQE/GGLKsCKJPABElq9CCjH
cVuJF7Yhl8Rr8LwGAnZR10d460buRn7miTQM1tsitGBpWBppikszZaB5aX0r3aurVgJaDrUuliNG
ZBpQHg0EskktA0e2cA7KkONcVkMkujah4FumhDdLV+R4V66pvBqjuGJOQ+RSm1eSg/1tWUIdrlLS
KDx4DMNaWAvBKff3DV8CdaCKdB1Zx9kakZACAMn+cAo3K3cGCrM9tHoVLHoSUHbYys6K7YIw2KP8
R+tS10A5mX8NhfJyXzsM+dVzyDjXi05aplfzBiX5qannww6GjGQa6Qnrybt8PVWFSRMGKD4MceYA
0irECYWFkXPeUdUb2TqH+fXr1dbkvz/GhBYu/xlb8tMGIb79q+k4g5oNU2zguAs0XVhRUUZP0tGf
sxR0Mi6VhQkVEIdWJgKPXX1fWstyEf+rdZxBBdxxnuu5U6REp0cDiLqOcGT7u8TI42csFSQs3+Yg
FSL97xHVcjToYiSmHWBzAppLpgRmi3IA2b/gHWFEk2kzVl+RH2/F7kkZiAD/KrQ4bdCP67m1IQ8N
pLzkPi3USh9OjV/qYShlVKMqTTPaw+4jeAk3xxlklI91rLVgMXMe/6Ef08PHk+vRAPvs8U68v+59
oFLvkVkIIIWjns7T0BFLscuX0Bqba5I9esp6Iun33+2itOZf6qufK1W+XPBCBCsptOcO/Yf70n2V
BDrLAW0XUJ9hoetm9e7LXo+D/XWV8kqEO/eDhv7S6cvj8tLClCBqiuIPvOiGS4QGwbk07n05QQv5
G4z0C1J40q0aK6A0jpwmLaTwI8t5fGrS326/EOeiYegfpIBWkfGJ9Gp0qA6601935R7D5yITpCWG
qSeM7Yojstni+NqVbohcDBPOyFFc+9EOA4fpQSyLnXx9tRpqixoDl9UOC1/3xidatPz7K6kWzseN
BobKxVMuQufWJduFUVTo+WjDm5VT9Redo05Pvw2WErDVCuxWsjAn3/VZ0M98ATag1tfcME+Cg3gy
fElMtvFXc1XGKhlAe1c/ecRkPh1xEVgYIjAEPfcTCyLttTpf50kL/QHoyEwHTXQxTdGtU/82cirt
DC2R1fUseCa2t4WbF2TqPwKinCNh1dWI9JcdXChqq5XafG7Ap6FGjjqL68Mb/Z3+AVVnv/XL/PoO
DdHv0se2wT/LQsedOo27PsrMtT1K7kNMf5zxlcnRSF0+vZCDvV9+ejuxr9+GtdQhvNT4a/MlXrqT
eFwkHVYWhXqzkCG8xx8IUfN561+Z6e5s+ba3IW/vtIqNA+Bl8l+xRDfRgARU5cnAqwbmyyfkb1vk
Z1fZKzA4TMXROTyIlh+F8XNkw4bZ49tBGtHN5OC5auH18XQ1noZiFkyFLuyXVU57Ffa7twVG5rbQ
heq6/euZJAESnpuvV55Yp+369SxHVnkQ7BQftp6pVIRTpc5WQ+9WqoOoDJK0bYGZA3XWK2Ivku8t
HRyNnXRP43oyUp8//7cIz8RldyOqLxV+5B2Lx3xrPQ9VMi0BYuA83tRnvtY2I6haMW2yvISdTKJK
upVpgIMV6AEUQpxv+GxK6ee2HaiZ5LWPuZLqTpg2myZmTlRgmmu1At4eBuWFqp66XKSuYKp6Jry2
3YhgmlCB+mPq1xFY+2iGIMgu1LfT+/rVSsCSJEqhn/HDWV3OTyIn9XwSvnbiGJYw/Kq/Ap1QAiPn
/KihqnlOG34cB4LF/BOdoHReRcsqEalP30BmiLDIFyeg8pqLD7gAOE7caXta5FwJGzvAURwbtu60
v2tzktL8aK4iclnxDEIrISz96z4iJFGWShY5q5hRtzGiOszQPBWZP+neW2ZoZeT7ZFJrZ7NYH3jk
CXsnOOoJT+qsSZMhNzJxsp5FS61xQcET+Cw4tjjUIOjzT4Q8zCkv4Fh36qjr3u9Op71JrnhCJOtA
Cld7hEBqkxbRSyXwD1Aecn+kEkNRiBzybWQb8/l2WEM5tdKQaTMRP+CMOsexNvI9o+NwRY00cbZI
Yy9mHe9j39X3rLQchO98tlfIcXan2daqSkLOrWCXIKP63sFgZwZ8wpGV3lry7q3LTBa4CxoAtuWz
jZRqCzc7qv1J3hSf9ASW9e+mgjDr8lBiC3Ja06To07UeLUpzQZhy8AgGg1TWdiY9IUERB8ryt9ZA
PoxfHHmo6JGNB8S7jBZCYzqfE1aHD9Zz7+Nn2B7j35meN8bqgDy3k4mPx4eMuvUMsCwEVlE+9zz5
Q28CDm8t0pqxQSxS2YXF7OYbCMSfyrfQu8G+MQP+jRQB8H8Vb9G2i2QdNj6BZa5P8+svF5xA14Ea
75mqjaEuU2p1CyfSkuK+OOYnfXYVLLEv6FrTNUOcTZaDdorSEVaKTzi97ruKbC6rCxq1dFt2MXEJ
BzrjhgoZ2HayfeE6PBiEtIEU2Bo+3W4ayjqORck0vrl/QttLBh8bbhDWlwKfY1XxPCcFOOBULhX9
2rrcRoEzPhtICOtDmm28OSP3KFP9M1mGbZanLIlNGiClT+KI6yKbBzqwgD7aibVMBoOmLhmJEWLi
zCriDFD9qFTJ2a73QhuZQKJycVzZi7eT8rNSJ4dGzxrVJfA3HKKo+erVADH2xuQTJWzuBb8dfsrb
fCsI5ac3VETDiU+qiwe12mo/sJGNkK6OM47yX8UV+9vJEDDl4gILegJvmBHBxu2RV1rOL/0OPj0w
t+xBe3d++M/gutunuDrYw5ydlL6LAP7s4l13bg4cqoD+D3c/LfyaVTww8Kp0/642K5y5tE1Q1l2g
YaeDT05pyFf6rmRM641z37bD8zogUrlamLpJGckoU83VAAdCO4+DQ8fmP/FIEpiM7uYxI0VSUA7T
0wqndTfNhojFIeF7KYUPZpOfj1kmEWZugV13l+J5TWzM/Koaxnu7u4Ze+Q9NIf6HeSIb1Oc+QGuM
N7mHCCVWJyvIRehL2qj5sFxFhprm90LLpDniN8/QI84wBKkDWCDCpDu9vzDwVBTz5TEkNoeo798/
RJdGzQRmRYV4vOmt4aPyokHPxv3Fg95H+4rMsYa32pUt2l1yXOq0EaoureZfQAh+MqEZlZAFSLcP
bJfNxb110TM2+w588LY7BJrP2FENO+Bz/j/UIn1g7wWmr+XRO3Ry39ELXzBDDBN/YPvLs4i0KFVt
ii/AHbeSIpCrPv/Ww/btL8txK4opYXLB8BYX7e9xcMdzhi+/Wu0E5vZmQ6MUkixfA4qV4y83xSTD
G+2HFojgK4HTNn5EmBDYlql4IOIjqQcxyBik3ASO23YcTcIAgSLl+xkr8Od7uhKg3YXGstYIB5P4
IZgOH0CKeXsW/HC4CKHFT009X2yo9D4hcwh8JikLKysQZevBDzp0qh+DG+CbAxBI8c812CeAfk7e
yZh/wV7I277TiC3pJNZ6EzVLy3DUm3wItDY+xfaN2ssFe9QIAdpFP8Je/ftZX2UxvhacTvPlpgSq
sIWPLSMYbuSoBCmt9VE1R5dM4/amt4bkmQvi6VPEYWh7FFbbrgJPf4fpRZrwg48H0JqV0ePjY8C2
Bxtdj+utGGOWXNKtPNNS1PSOBsunukDRsZNseR9zCMJ4g+77baG14fY3nWwOz3EuFaDhFY9BhXHP
9+SiO3bYKG0YxYujWt3hr1QiyE9JgYoSRz/cWjtuMlyKdPVlOIOob4OooaYn4h1MI4rcN/vX6X0O
SuJVP0J6bBSn6G3N2rHyK+YbySFF9elMRb5hxkcI3EH+yARA9zyONBD29thYhLIbN24TnFPlO3wI
2eg/1C5xCxncP5+4YCO26Ki3GVYET1Ysc/VhVvmqySmFt0FWE5suIw2AnWQ0I3vZQBTQhjRCR78e
Fxk5hqJFXsuH3GBHwka1mTyKy1SWYgiX+PYIZR2LLxgHQOS+i90p9GNFeUFED0W3NucYnKT2YF68
79X2KsuHBQQydA5A4LcuickuYNmwlKyUjgfENrnFXc014knTGUrZBD8n3azbMd11qAjyJhbD1va4
M1TYQv6O90mOcNBjsf2aA+zBm00FeoKvbipc33sQ/sjN0aFM6Rr5Z1qFITU+YoNcIX7ZeA/u5Yux
pkjj896B4mFL2osYcDsww9dixzhwmqwLATwYiiSfKdDlnTHIZOeazOKEFMuOYlHU3kVj76nHklyQ
QfNSonIUIkSSLuiEZv4W7Ei+1YDImDS6NY50eLqpWXLzfcp4P0LnF0YS7tWW0y+Zn1/VPPDLI+zN
RjDkiP4/n8FmaV2HqJwsISWbWRBdGhZuEGN1bf4/RmfK2Vmju/ODi978TdN3g5+yXK56dQ6ikVuI
s9+76kiN5FbnNE7SNwcY9tI7ohE7itMgTvXcb5SMaDdjRxNTI9KdkVEKgUV/xU/VD/FRlo1NRheu
dEH2ys0fpf1gl8jbTzFhHEfIgT6kfNO+Eusw63F8dJY8RlKjwGIEHhIvJ+rKqZf1083yez6br10i
B1EeRxqNIyzUplXXtjjgQR6FY+NiD8rrBsvgkeO0xQkmMxZmtkYIgD11m5j0InuCUbwkZfCFDTXZ
OKu4SHjYiq3/4XJPHU80okCMp8elnheUKYGrSM3h1ZOUGTkffpoK8i19SJrBHWqxJvTFP+92mqCU
+ZR716reeEfftFEzcA2tAlSA9//WbabWuYCsxjyIhFf0C77rnouv0a7iL+PEwJfdmONf5gIPab2h
WIonMn0ieU2EdjgLpSi9N0KNxItMK7mv5MYite9dIvDEWWwU1tP8YUPC78HqrGr7cUI8mvPWZ173
4U+W/T6+TuXlo5Nf3dy41QGEP7pYwlEmm1CGZt2n09yxuS3gZ6cp00Q9Eo285GxOIANsd6oAAGUa
w5568ziYgNdaQ1ntG8a9NNyNnW2LhhN68VsAvECi/Xo49VdjxbW72D9lS+ZqWIEg7nQE7RMU6jlK
zQuS3IxV8CJE5+LfzbJ64xw9+0eqA7nqyFV3D6UnF1NVzznnNjLW+sfHvxxyIfa9R2bv5uMo5cZa
0xcRF/J8CyKh6pf138E7mJ3GxZnfZmuMTCR8IpRUNCdC/ZEzAieTlnpc6cURA87m+ZMCUD+WZec6
hsId5I/Dzd4TUnFEDllnxFU+/v8XfbEsgaixaHvoYlyEKJCkGHuzlX0THWVWV8lsJw5+x6S4B97V
pG50IcEaqpfo82cVIuxOWdj4e5mI24W3LWRMxBYU6W0ZDYMr3teIwakqKZP9I5MYHLNEVdkhpPOY
eAKIdCIjGZMq46cremK/vUYGgSZ5+kZsuHNNeXLrx7d628QdQVcK+NhBkqb1OKTJwI0lhGXBjGq6
yCGEM+IY0AulY/du9Fh68kTD1SSu6GuP/UdXZce6uzFLreb9TPLwNdVl9N1XFHGEq1DDr64d9G5s
cIQ6nirw7v9ytJRumcgi0zYEWF0mnAB53ohUXVHAeTn2seoYBMqG8bXZDIbLfuH1vBIrl5GvSIOU
aABWGmW1ZtDWaNkfvUzILjcQD1CBHtFT6SVcKLqShojCHbG7d4B4giuHurZYkg3P8iJkalywpwLa
jvaWA55eE5FHQGLQUVvpBorl3gaz2g5+kptQwVl5rodUM8DTIQZSbkKrSrUtLJaCNoDc8Xv1ZS0C
H10NzNdxbYWXiVDp8dg6CmDiOEh+F0nFTttE/jSBRskkM+nPB74QqgWKmXDpC2iyLZQmtTxm/naj
JGKsIPeZTIgl85AIOOrftY4g/R/8Yfi+w0xELOi/8ZDFCO+RzZgit4g92mrBudUmAdrQspwdX5zn
KbbZXX5TgI6rk1P12cqH6i5ZkejRNj8EStO6y8q67f+At/POLeI2RbxsZp2iN4eN8spbriK+0YkW
H5yiexymIr+UIG1NYNWa3Efqt6Gi1o/6GnQjPYzoaw8mlKFQVB/TZYGqFqiroj+u/5AF5i5wct/R
g/tfD3bEXt3hrFoxAy3axdtJb2HkoFxUlH3p9R/IJMz4Ek5N927F5DjFiqX2TvdFYGATGcCRJjN0
2hJlYWtLAYhEljZjpgGzJlmEFhmjuAGDvw7ud9ohDcLDGlQDrC8B8uJvzDi8SmWF1iFxc90zyZVe
K5LXlX25rUw607EQcMAOqZh1kp+ZhtgfUoGvYX4xZPT2kb0b8TVteDezdMrsD13l4aLtlRY9slNH
NpEkMmGqEG/sQaaL/MgZwNiASdntalXhat8BN+j0zxo88nJ8NKjL3O3bF8QyXKUK+SkksgRFZD/N
9n5v7FUReR1VQdMOaGCi2whjnasaX7xTRoxj9B08vQkItb5ywNZL6Sn1Op0Zfl8xdW4QlMNOlLV/
mm154Qhpe5hOJLkhRi17WHexTE/nv6N3/+bz4IWiGGCWP77ct5fXKrDJGl0bV1yZDNw5Rl2EFpZu
Xz1qhBq8BeZIGAQMv0ZiR2mDkc0LLs0gN96nGSLGcZusns3zPmcBzF9GaIPkjVzlXaQJGZJJrvmK
+5UMV/fuxXgn/MjT/Yd72J/J1m5w7xn38iAS3JY28h4GOgOnHNFj4P9IrZ4koa685avrftMXgd2a
wHhhVUcPzS1p78tD+9+a0b8arb2pYaeuiXyjJl5RGx5T395oua9xzVPBv1Fo3QRQWDhj9FB9FN5s
H6poPVrVMhNL/wkAppTHkUEzoANj77WPNi1d4WcQfgGkCZtZU/DOcpddLlMJzNYd2xqD6t6bmVpb
DiILzxB47+60kO/fRoScerVNjLW4iB9I61wEaQwXxZ9ubX/6GO5GsbsUM8g8tLDdxrzgM0a7qaXM
0IW6isDFqm1KIf3ST9PcPAerCA/04+JHrgVnGlDeVRdmbEmpLclGbpJ5X8YVEbpTs48vhE6VRmMs
Z7m3985V4zwXasvRezkPzT4f0K4tKzl6NLv6bFK3P3upOJ7IAU4KRTH8XCc7UIBk9wzSwxAsOyfV
nVPwUckfEu+Y8zG+bUqTZvc4JoD1Vydys8UD4kf2IDGupo8Q9wfbLsmQBOv6iaK9a4bI20eka9yu
D7o7sfWAJxr2V2l/xLEQpdg3SedTTQRTBnyYVX2vDtNr13s6s1Txihi2xhji4ttnQ1JeZEwq2g8M
4jqcfEHcriuTNYalMHSRx6f6WTfSFvz6+i975ME7OODxByBQoCPw8/MRBA3mDY5+ah7D7FAvGX64
vqsuwCsVMM18GPlTP3OawsmBK+2EiK+hvnHwu1vf5LUY/xnnGwtRaOEhz8Lgx0S+MGHULL//H5bb
vE5LuNe7YIdlnA7rBzGSGNBnSXXlRZS8neaQZd1Fut8ZgWsdxPrV7cIbbcpVDk3kNWYow9LEr3VL
rhVvZoUT+CXi1NZ/9EQC1MZDqF/meDQ6AQ+mybUADLhp8rZ0+L8Dt6Rj+2kaOU+HEYxqzymUODha
IgRy0A3NQ/4wypWFhwh59DRQGgIlyHtYZqX4QBwXS/gxa7XgpbyWXsegKs6I9Pylhc/GP7W/sd+g
wjhMpOx4RdeZvtwkjFsog+GSB957U1YHfxE4RkNDFdfFxz9dlwurq+6CXXuHM6x0lEzOaVzwrc62
HKmP9OFjFdGOVWogBiv5TUmJz29QaQLSoXqqPwnlVaIUQcV3D/+2hFBJBbTbGgIpAaNPrGan6xLN
5I3YI29GkF7xR0QPVoSzNLDdMhp08gIJD4myiqTBeNWm9XaxRGdknG43tSchEwzn11Qu0m1gvngw
/FZs33o1LAn7udQ+m/ec27erOJ5g2hEdOjXzWyNYfsJd6jDaftmvhaSRUQ5l6ZpsneZAd6dpVZoq
BQGFiYNvDhReTS7B8CEOWDXAIlJIA3rB3laqGkurVygL7bqBYYE1COhMbdPHL40ko4/XOaVMl4jH
FLqkgFbLWKiGfqRdnS+33SX7P+zUiXgJbqju5Z3vmm0QLslt242I/vI87xMWQfqUVb7rf6u5ovu8
sVXiezvG4J3uKFlTtLr/YDNNz3ouMlzCIe8EbjB6E22UshmSsBFerV8zpTDSVEQT9YR7VrmtfCv9
u12ODAbyHezdE2ZYOp3yhCFCm2gTcjfBHdjZOf2r1XI5sllgucdZEckjXjn5xgS0oDmrBWQW5HuB
Rkf3D+pL5oqeraEDlaKGCXEhy0TmazGDy4tQWRg+5T0u3P1ktdA4/NHYVl1FcV35s47t5NCO/vAK
0Z3JcR/+nsF+2bZ8sr1v1QlA7W4zyxnkJYJklM9mshqWn2S6aPPFmY+7SwDM9v5UX9iBv3zTmNm8
QdbDwtffXXjsiAYptthxAWIPjdEjaTdowLgodldUSuyQ8FYTF7LlG8uq+vqVPMxxqcUTNt4vRggT
yVCO4ipw6tvCzZLNVo3LW4eyJmOjqOS2RfvuMdsqRfOkBb6Hiyac0WaC60vheq9mmruvkjCZXc/x
xt7TLBSk3wE1NFI8ed8htvcdNPaMzd/4HFl+hxrPeR+sKx2P5SJbltTT8uAJPVx1XsuThz4P+/48
vioOhZIEfQIiSXnPlcE5geBdv8dkH/1cL2zlmX0ZYCb8XjDzIT13shhYX2MZXFCeQHDbTQJ49Fyb
sLTzzTVZx/9nfZZp+CYXu8tGdMNW153Vx1QMdiFvPmX3YN9yhA8JnXVweXmbpYbZsosxi8dMdW8Z
EYG8kcXiyBT9jNom9Ru4qXHWQe0R9fLezbD5tThh/TSb9pvPBAPp+RaEMvcKBK1QkwxzTYL0GX+Z
zTcHM14lcDZcVc0etF634dfrUCMJ0hotTmFbhMiL0ivfmKKMKAscfEzKvTSYwkCSM43tn0+0Cskg
Ln4JRgBlnme358gvaXdvojgMIFCOYURPhUh7hlEjQDpqTiqf0YR+6X0q2lC02aEXw0E+z/DInym/
2Z3DOJDoDpD9jor/gcPDFGb7B+Sd8MRolOg2ImGFDL26eEMyXAWtwcqtpvmFMQj6f9l4CHEXrb+f
hJtHHiroYwtBmKHf+nM81cMzqPqIqUwBtt0tdGAmisxmFFbv08UZy3kjlDXlWO8dkf+m/XxTLzIG
JxyRFcnYr68/goZdZio/q4fOOGzSNBL4kbZ9RewOV5C+fzRtZdWqhj/7B1zNTSpYRBuOesviKCyI
Vwc4P+WujpyMsy9x3s4IyeKba4DSpoR7hYKCA2u5kTG11atg7IxJwe31IiWqj6bnv5xQe3z1yKT3
wGM90h8r0k+Z9j7jKJfaum/lCv02nBACPNpiGsTbn1TddAaoJ0WkEROLcXWplIa8as3TLc+xGapw
OM0NgUQkmQtSp56Gg39oL7b7uNr2g9cgUXQjPtmJo+Ax2j0zzQ1XgJdI6C9Lb2A5yFEisT0b9uQ8
1zI7aDFW7+dTiPHjyQe8KmbWOGpK+zioyso4pgCp2VP1ThiqAk7UudDK7lE2ftsJHsy5kymEmDEo
6fc8RWALQjANfq6j2bSdaMYrE7oChgEava9uHZdeSYgANn+nC0kvSEJCUdTM0vMBL+YRXFnjafoJ
O9IDX11Jj8xiia1HDr4ImqJY+qAKG2acwDrCTm8ouTv2k4KCBFGBbVPgVXBBlL1vT/ah4yZqRljL
qXHgIjiXpp/8x08zJnam4x/36qUK8xpc0ICIbD6qiEyUfcEmCu+eqPMB4qZmMZ0MNFYJpWjVrJqU
tS1tB4b1YtBYjKjJ1Tga1uiOc6tOJYlMv/lEpAd+2+Nks59NvscRBXVi8G6zg344WDGSIBAjFd0i
CJxlg+W7GyEJj/FAGVIfOW9LB5Q099YJhNiwYK8fboc5MC9iFl39DWGitCyHChc+yPOn1YYHs62H
ypYGxePszrYjN8hq1citPV6COFHFyCji35B42DNZyT6j8cnMtsgqcQWtWG8iTYqtPxis7Dwc9+QW
92dLi1gZlEw8kwOowav3i3wg2dweBd1t9b2T1cjzIIsX1gunGkmBlelVmUJUeTthDxWhgxT/gVXW
hKUs2eibrrbYsuEyXZ9NjMv0j4SOEzff6myr1TfPaCcM+AlrSoV8LLsfZNuhdfwpAhp9t1RkWMVU
99b6Mv72UbI0ajtdO1bVkC9UTyndwVvEoxBfmwJFxDLDoQdOItr7iFn0WfN8JiLYG3/lYyyU8X+P
MxMR6m91ngwyqwRm0519VrDuc3ijAKFviEzy/5+qUTSgYuX+7yv/WKZtlf6lSrkPBNg+yKO4vCNv
NfpgVV0pGOS0atqRiHg4j9HIo83lvnqRc0pYC1EIMdMf2ey6bDixv01BEAbeT9OgZw+CpX/Jl0Nf
MrZCBLwbrexQYVQmPCPGgYxq2gIzAVzdJ/soxwDMRYoswFYzk9h3R3QFzGL8qxFAa7vTcsXHYB7P
q/tOOt3JC49uy2etEap0Ca7rrLz3H940gA2Cn6uv1DlraOveGo0nYgcUpCaGyRZ2mIzWIXSlrizE
zboGVDjfMZgAfugxgj73kROBMk6XdC5mQOddMiNAo5ACjD/XyDQPhiE2z/CVm+7rF330f1704qbO
j2AXreLNj7LzP/5uF/sVooHiPgU4pScj3iRmf+7P86Bf/QKDZEeW/Pn/1H7s/yKWTaL0Agrnrx/a
cMk9rTbreztqw8gUDxwf26KjKF5zEQOQ3DC8xjFy/qUekd4FOfvRWp7CnL/RSI/7T69gMXB4x0fL
v3UUPupKOQoY8eEN2it0PUqKg4541SpjpXY1Ud4iny2Q9EslZ5glj7kQlqvEfCjWPhD1yljVLI3O
auzGRi+RBSZFfSDqjCWeGjDKTMw2tE0FeJY3lBByZ1DnSCvn6zWH1wMgrJiieJmJD15C2Bg+vHpg
CAnsmyYd1wn7XcPU5LRYQdjNx6r/bvYw0GF4m89H7BX34WLZI3jLjm6eV106oZ2zQiHD0KJ2PLnq
8WJzNO5+x4cHGBipoNneB4sJJoDr66wiA8FxkCGyjcSyd/9pP8VkMR5EWh44kfe0kQo9/mzVVHKJ
ZYL7YmSd8OhxY2PxbFg9QvFWYzlu1xzBa4okjCXKNFGqFX21IasUMaujBE3dVno1QvZQ5rR+9mw8
NBOpgCUCyEDnQLFCPbn8JBMfn++Pr/Whz8ww5IZDrwd7lSVDsBxSqGCckq4mz2XotBe121HIu4Wj
MZEFcXbfKWDS9OwncXZqu2E3uv6xEP1P/E5XCBmyYVGx8AViltXacGj0P9ujBnkUdNXT5xVbJGbO
Cx6B/eUWnZ3nTPAfH6d/fCqeHhOASpR5nzeicLWQfdQJ50ypqLsycDupoeKGlnki7i6UY+p4QvMh
c5V5xA76ALSCR54umVlVHwoi39QtkDum927EipLfzhb/Odm1Cvr5uWpTF5fIC8n1oMb81G8wR1OP
px9YQ48IUZLa0jLOJGNHRgcrqqY3uzBSM5Xc5BsxRCr019i+IMG62Fg76KdNQ5VrTavdynHa3gQm
ybeL8qrF/E6kIhVjxn8MlPsz+ygg+QfzzJvRoGNXw8h+tG0R5Cu+K0mbwjw4J5BdwiRHXqLLHWdU
4AUaZf7ymCV2ZxV1MnJvICxLmmByTEQ2bXQf4OiX3apJUFT9ZJSFOFBZiLH83Jy7AICn8v/c0zqH
JKHBEScIjzwrCUJLwaVlZ1vJ6lnfEgXk/EGrkoT5TbOASX4Qj0Y7xlsdarvc2jMpytbpxv3I/x+S
IgkejKgQvf95cJhPsg/Dlm5/5xWbl4/DKVJoRNohWF0feJQ+UbF7kldai39HYR2dI+0Yo2SZt637
HyBXMKK0ZQnCjJcpZC9rp5D9f03OeONR0gKUMdzL5in8aIUSjgoUliTN4+UAPz+OnUGn13rBk8l6
0dM27KFRnXpNDZpJw8T3Bpezkl60p4HEbGCwbJFY5DlWiXsocItwKBQ8J97VIoP0Y+51wQZ6Kkhi
+0GkgS5OJW5fZI2S5u3mTPh7EbtfyTm+0AHvOIC/BeQ3R/OqG3A7MfKKFakCBuKHVj1LuXJjQ2I7
bMC4DGwNkgq8h78ITcywxACEqL1nLQv5D55h23rpFtF0BU+0srNHU6ROm+KIDM/UqPGInx81YU+u
8IRKLmLf91AlrFu59AZSXJk52tXGNOEsTvwtDDWs/nm8WcGEetaNl+H+k3o08Hfgeb5Zppx1gevs
xpXyj/4B0NhtVMJI1cJuRdIqq03GA4ymZMky3Q+fQoE08bNL19nu9ES5+tBSsycHdwdVVr5KtAlI
Var4Z87/B63RMKpi/9uKuR9JLy34zQCRvUBDbTqGtLb40zs7BSJposv9a26HK2ltbbD5Cenh0zz8
gedFFVX7OXkQRNCd/PwXOfZ9VyFgcEuxRRGsmbyRfHwLcV5yGK4+cst8WcX0Ec5bYrnW6X9mUtWx
1F+oB0ZZRQOa0ZVkpodCRoiScg8N3vNWjH4yW504KO61bOF+mwZ5pzLonSpakP8AmXHyDeWGjwih
NBvY9c0irxEyi/ewcBJ6lidL9aIlyNpcjzDezQXM3SJHRvYraWK0sB46oMsZu5NEnPm3Hsd2G2qg
kweLuGQEDaTWn2vyby47WEV/HS68U1+FaQJEXmtb6xY3CFOrhFWkHC2kjG//AXcgk2MlRpagnZ2U
TjofujB2S7n825Iy6nIEHCj2R0jZyHYsHhRqoRX7Mi/0J6AePjuW1JYoHiLYKvb7a1dm/RGZearO
5JiFM15rE4m906iO7KWXF5QtUS2v7f43nveDpgrca3qbmc9kON40Ug5+YEKB6qRJD5726MjDXo5X
2AOFRTsWj/SRiN/XSqXIzvFaX0/uXCAQUxEEst8KRFjspyVCO+y6UOqaNuWMXpNYs4uRxblLBYFY
+FumQNv7AIQFRg7l8lMh619xo/YQ5y9P8/j2bI0Ec2LNwjPU4N9BdIQ/TVKurmJKfKRiBqzdKASO
xMX9D3TGtXKy7YaRVpJr7pejhFK+yGU2R2G/VtjGZuHK0JaHbYGW/X91MUKH+t0lggxrEYh70xj5
x2ta9QiSFxj5Kqs5Xdrz6RfceJanCGqGUijVaI0ccVY8mYwKBUtMGCMjw3NEPoszD5IoBLwwDrt8
09Qg/5j2YJBjrWvvYFcE3wKfSmTCaXx5NkuQQ9lwEG7k1C5fnMOApiPoyKWuHzU4I9lC8xL504cy
qqZj3RUmPpkECT+t7v95z6EylH1OL7RSjhs7nWTcnAVO82pz2nd3C/a079QjaCXVbDX11VUSXc0k
vytiCVMWxt00e4wj64Jnx2d1HUKMxC9WuneNwEcVczIbIlTku9X1erfnzp7JPYitQtkjWQm3RvgT
A/hyx55nReS17Q5G8oHjAH8Mzlb9bD7BDWMQvlikVpUFxC0StFpABHiSuVfzeE/rVvc9wTbN0BKN
A8SZlmHDTKa5uaffXYdZd9Luy73lp2vVy4wLZZovjoyryt6wP8f2MncMPjwpjJjd9e8QdM/7meLL
ZyHjgQGGtijZzTETqJmdNOWogkWq6oN4TsO3FIIQcEhbngZ/FXmEauFuTt3mLYxdL6KHmWnscbH0
i4oQwIN32Sb8RRT0Gj2rdSdRf+sceqksk68f+FgZE+SpzvyMbCiSfQ51MN4YIWHLJLX9XlhV3AOU
+IoVQNLLG5XC/PWvQ1Jce/s87hZBIT86CUgnGhzcd1Q7hk9zzp0YdY/ydHbyJevSkPXP4NpYnf20
K+RoNYDkVmb0MpWutc/dlTAAhOiS6r8JlEggoqCDjnmgiRXmSHOKRwU+LhPxHgvX7wbdtOaAYkEB
VZj/NOXiL5GWIIXCicRrmrOAwrs5nvnhS4KhugojRZaFEUtpjH+rZc7KruMnexHwFY0WCrZx257l
PiMoOZKKaj6iLi+pLeUEk8rH2/XaGb9Ef0VRq139Sj+SASuQ/PXtl9JxBpdlflOuoQOeGUGGMCZ+
OEuwRU3v7o6yOQgwKmSXoCUcXrxAS9deVF0nnBSv1o2BsyHBrsb956LlRDKRuiOWrt30uv3k8Qqg
JVk+kprEs27DWf0eF7plaMTwcqHxMP0dJgq6dJ+d7CWob3iwda4dQEpL1r9nCuWE/gRD19i+XZfF
TU09o0CKbIwILK+A5rtr4qSlqz1CMVRYQ+Tq63jl2F46miQ39w0AOpQPM/DIj6A61PKMloiLQYN7
tDyCRnVJ4cvRwtIy90SXgBE5DcdIRPsYiHSjN34+9Lc1eXbz03HwqU7xb4PHo/o1WJaZSJBRwaRr
85EulIokGFRkBp7Y+r9mmSmcYy3/k21l+OIOjijDNJTwKmKCO7JMF5apn7j14DF9EgShYj+h7BdH
2w5MFujThpT6jNXpYAtauCmIRAKgFslEt61AvLuSwQf6tkZtnQUrQxWpbv9a2jT72kQu4EGPBuGt
oCVhlLMdsqzmz875qri6JQqqx3F8fJPidr07erbta7c8ihPUlUqaGnoQ51OxbOx6HcfP4DxT6TeJ
O9r4c5e0BF0b3jow0G4plogqX1tbyKaAZEdZDoW/S1RH0cGz2vOkLdN0+kMTYRl8aufFI5t6f3q8
ZgAiy9x1ss23qydQ9OLitZodDdgnzhDSUDO1JTMRHUCDGc7PO8MFZhkFxlZrhUuiUc9UrvbiVPFQ
WEqfgA3BpDXhdHWmkztpe6VFbqQlgSB3426WhBRisDA4EHsDHsAtucaBX0QNcjkhHjxgfAW616gQ
jXSJP/c6amP+j9xU6ec2NlKgo8nq1KEgRzz9KkaGDyiNK90mnwEaHwfQ9PoBgj4W6Idgs9TmPi81
nwe8GN8C1A2zLWoR5EiPs8EnBxjAtZYMXoNnOlST718A6Zf/Yb0AFbSliNnyvt1DeITyBvD0WJ0G
vFEWWU3S6e56SEJRBgXXihPJ8g6D/KhtYlv+GG/pjJo+LCxCeNFP2QUO9RdwW8VzNFMlHC51FaL5
edqhnWzVrNnc54fd2xTe7ouDWSAJKDRTnb9nZFYmGiAJGgkI470Ni/9Re1H09gnlQeh+whfVtXoD
PtA/oLy0X+HM+usOtwHUusbHb9DbVWqXqFZStFpRSl+DtsWGCo7k3wvkkGzF1FnOp01ODlNG5ksP
owY34C3Vwu5br37RWGveRH9MibKfumMSEixUPuC96wMNNamn7BPzbvYb4OnMComT1H1w4H2aYLYq
lIZd6iA9/gcHn4CAVrNnolOuPdR9ETTN/IJDleWDhxx6z2r3tlFiDf8Ow5aslZ/zCNipSAZ5ITte
GkqixWzRTxNQbZGNABvflc7fdp3kvwZ5K/1crsjqwNVOVYmmlq7vgq9P8/ra/Sjr/pWEevskldMY
sAIKUh+aL45FGAdBzwmQq3XQ5rzkYvASs3YtDwUejtDnEw5zb+doKqAqGOqejtci10jbf1Ll2SrX
GHMFCHDn0djwcLXnm4Tco6CyfQZnccCLFgXAn92oEnj/8B0qt5bSsQlWUUBemXBuhYBogS0q4zjH
5v57E2vGbVgU2AxdnQXgF+yOS67+cUnG6sPf9e5RC6NOQDiI+7hPwaeFQ4ExrAx4p4EfvmLfsgre
zYogMIKWbcdn2n17DYJvwlxDDqXiUffi1HwXakpxz+cMOvwT60LFy+bEnAUHchj3q7HSKuzOhE/4
3heP1Ok+x+Wlpouim4UQUItZorpVJ8zS9Rbx5mU+EikbjHJFMeOJJ/Ri21xi1aN637qApR1ffzY2
4PtlahRRpieg6yduHBMHZg/zws0CGFxsY6OwoadaooA8TEg4UXRmNgC79u295gEKoT+j5xTRE+hi
EoyDF4uodwoxWx+Xg/rmO3nrpF8DwHcuFP6h6yPIARc+ANSHtX+Qnro/mdvglzmm5dmzgLcxp6NI
8ejaHFJyzEXcbhKzSE4M046nKcyKf63m69tdh03/9GSY0Q4O7pgceAO7eohkW0dPSj2Asfh4KHka
VG1m5RAi5sMwzl2OF5s5abswLB2i6qMJVyRqGIWGQyw0MkaziK0mL2jAZxSk5+a0eIPK77nHkr6o
5L18+OoHCfyo53shYSbYqDfDktj3teTsBWwfKCnNX2tt9lTh1WPV7VaJF3tcoRWCMr+fXr3ZhbP+
IRZKkqr1eL8mRwJhuPEYOGvmN5PO/1vU6oa3enVBG3Hkc8oQZGtzTE5KY5Yx4rHGK9DYMscXxtW8
0hHz++5ZPIv8DsvELWuifhxL92BQgPsgrGvKpIfBjZAMHC0/pu/+4snsSaQo9baajFlXayRaBuuu
VrpAw9Qc4x7a030wlOA+8GnT16Zdvtz+w8OUI5o4p2y583/I2z+XAyKITAQ+T8NgIfCl5JsS/bKR
Ab5I3ef5P+2heHNbraj7S+xrhuHkJtmSMDj/LJ5UGQMCSyZgQedWOWUqWv3DsO0bgbQ3SZjLpoKU
cjfvgnHsttvsUW32gUjQzajdhKvK9Y2Hs/mhwWgV7xgDd5W4jva16ehpohDG3KSL/O0MgemD1eRu
PoVZlwcHGGbmJ7al5scp6DGY7WmAMBC4oyhCotowXiS1KtPeW0IEkDRsJDAgUAFDShFjIvcVMqY2
RAJVow4x0qQv87aZN9UmY8pS28aohSkrMsSMP2T6+IFl8a1bBpsFXEqy1WXA3Fmu5yjetQJ5PYk4
6EP8YFe7SAGgiUmA35YtZaP9ysXzPiuKLfNsIjy6BIPVFMVfG3qWFyD/05IwacPSOjDqJshXpq87
k6aS+Y6xtBNLCeWt8pD1l1WoFwlKeaH5vGutC8f9qfuiAUsw8efspxR2QMdAHRsw6HVoFtweU6E2
7WRzrNLNsu8/sElqw+4V0jlBeWI6D7QPkNT3xMrtMgK1On2+281uJbhl37jzl1rF/PSKbzFC9Snp
X1nzMhQMI5IFM0flDNiUFQryfCtvodtvxK3/EnyUy1Alp80fiLanETOu7+chavVylyDFHekMqh+r
bI25rzBfouPB/T+k4MZiNBubMjoGXmm3LEMVMzr1iMKltQZDaM/HLp0GPJWbRBajdtMQi/yWEv9r
lJkyY5M9yB4+ux4uHAaIQBpUE9MP0qKPFuU1/jCACkxPWnbGzdk/81vy2Yr+nyB6moz7JBU/wJGa
pwf/GEsHJD32SeVgRBy9hwQVx7NS6pLpRoXGQVikKTop7VPCObP4v1yD3rmTe7sva4BM5fDiegEK
ekaoWylETQuRoKtmaOep0+aHIObCsKEnzu2yurN3ysdyFLhLNjoLlLvrgchUFeXCqwLBsvmP5xjy
1Ou2MJwux9d/UQY5s2qORLj9rJVHnvfOPrUaW5T6JsNr/QQWJWM/8q/sMKK/bT4oVT40HXAsBzWh
AKINTaz+XQcCV4LmANNf6qLelfnGE4Ung22U2f0tLeQFsyWCMoWTR9VzWQKEwvGnT1q6PiTCEPhO
Klt/KLDP1S0Y9nEz9Zihd9pHcjtmZ5HsygZlSxdGM3fWpaAwf8sW9sIE/yInr+COrvtvS+i27z4q
iNp1+Jlh3I0vQY5yPNQI3ZPJZQ5EBOi4Xp5otyknjyJEeF0KocBwlKtVgjZ09RVNUxczaARk7dFN
yZAE2p069vDc4Ahn9jHC224+U7TOBcClO/wDqRmLlboS6aZgfOE0g0hIvy1cM8nFvgtz3Zb4Fp2o
9WHz9dcEhyepyFkqwqCjxbFSIeV7MPzDTYEmgK+PFlPQsV+B10NSJ3zTBF65h/JI2Rv9/IbPuRkp
tbsy2FsTF4hRH0goSmMVtev1mx+Ax6+lzqUgCw1l41iEX/ZOM7QE9BDYOvGWyj9O2Nm711FDFRxa
kE0MvW7Waf+34pYoXgQ6s3LFA6wCg3GLD1ixBVeyvMl4bq1mL8NDoSw08qOpoaeFOZUp8CzEr1nk
0GUQAK1Z7YKAx/1TcZwEXWZlLKXu5VQK3OSaQnTIdiiL1cAzbVVZYegbyJYvE0nz4nlZSzlqT5na
4HQQJF4vtaZRgSz7qnKNt5WNHtUDFlNV1mkre5Y1U85D7uy2OkT1aU2KWDRBu1v/1O9zzDheV4LL
m6mgwZ3rK/LUnOvzag+dyvQN4fWDxwUn5jTnJpqpQf39zthEo8nv1x4p4BBKRGs6TM4DL1cpBr9k
04U2vS8rgrlyqA+03phkG+ksbptGscq3gVvnaUdNzmyIqkm14NRx+HA6phiThVQcXh54qwiF+aPi
ICujeNB9sslwLSDRNEnL2b6cQGN3Tf7pMjBCYNmA+7F8AOL8LZ/0K7Kc+nausxwq1OAn6xZVe5aa
TzvbR3G1BILlW0lqPyjnEVUlgPJx5vCvsIGwH5g5DaNQJ0Bg7TTg/DVfQNoP5UKONXqfx83SX/up
Ij1C5OU0uNS5xA42dBJTxNg3QyRqPW9T17nO3fL3bahtwwViBbPIZWuFtfunKR++rIXFBgv1bry+
zuGGuEnHJZ6B77A/xo/W/AKa9mYvEw9ocRKT1Rf5yGES0hJvTlxrRmUwKj0wNDARLMgZT03MXID5
y4zkUBpddRi6CQxZNf4SCZaD70ly2l90e70zVaC0tcjABhbNB60YPL7nLJEyEUskurZUnKTc8tbL
Q0Ql28QfHlqWJz+dXIsnUU9R3tyXCuqpAVEQK/1w/MBNXiqL/yaJZIi+c3ZV0onZPJEysnN5ydL5
erj26WrsHNnOx+9FaOvmft+VrzNYZ52HuUxGjXSOrKF4tty4g87eHUbU5dUvd+PcA0KuwhvcgIye
xpcWyIArcCbrr75pwhrR334ypI5PJP6hgLpuoGaB1EpM+oiKa08AyGBDuXZMzgkOxm6QN0BYVuTz
yvDwjlX0jAXS6sQS9BPHIt2Nvhaum/5jFgmNNRG1qOZv3+/lZRc3wZhbKdbSg2FyUk22jK/AnjL8
rfH0RAphsfh7D4UDyvbWE9ivuE1hh+FNmTvGSuTgz5tYhYINVSDTcAJwRtpH+S5jb4H7PSkwALot
hyjITrWYUVKYmUBaOu/pdHyNCLQAqCLLSdOsvc7LcqNDWiOodmBiZs+oLjxp4Qjihd82pgYnEagx
auGIaLKJcn6GQavM0IEsIoUng7Cfd9TT+T4oIDJ/aA7EkrDvBDO3JTx4mNUVdy2vKKaBs6w53T7U
3Hqje9LlPAnn38bY3a47/fmYejvy1vJw4UBCbBVJBVKBT/oVL/m4RA1I0O6n4Xp8cmJX/Dyy1agG
ohw0Vka6Z/eSBe8FPWpeBjQ+J/rCrK0W29AyVFDzhmNv8mcoAikyKMwQm2Da0buS3JKNk3Q67xWX
Ee1/253lO+X02RyrbnAwrehaikj2jygsXGSvdiQMXqZ9Sj3UL1+cqxCZDbbtoeaG64s9uTWTKzWx
RD7juSLJ0BK2ZW+oGy56UUhjJk+hWviPu+r4K+nMkKqwT8Cq22o3ypBBqstUqWRFEt1TT/BMx/3m
iRF2l4hZ1/sfxLmUnTfu1nlFgzb3PNB/HSbD6/g/kGSyp+AaoS57cImOKbXauiGG9WpUp+NoYLCQ
orpMd1ryIELF8ZXXWdJd0EFHbSq9IOda1nI3HapRiTPaFYO88s+xJNgZT7HyVX+0gNs6Cv8Qm1CP
eIXp1Q/7G5Bd4ddOqFddJyJ5aUxvPz4+GT2Y9ljh5Zw82iELApRgumnpHFO9MOMJZn2300ZmrCb5
orRsOOpoAMMMK7rf7RjVYwnPWUlppoFXD8VakHgACQjZrYyE6A4WRAuOctX2sye+68ww00908pnh
Pg9AzXRI2vr3JVfudt30LPMzvnd4Ye0BjMT+9hXWGfhcn5ZROmqi3tsx6QphOO0uBbyH3iptsFYW
o11Tr7MZFPT/kXXFjDAkgj7yXDAeVV/bmyleQjrikksij0qCvadpojjoAWgoW9eqroZ6JYIi/uX3
ivShOr4HlUK4AGnLhRqLZzDZKuLFFsuE4RwhPiXDcaxshf1IgP1wue1BTkNXuc2Eb5QgvAssJEPS
SBUjXUVi+62JBRjv0+tAdEz4nazCK6Yu0+LAJ6nCbSATNKOIryv8Ev0Xxu72KC0Nm195l//MkoMz
8CvpmkYMJRdYGnf+iOcGFNrx2lqkSoBk32ET7OTXt4WSDkdUHxP2coMrNBHIEi112s9KkYpjEK02
gX4UcjlBjMPbLfTE7HkpHfGA/1TXZWCHM4K6mN6kdixspbyLNz2QqJGDv/4y0wGbumIT3LlNgKiv
n0lhiM3d+8LsAxpa+gb5y8sjpiNmXZ+4k1WyoJwqkaR6/1kRQXfIjHwMzNoX0zoUv1MrxtUOUjSC
I7h9YCzriZCHfJOYUZWBrbq2d1FF1hi6/9+noCZKUQDdelA99s6z3U+W6inRsSsYkEeSmxc363+7
TYRLUDI9uu6rNQDg0WLo1ZQFYRQkQp6tkdqxRf/ujLU7AJFnJD2nc8ZhFJ6MOWRqE7lBuMI/3Gvd
gePm45CxyT4vUkwKOvLhpelADvt3XV/SaCPxNqI2AGbegEPtj08r8vEYTuFrKBs7BTyPIO9yCKUi
mE6rhPcEmXbUGXE/PK5IZcN8xqr4E88g4EV6w9lYe7qttdTDTNqmaHvWJYUG3wyk2f88LLVvFw/Y
Lbxh+fA+RHe7WFB6Zm8XGZ2Qd1XlJyAZIro4RJrkceN3JHM1vqIjSIRYaHw097BDw+jYR0T2ZVp5
uEJLMFQ4om8yNYJ4uqQtIlScDEClNX4nXF78m8ogHtcG8WM9SkRb9RYe46Z0k74n20OoylUPBg7o
xlXQF0gN1+GezFKqnkFNgqtUCHbN+PZV7jzlGk+lbBiBpV9k2fsDtQUOiB3w0PGCZoT05TtOSSzM
R0XSLjrdPieZodLoKqMmnxDn1aP8esmC28bmwrlcurvu+QGVtxbfMDLy013A1e4cs3am7P6Auf+b
doAnR+K999JJQCKoRlTEyE5O3w6M7AyNNXwqpcQWNnUItqfA1AWsGIhHFnKZkiWA0fye0o+tp9r2
8risNrzvjq7FJr0xGxH7b+yEvL2WwKXPRHGiKodeUUtn0OA1PJkTuVY30gOc5YFytWTZKO7Q5QJr
2+C6ArcEHiSEkxZoPPcUgs/mex0xPz7gzkS+MfCJgsr52glvb1KnQXeZvqW+YbspcK7KQbNzQgi/
4SN0KCz9CB/2CC/D4oFCOzroc2FTivpJtlbNxlT7nI7cQRvXFjssiaGaIYHSyaROsMrPmqY9lg6F
OiyM/fhyc07n5VJU9/ffVsKtWLdwhcdTOaYk54XM+p7p/AnCLLYkI5cWGI72ikmJcB/dWqfcMycR
3P/Fuov9t3xUKV8PFPyg+wkV4cBu5HKADNmk0CvN9lkanfMeDsobGtquyT/OaUKvxTUquARC7pPd
gZBDl4MYP/5GWocLJJcqcERxXhaQhLVOpZcJuoZlHyO9KssxejDR/zSUjRgS9vQu3ta4v1UjLb+u
r9q5wPmyFv3gL8KmesA64jTVIpbotf31fX0+tDmqiOu8nD7lfb4VoZqOuDS4rwKP5e2PaoqDHXOM
wzdvTp69fRVax2nRRvIPzek/iqm97SJ55qsPJ8lr1D6wSt+ZCCLUNi7syFVrUOVei72gb5ISVvId
jP7YPTxg0IWKGEtjWeqcAW/52Agz6zvtVIg9YCv+WoYcoE10mbDoVIscz69cBqKeEPfx/IFghDou
389DbadW1LhbUGYVWpBXxmQev/AWwEsFAGqGqu/G86GaQUsKCf0o7hYGNQqiCnLO1OHcUnMguVBH
CwrXkxyhG/7WKbzC5+Il5N4IIrHi4trJWCSTD8XMp3QwnEmGyUbvn6tSO20jtlQZMz7U8IznmH5C
LSwT7pMDenq5YxBKXv/neTsMVTnH9Ibt2rwlNxR4ascvSSPPOtNRGBO1Afgr9caGf+1vnDbpZ+JD
U8vhPd0NK5+UyN+Xafk9axCN2f7bo8RSg8hUwkpB/g+NAmXhsIMNOVCmgjA5BVydTMsOM8lgMbd8
tlqmJp58ok8+UfBCNnOKVLuXyd77DhcIILyBhauqs4/g1iy7AdsUFk3nnr0p75/4YG0YqGP5dBGb
a3CdvEyH7b6Jb6Yja4+WjXmJ1AoyxFogTA6in/BMLJMKwWKAt3JSiE7bf4MSpwvOUZHfE2Whti85
HoT9XTmBc3mFnanph5Dhq3xPMcI3jPv8KhmV1/L99US1fO1n4YCXHV6Z1KHTtGHxExHzyT8hV7b6
KOOZW7zkXGVuOPPZ6JhIu73dXfP9FahITPw2qhG1CsdoaR9idQi1KRmOKz3NRxjSw/wjFu1xtSoj
2fCiGWarnZ4mDcKwFpr6TPhz+uDTDXGbEBbfa+oxnO2AlmB1YjbRIhefuC9hmLyC38OaocHAb80g
+XBO5Iq1BbJnKmF3GNXL6M64Z3iH+99dXULc332CQeM4mgiAYye3jCiTxa+kktDkXpqF4maQImKn
58oVnm2q3bnwtKbCowQHJNrzvHk+Wn4r8pitkXooq0aJG/hTQqfLGRglRTE95VE7meKtdSiPpyiQ
4Zyc8k8hyLMDsczo15hWUXiFRM4vcRz8MJMp6w5Nu7MRQ+LDjkbWl1Vh1aUJ6MohhAA9OuPwgmW7
8/Ojw5qCZFDpWG0B3llZahA6ZsxDPgvH0H5DlRwLUYxRTkxGOORMQYuMQWS6S7dSmhc6daw8IHnJ
h16oBzecQSPzTCHnjsgH3jIB2iNz//zykEPZ4sYNcu1sIJX3VSiG7lD3P0wmTuJuhnDJVV12Sz/N
6206jczO3AlMLMWKOoql6+RykZDXfnz1FI+RmaID6qV6OcbawtLymQbsxsw7aryM/EfE0sT1CD8m
fEEMrnrp4vuj3A6MsDmtadAEAZla5kJLjAEHjgmlbx93AQ1WKrxYVpMQz4K18mHIiUE0u+kM6+E+
oLIEQbrLwoDJmJd2rvLVs6hg//3xuuN29n/0cXrjTLP66eRv/NB64swj61JulxSjKC0t+fLcQ7J6
sKX5d50Jqq52g4yuY4xS7xCGHgnKA0XgHB4gXIk3EWXzw253KSWkrfS6DWdThNeb6+fReKF7vJ4r
1pJGre+h+TL3rvwFTdAOeGKNLomrsjEYjryqx5SnvA93PYJ2NY78PpkD2oe/lafAQQTyRmQ494FG
bWodLFTkGrXl0qWcfYOGnFuy0Bb17tx29Mvr5Zny2MbylKJsHOo/eZEJRrYwDVVSnmtQJdLLXP0e
AAjXXL0bS0bw4TwD3KImOJw4hhCbW+qARamofC3fNODUsCwQcAWa8Otmbd7BSEvluO72AZaGMSPn
4JtI7+nH02oEqZW6cMtaFCfrGqaHlmcBNO12MMEUvC01+7byNagvMk1YA30tuRTGSYUtsjkDY1Rt
2h1AGZDgqlLzaU2rcrk20kOCdsrKeX62auBCVZQavX403JXvsNOX4iYmCVMm17hd/WSfbdrPIoeu
5bwVjAIBd6tJwPCRxwQ7NxgC84QbX9xrRcUrJ/b8Rk8YUDW7g6BeS4Xjxbyl/fJeeSdjALEOqrO6
bXr6RnYP0OiTH9QQx4EGq2u30IdwCBNzDbgnweWwfWkfEfCX4uQYQHoM5aB42IvNhHReiDsIKwEd
gbl6XIMp6piy6W1kCLfOG2tUbAeSsfo4jIwpZfyp8R6tohQ+UIcdC68WcpBVnxnVs7ouCVi+yXfi
mnV/XIRbdJgjELgzqAmdxAxbE953aXSZNNJOrLhkCq81Bc5Vj7+GhRha6mNw/ISvZhDfNL8jm46e
1euWphLNzpDWrxZppUcgX4iEKUfnf0NnULbulTAJsmH+kSrvbQmqfXClkweX5obkUP9i0VMbkYN6
dr+Mgp71b9suqp+OHTqGzDkgUR8MlNlvcIJ9y/gfx1EP/q+qGug4YpcVVMuARkwUTfd/41aTS95/
A4vBKd7lNJ5CiYoKokDXNYngi7kuYXvxYGUnm7CdM8iAC22ky5WcrAQCtdH650GgPJMR4tUr7XLN
8/+XdTh+3JsQFC13JHXct1uPm1xdutLL4UlzbMC0vpPIm7MFgfpRkk6SviJoBg5YZBmDSS1Egzt/
MiX3Vy09iLGCFIPAkmlGYxw6zBH+ZCLs8kw23UAE1VMdpJyyq1JEnatxvyHgqLnKQ5fMb5WWOJCn
SYgAH8JMXmmC/r8prAMSCoZJ03F7fsgi5nwQstmvlA7Lj7HCjibZt8AMPPii3OLNOV+7b7oY/sTk
sTIx14FpZ3LOoqsAOGyyHIJS7VUGtLC+ruvMWO+t5gk6RWcNQhGpzfbtxg550vquLqiDz9i5b/bO
ROspiBd0CCMudXb+QRyTNwh0WPg9pNuDuRtVALH/AR++sHAiA3Lk1HZnlYPVdNf07Qdlk+HDYv1q
DBwxgNppdMmh91c5Cuk/LQ/owhxUAPOVv0b+F1fkBcRXSy+M3AdM245ABACPtXNYKQRYlG0kJ34r
spGKgERL6XRsik7n5O6twnkJ4GPfNUpM7eLv4IfaCRYiUWyt6btRAJU1ieRs/XuAoq+XNxUvzwTP
TNXYc1r3REJqynjtYGExqpaN9uR1CfvAlC4JYVbF1+Je5npnoiiZ0o7vCyYEKLdkOU6zvJvWV54=
`protect end_protected
